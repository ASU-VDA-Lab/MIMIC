module fake_netlist_5_2377_n_1706 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1706);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1706;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_73),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_89),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_97),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_45),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_5),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_34),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_144),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_26),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_68),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_28),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_42),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_20),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g174 ( 
.A(n_111),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_57),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_54),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_25),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_96),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_6),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_77),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_51),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_50),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_53),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_87),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_54),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_70),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_55),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_50),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_10),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_11),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_5),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_33),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_40),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_45),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_24),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_105),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_85),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_58),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_33),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_75),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_101),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_137),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_10),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_27),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_103),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_48),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_12),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_149),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_37),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_106),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_18),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_126),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_102),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_92),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_95),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_56),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_93),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_48),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_30),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_43),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_141),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_123),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_59),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_41),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_63),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_44),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_142),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_19),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_121),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_65),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_148),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_81),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_104),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_49),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_138),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_117),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_79),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_14),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_11),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_124),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_13),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_127),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_90),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_19),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_78),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_18),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_24),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_21),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_39),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_72),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_146),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_82),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_131),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_4),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_61),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_56),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_112),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_135),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_55),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_69),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_38),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_29),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_99),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_114),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_21),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_159),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_160),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_0),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_154),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_181),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_169),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_197),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_168),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_155),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_169),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_177),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_186),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_177),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_190),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_156),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_169),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_157),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_194),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_165),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_163),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_179),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_251),
.B(n_1),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_194),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_228),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_190),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_187),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_255),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_212),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_166),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_212),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_228),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_215),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_162),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_253),
.Y(n_349)
);

BUFx6f_ASAP7_75t_SL g350 ( 
.A(n_249),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_253),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_173),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_215),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_175),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_176),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_185),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_216),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_191),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_265),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_279),
.B(n_1),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_192),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_241),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_241),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_193),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_216),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_195),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_286),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_217),
.Y(n_373)
);

BUFx2_ASAP7_75t_SL g374 ( 
.A(n_249),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_199),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_298),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_241),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_203),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_255),
.B(n_267),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_251),
.B(n_3),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_325),
.B(n_277),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_267),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_307),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_289),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_309),
.A2(n_223),
.B(n_217),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

NAND2x1p5_ASAP7_75t_L g390 ( 
.A(n_337),
.B(n_251),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_316),
.B(n_289),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_251),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

AND2x4_ASAP7_75t_SL g395 ( 
.A(n_314),
.B(n_182),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_311),
.B(n_196),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_309),
.B(n_263),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_263),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_196),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_158),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_305),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_323),
.B(n_294),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_331),
.A2(n_227),
.B(n_223),
.Y(n_415)
);

NAND2x1p5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_220),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_323),
.B(n_206),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_380),
.A2(n_208),
.B1(n_243),
.B2(n_301),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_374),
.B(n_174),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_336),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_367),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_330),
.B(n_220),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_367),
.B(n_305),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_330),
.B(n_219),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_349),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

OR2x6_ASAP7_75t_L g439 ( 
.A(n_374),
.B(n_174),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_354),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_368),
.B(n_221),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_226),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_377),
.B(n_378),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_317),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_427),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_426),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_426),
.B(n_325),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_306),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_425),
.B(n_310),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_407),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_428),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_428),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_395),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_425),
.B(n_320),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_434),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_402),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_415),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_378),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_407),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_383),
.B(n_329),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_383),
.B(n_332),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_415),
.Y(n_480)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_434),
.B(n_334),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_344),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_336),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_387),
.B(n_352),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_396),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_407),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_439),
.A2(n_365),
.B1(n_391),
.B2(n_387),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_394),
.B(n_356),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_450),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_308),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_382),
.B(n_357),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_395),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_395),
.A2(n_342),
.B1(n_283),
.B2(n_260),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_444),
.B(n_335),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_395),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_439),
.B(n_324),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_400),
.A2(n_342),
.B1(n_365),
.B2(n_350),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_382),
.B(n_359),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_400),
.A2(n_342),
.B1(n_350),
.B2(n_328),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_409),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_385),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_410),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_441),
.B(n_328),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_385),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_385),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_411),
.B(n_363),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_385),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_439),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_404),
.B(n_366),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_411),
.B(n_371),
.C(n_369),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_416),
.B(n_375),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_379),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_397),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_439),
.B(n_317),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_409),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_414),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_397),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_417),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_416),
.B(n_277),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_439),
.B(n_364),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

CKINVDCx6p67_ASAP7_75t_R g556 ( 
.A(n_439),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_439),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_409),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_403),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_424),
.A2(n_376),
.B1(n_372),
.B2(n_161),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_397),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_410),
.B(n_431),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_399),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_403),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_429),
.B(n_288),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_403),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_413),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_429),
.B(n_222),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_405),
.B(n_327),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_405),
.B(n_264),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_399),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_446),
.B(n_324),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_406),
.A2(n_347),
.B1(n_327),
.B2(n_244),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_431),
.B(n_347),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_424),
.A2(n_282),
.B1(n_248),
.B2(n_237),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_413),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_431),
.B(n_358),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_409),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_409),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_399),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_446),
.B(n_326),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_429),
.B(n_224),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_429),
.B(n_229),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_413),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_429),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_413),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_416),
.B(n_326),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_447),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_388),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_388),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_416),
.B(n_343),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_445),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_390),
.B(n_232),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_388),
.B(n_318),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_399),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_388),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_445),
.B(n_164),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_399),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_390),
.B(n_343),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_588),
.B(n_390),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_452),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_472),
.B(n_390),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_406),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_570),
.B(n_388),
.C(n_319),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_452),
.B(n_406),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_532),
.B(n_406),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_506),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_589),
.B(n_447),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_516),
.B(n_406),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_504),
.B(n_388),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_498),
.A2(n_393),
.B1(n_445),
.B2(n_238),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_504),
.B(n_170),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_586),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_534),
.B(n_393),
.Y(n_616)
);

OAI221xp5_ASAP7_75t_L g617 ( 
.A1(n_595),
.A2(n_198),
.B1(n_373),
.B2(n_355),
.C(n_362),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_453),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_600),
.A2(n_178),
.B1(n_270),
.B2(n_262),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_457),
.B(n_393),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_529),
.B(n_393),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_534),
.B(n_393),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_492),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_SL g624 ( 
.A(n_576),
.B(n_172),
.C(n_167),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_453),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_451),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_455),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_471),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_534),
.B(n_162),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_557),
.B(n_162),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_529),
.B(n_445),
.Y(n_631)
);

OAI221xp5_ASAP7_75t_L g632 ( 
.A1(n_595),
.A2(n_373),
.B1(n_362),
.B2(n_355),
.C(n_246),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_557),
.B(n_162),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_557),
.B(n_529),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_471),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_483),
.B(n_484),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_483),
.B(n_445),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_591),
.A2(n_590),
.B1(n_597),
.B2(n_562),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_492),
.B(n_318),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_496),
.B(n_502),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_484),
.B(n_408),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_528),
.B(n_180),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_578),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_487),
.B(n_511),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_545),
.B(n_340),
.C(n_319),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_487),
.B(n_408),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_500),
.B(n_184),
.Y(n_649)
);

AOI221xp5_ASAP7_75t_L g650 ( 
.A1(n_515),
.A2(n_370),
.B1(n_345),
.B2(n_340),
.C(n_246),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_473),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_511),
.B(n_518),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_518),
.B(n_408),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_591),
.B(n_162),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_475),
.B(n_162),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_539),
.B(n_408),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_476),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_562),
.A2(n_396),
.B1(n_303),
.B2(n_226),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_475),
.A2(n_303),
.B(n_280),
.C(n_262),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_539),
.B(n_408),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_480),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_502),
.Y(n_664)
);

OAI22x1_ASAP7_75t_SL g665 ( 
.A1(n_477),
.A2(n_231),
.B1(n_188),
.B2(n_189),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_480),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_476),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_541),
.B(n_396),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_589),
.B(n_447),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_541),
.B(n_396),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_488),
.B(n_396),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_462),
.B(n_396),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_490),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_482),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_456),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_456),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_573),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_598),
.A2(n_396),
.B1(n_235),
.B2(n_164),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_575),
.B(n_345),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_575),
.B(n_370),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_535),
.B(n_200),
.Y(n_682)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_477),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_469),
.B(n_396),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_555),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_508),
.B(n_396),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_509),
.B(n_432),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_527),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_542),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_548),
.B(n_432),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_540),
.B(n_162),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_552),
.A2(n_233),
.B(n_302),
.C(n_250),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_551),
.B(n_432),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_566),
.B(n_432),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_599),
.B(n_432),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_599),
.B(n_438),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_599),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_598),
.B(n_600),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_571),
.A2(n_233),
.B(n_250),
.C(n_236),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_481),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_481),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_559),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_521),
.B(n_171),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_573),
.A2(n_257),
.B(n_302),
.C(n_227),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_571),
.A2(n_281),
.B1(n_258),
.B2(n_261),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_489),
.B(n_438),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_481),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_569),
.B(n_438),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_556),
.A2(n_242),
.B1(n_280),
.B2(n_300),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_524),
.B(n_538),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_521),
.B(n_573),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_573),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_556),
.A2(n_271),
.B1(n_239),
.B2(n_240),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_463),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_521),
.A2(n_296),
.B1(n_278),
.B2(n_287),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_553),
.B(n_162),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_582),
.A2(n_270),
.B1(n_247),
.B2(n_300),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_559),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_495),
.B(n_162),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_510),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_510),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_463),
.Y(n_723)
);

AND2x2_ASAP7_75t_SL g724 ( 
.A(n_522),
.B(n_560),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_454),
.B(n_210),
.C(n_218),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_583),
.B(n_440),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_582),
.A2(n_183),
.B1(n_247),
.B2(n_242),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_526),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_467),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_478),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_536),
.B(n_418),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_479),
.B(n_201),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_526),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_495),
.B(n_447),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_467),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_530),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_481),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_530),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_486),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_495),
.B(n_447),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_582),
.A2(n_275),
.B1(n_214),
.B2(n_171),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_531),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_531),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_495),
.B(n_449),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_584),
.B(n_440),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_474),
.B(n_440),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_474),
.B(n_440),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_486),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_533),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_521),
.A2(n_214),
.B1(n_183),
.B2(n_178),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_512),
.A2(n_225),
.B1(n_304),
.B2(n_235),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_533),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_493),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_491),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_491),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_464),
.B(n_244),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_474),
.B(n_485),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_493),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_468),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_494),
.B(n_202),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_495),
.B(n_501),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_582),
.B(n_418),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_485),
.B(n_519),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_485),
.B(n_440),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_497),
.B(n_205),
.C(n_204),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_501),
.B(n_449),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_505),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_461),
.B(n_207),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_523),
.A2(n_594),
.B1(n_574),
.B2(n_470),
.Y(n_769)
);

BUFx8_ASAP7_75t_L g770 ( 
.A(n_468),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_675),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_610),
.B(n_519),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_676),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_675),
.B(n_501),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_698),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_659),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_611),
.A2(n_466),
.B(n_577),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_608),
.B(n_519),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_611),
.A2(n_577),
.B(n_564),
.C(n_567),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_547),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_667),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_601),
.A2(n_466),
.B1(n_520),
.B2(n_513),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_676),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_640),
.B(n_468),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_621),
.A2(n_460),
.B(n_459),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_675),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_620),
.B(n_547),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_604),
.A2(n_460),
.B(n_459),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_657),
.A2(n_587),
.B(n_585),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_700),
.A2(n_568),
.B(n_275),
.C(n_225),
.Y(n_791)
);

NOR2x2_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_266),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_641),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_631),
.A2(n_465),
.B(n_460),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_614),
.B(n_421),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_603),
.A2(n_459),
.B(n_465),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_675),
.B(n_501),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_623),
.B(n_547),
.Y(n_798)
);

O2A1O1Ixp5_ASAP7_75t_L g799 ( 
.A1(n_711),
.A2(n_554),
.B(n_558),
.C(n_580),
.Y(n_799)
);

NOR2x1_ASAP7_75t_L g800 ( 
.A(n_646),
.B(n_554),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_703),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_603),
.A2(n_465),
.B(n_525),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_677),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_700),
.A2(n_711),
.B(n_717),
.C(n_632),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_649),
.B(n_554),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_L g806 ( 
.A(n_613),
.B(n_643),
.C(n_732),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_657),
.A2(n_558),
.B(n_505),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_707),
.A2(n_525),
.B(n_579),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_613),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_664),
.Y(n_810)
);

BUFx4f_ASAP7_75t_L g811 ( 
.A(n_712),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_695),
.A2(n_525),
.B(n_579),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_634),
.A2(n_579),
.B(n_580),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_719),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_702),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_756),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_615),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_680),
.B(n_266),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_717),
.A2(n_769),
.B(n_627),
.C(n_636),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_649),
.B(n_558),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_656),
.A2(n_507),
.B(n_580),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_677),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_656),
.A2(n_507),
.B(n_581),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_634),
.A2(n_726),
.B(n_709),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_682),
.B(n_491),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_617),
.B(n_491),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_682),
.B(n_491),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_745),
.A2(n_503),
.B(n_499),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_626),
.A2(n_304),
.B(n_236),
.C(n_257),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_606),
.B(n_499),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_754),
.A2(n_499),
.B(n_503),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_644),
.A2(n_234),
.B(n_292),
.C(n_299),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_637),
.B(n_499),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_681),
.B(n_266),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_685),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_602),
.B(n_266),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_688),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_712),
.B(n_501),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_639),
.A2(n_499),
.B1(n_503),
.B2(n_565),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_618),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_653),
.A2(n_234),
.B(n_299),
.C(n_292),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_629),
.A2(n_596),
.B(n_581),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_645),
.B(n_503),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_755),
.A2(n_503),
.B(n_514),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_705),
.A2(n_596),
.B(n_572),
.C(n_563),
.Y(n_845)
);

OR2x2_ASAP7_75t_SL g846 ( 
.A(n_624),
.B(n_358),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_759),
.B(n_543),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_712),
.B(n_514),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_678),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_616),
.A2(n_514),
.B(n_565),
.Y(n_850)
);

CKINVDCx10_ASAP7_75t_R g851 ( 
.A(n_683),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_724),
.B(n_514),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_699),
.A2(n_565),
.B1(n_514),
.B2(n_517),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_SL g854 ( 
.A1(n_661),
.A2(n_572),
.B(n_563),
.C(n_561),
.Y(n_854)
);

OAI21xp33_ASAP7_75t_L g855 ( 
.A1(n_732),
.A2(n_760),
.B(n_643),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_622),
.A2(n_565),
.B(n_517),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_622),
.A2(n_517),
.B(n_537),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_652),
.B(n_517),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_724),
.A2(n_561),
.B1(n_550),
.B2(n_546),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_672),
.B(n_537),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_730),
.B(n_543),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_605),
.A2(n_550),
.B1(n_546),
.B2(n_544),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_762),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_770),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_689),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_674),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_619),
.A2(n_544),
.B(n_448),
.C(n_421),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_760),
.B(n_422),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_757),
.A2(n_537),
.B(n_442),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_763),
.A2(n_537),
.B(n_442),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_618),
.B(n_449),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_625),
.B(n_423),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_713),
.B(n_422),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_768),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_625),
.A2(n_435),
.B(n_437),
.C(n_448),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_628),
.B(n_423),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_692),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_628),
.A2(n_435),
.B(n_437),
.C(n_245),
.Y(n_878)
);

OAI21xp33_ASAP7_75t_L g879 ( 
.A1(n_768),
.A2(n_276),
.B(n_211),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_725),
.B(n_765),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_714),
.B(n_254),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_635),
.A2(n_285),
.B1(n_213),
.B2(n_230),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_635),
.B(n_430),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_638),
.A2(n_436),
.B(n_433),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_360),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_651),
.A2(n_663),
.B1(n_654),
.B2(n_666),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_629),
.A2(n_436),
.B(n_433),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_630),
.A2(n_436),
.B(n_433),
.Y(n_888)
);

NOR2x2_ASAP7_75t_L g889 ( 
.A(n_651),
.B(n_430),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_630),
.A2(n_430),
.B(n_443),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_698),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_654),
.B(n_449),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_704),
.B(n_209),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_633),
.A2(n_443),
.B(n_419),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_666),
.B(n_443),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_702),
.Y(n_896)
);

O2A1O1Ixp5_ASAP7_75t_L g897 ( 
.A1(n_633),
.A2(n_360),
.B(n_449),
.C(n_419),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_721),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_722),
.Y(n_899)
);

AOI33xp33_ASAP7_75t_L g900 ( 
.A1(n_718),
.A2(n_252),
.A3(n_256),
.B1(n_268),
.B2(n_269),
.B3(n_272),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_670),
.B(n_443),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_746),
.A2(n_443),
.B(n_419),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_704),
.B(n_274),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_770),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_670),
.B(n_443),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_727),
.B(n_443),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_731),
.A2(n_419),
.B1(n_297),
.B2(n_295),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_747),
.A2(n_419),
.B(n_293),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_764),
.A2(n_419),
.B(n_291),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_673),
.B(n_419),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_741),
.A2(n_284),
.B(n_419),
.C(n_7),
.Y(n_911)
);

NOR2x1_ASAP7_75t_L g912 ( 
.A(n_665),
.B(n_62),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_702),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_761),
.A2(n_151),
.B(n_136),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_660),
.B(n_3),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_728),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_642),
.B(n_647),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_655),
.B(n_4),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_658),
.B(n_7),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_750),
.A2(n_9),
.B(n_15),
.C(n_16),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_684),
.B(n_64),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_662),
.B(n_9),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_702),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_751),
.B(n_15),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_733),
.Y(n_925)
);

NOR2xp67_ASAP7_75t_L g926 ( 
.A(n_706),
.B(n_716),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_691),
.B(n_17),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_686),
.B(n_67),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_761),
.A2(n_66),
.B(n_129),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_668),
.B(n_134),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_696),
.A2(n_122),
.B(n_120),
.Y(n_931)
);

O2A1O1Ixp5_ASAP7_75t_L g932 ( 
.A1(n_691),
.A2(n_113),
.B(n_110),
.C(n_109),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_751),
.A2(n_17),
.B(n_22),
.Y(n_933)
);

INVx11_ASAP7_75t_L g934 ( 
.A(n_770),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_751),
.B(n_22),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_612),
.A2(n_697),
.B(n_671),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_710),
.B(n_23),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_715),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_687),
.A2(n_100),
.B(n_94),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_708),
.Y(n_940)
);

OAI321xp33_ASAP7_75t_L g941 ( 
.A1(n_693),
.A2(n_23),
.A3(n_25),
.B1(n_26),
.B2(n_29),
.C(n_31),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_690),
.B(n_31),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_694),
.B(n_34),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_723),
.B(n_35),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_708),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_736),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_701),
.A2(n_71),
.B(n_88),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_738),
.A2(n_91),
.B(n_84),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_720),
.A2(n_723),
.B(n_735),
.C(n_729),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_729),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_701),
.A2(n_83),
.B(n_80),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_734),
.A2(n_76),
.B(n_74),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_742),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_855),
.B(n_609),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_874),
.B(n_669),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_809),
.B(n_669),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_825),
.A2(n_766),
.B(n_744),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_827),
.A2(n_766),
.B(n_744),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_780),
.A2(n_740),
.B(n_743),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_868),
.B(n_806),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_793),
.B(n_752),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_886),
.A2(n_679),
.B1(n_740),
.B2(n_737),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_840),
.B(n_735),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_886),
.A2(n_811),
.B1(n_926),
.B2(n_852),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_811),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_816),
.B(n_749),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_863),
.B(n_767),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_865),
.B(n_767),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_824),
.A2(n_758),
.B(n_753),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_864),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_877),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_783),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_788),
.A2(n_758),
.B(n_753),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_818),
.B(n_748),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_785),
.A2(n_737),
.B1(n_708),
.B2(n_748),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_810),
.B(n_739),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_834),
.B(n_739),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_923),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_SL g979 ( 
.A(n_941),
.B(n_737),
.Y(n_979)
);

NAND2x1_ASAP7_75t_SL g980 ( 
.A(n_880),
.B(n_39),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_783),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_777),
.A2(n_720),
.B(n_737),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_927),
.A2(n_708),
.B1(n_46),
.B2(n_47),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_804),
.A2(n_40),
.B(n_46),
.C(n_52),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_801),
.B(n_52),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_814),
.B(n_53),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_885),
.B(n_835),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_778),
.B(n_826),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_819),
.A2(n_826),
.B(n_927),
.C(n_879),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_950),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_837),
.A2(n_817),
.B(n_937),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_776),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_772),
.A2(n_789),
.B(n_805),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_820),
.A2(n_843),
.B(n_833),
.Y(n_994)
);

AND2x2_ASAP7_75t_SL g995 ( 
.A(n_937),
.B(n_924),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_836),
.B(n_873),
.Y(n_996)
);

AO32x2_ASAP7_75t_L g997 ( 
.A1(n_782),
.A2(n_853),
.A3(n_839),
.B1(n_882),
.B2(n_933),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_866),
.B(n_861),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_878),
.A2(n_852),
.B(n_875),
.C(n_911),
.Y(n_999)
);

NAND2x1_ASAP7_75t_L g1000 ( 
.A(n_775),
.B(n_771),
.Y(n_1000)
);

CKINVDCx6p67_ASAP7_75t_R g1001 ( 
.A(n_851),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_893),
.A2(n_903),
.B(n_878),
.C(n_943),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_875),
.A2(n_911),
.B(n_935),
.C(n_919),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_849),
.B(n_795),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_781),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_920),
.A2(n_832),
.B(n_841),
.C(n_829),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_849),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_858),
.A2(n_794),
.B(n_796),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_771),
.A2(n_787),
.B1(n_775),
.B2(n_848),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_923),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_889),
.Y(n_1011)
);

BUFx8_ASAP7_75t_SL g1012 ( 
.A(n_904),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_893),
.B(n_903),
.C(n_900),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_846),
.Y(n_1014)
);

OR2x6_ASAP7_75t_SL g1015 ( 
.A(n_792),
.B(n_915),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_786),
.A2(n_936),
.B(n_917),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_942),
.A2(n_943),
.B(n_859),
.C(n_881),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_945),
.B(n_815),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_773),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_945),
.B(n_815),
.Y(n_1020)
);

AOI22x1_ASAP7_75t_L g1021 ( 
.A1(n_850),
.A2(n_857),
.B1(n_856),
.B2(n_887),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_912),
.B(n_898),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_842),
.A2(n_828),
.B(n_802),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_899),
.B(n_916),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_800),
.A2(n_953),
.B1(n_946),
.B2(n_925),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_830),
.A2(n_808),
.B(n_812),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_848),
.A2(n_891),
.B1(n_838),
.B2(n_798),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_784),
.B(n_803),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_944),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_896),
.B(n_940),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_918),
.B(n_922),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_838),
.B(n_871),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_860),
.A2(n_821),
.B(n_799),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_822),
.B(n_938),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_872),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_871),
.B(n_892),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_876),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_907),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_923),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_845),
.A2(n_779),
.B(n_949),
.C(n_906),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_883),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_791),
.A2(n_892),
.B(n_867),
.C(n_930),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_930),
.A2(n_921),
.B(n_928),
.C(n_854),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_923),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_860),
.A2(n_870),
.B(n_869),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_910),
.A2(n_901),
.B(n_895),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_940),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_774),
.A2(n_797),
.B1(n_862),
.B2(n_813),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_774),
.A2(n_797),
.B1(n_896),
.B2(n_905),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_921),
.B(n_928),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_884),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_934),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_940),
.B(n_913),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_952),
.A2(n_932),
.B(n_888),
.C(n_897),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_910),
.A2(n_909),
.B1(n_908),
.B2(n_940),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_807),
.A2(n_913),
.B1(n_844),
.B2(n_831),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_790),
.B(n_823),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_854),
.A2(n_939),
.B(n_931),
.C(n_890),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_914),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_929),
.A2(n_947),
.B(n_951),
.C(n_894),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_902),
.Y(n_1061)
);

BUFx8_ASAP7_75t_L g1062 ( 
.A(n_948),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_874),
.B(n_855),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_863),
.B(n_795),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_809),
.B(n_608),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_904),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_825),
.A2(n_601),
.B(n_603),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_865),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_811),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_783),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_783),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_809),
.B(n_608),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_809),
.B(n_426),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_809),
.B(n_874),
.Y(n_1074)
);

CKINVDCx8_ASAP7_75t_R g1075 ( 
.A(n_851),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_809),
.B(n_874),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_809),
.B(n_874),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_783),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_855),
.A2(n_804),
.B(n_878),
.C(n_809),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_874),
.B(n_855),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_809),
.B(n_608),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_855),
.A2(n_806),
.B(n_804),
.C(n_819),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_855),
.A2(n_806),
.B(n_804),
.C(n_819),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_874),
.B(n_855),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_783),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_855),
.A2(n_806),
.B1(n_608),
.B2(n_601),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_863),
.B(n_795),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_809),
.B(n_608),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_825),
.A2(n_601),
.B(n_603),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_855),
.A2(n_806),
.B1(n_608),
.B2(n_601),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_855),
.A2(n_806),
.B1(n_608),
.B2(n_601),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_855),
.A2(n_806),
.B1(n_724),
.B2(n_926),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_809),
.B(n_608),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_989),
.A2(n_1083),
.B(n_1082),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1081),
.B(n_1088),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_1016),
.A2(n_958),
.B(n_957),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1017),
.A2(n_1002),
.B(n_1086),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1001),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1079),
.A2(n_1092),
.B(n_1050),
.C(n_1013),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_995),
.A2(n_991),
.B1(n_996),
.B2(n_960),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_988),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1067),
.A2(n_1089),
.B(n_958),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1093),
.B(n_1073),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_957),
.A2(n_994),
.B(n_993),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1064),
.B(n_1087),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1063),
.A2(n_1084),
.B1(n_1080),
.B2(n_1077),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1031),
.A2(n_1079),
.B(n_1038),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1010),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_964),
.A2(n_1040),
.B(n_1043),
.Y(n_1111)
);

BUFx2_ASAP7_75t_SL g1112 ( 
.A(n_1044),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_971),
.Y(n_1113)
);

OA21x2_ASAP7_75t_L g1114 ( 
.A1(n_993),
.A2(n_1033),
.B(n_994),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1029),
.B(n_977),
.Y(n_1115)
);

BUFx2_ASAP7_75t_R g1116 ( 
.A(n_1075),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1004),
.B(n_987),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1074),
.B(n_1076),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_972),
.Y(n_1120)
);

BUFx8_ASAP7_75t_L g1121 ( 
.A(n_1011),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1064),
.B(n_1087),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_974),
.B(n_1024),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_954),
.A2(n_983),
.B1(n_1014),
.B2(n_1022),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1008),
.A2(n_1057),
.B(n_1033),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1032),
.A2(n_1036),
.B1(n_956),
.B2(n_976),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_967),
.B(n_1037),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_981),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1078),
.B(n_1085),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1070),
.B(n_966),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_L g1131 ( 
.A(n_1006),
.B(n_984),
.C(n_1025),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1054),
.A2(n_1008),
.A3(n_1048),
.B(n_1045),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1043),
.A2(n_999),
.B(n_1003),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_965),
.B(n_1069),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_965),
.B(n_1069),
.Y(n_1135)
);

CKINVDCx11_ASAP7_75t_R g1136 ( 
.A(n_970),
.Y(n_1136)
);

NOR4xp25_ASAP7_75t_L g1137 ( 
.A(n_984),
.B(n_999),
.C(n_1003),
.D(n_1042),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1056),
.A2(n_959),
.B(n_1058),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_973),
.A2(n_1045),
.B(n_1021),
.Y(n_1139)
);

OAI22x1_ASAP7_75t_L g1140 ( 
.A1(n_992),
.A2(n_1005),
.B1(n_998),
.B2(n_1007),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_SL g1141 ( 
.A1(n_1042),
.A2(n_1009),
.B(n_1027),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1041),
.B(n_1068),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_965),
.B(n_1069),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1059),
.A2(n_975),
.B1(n_955),
.B2(n_963),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_959),
.A2(n_1058),
.B(n_982),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_985),
.A2(n_986),
.B(n_1000),
.C(n_1028),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1015),
.B(n_1071),
.Y(n_1147)
);

AO21x1_ASAP7_75t_L g1148 ( 
.A1(n_1049),
.A2(n_982),
.B(n_1046),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_961),
.B(n_968),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_1034),
.A2(n_962),
.B(n_990),
.C(n_1035),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1061),
.A2(n_1060),
.B(n_1046),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1055),
.A2(n_1051),
.B(n_1019),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1053),
.A2(n_1020),
.B(n_1018),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_979),
.A2(n_1020),
.B(n_1018),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1010),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1062),
.A2(n_997),
.A3(n_980),
.B(n_1030),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_997),
.A2(n_1010),
.B(n_1039),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1039),
.A2(n_1047),
.B(n_997),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1047),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1012),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1066),
.A2(n_1092),
.B1(n_855),
.B2(n_806),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1052),
.A2(n_969),
.B(n_1023),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_965),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1168)
);

NAND2x1_ASAP7_75t_L g1169 ( 
.A(n_978),
.B(n_896),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1065),
.B(n_452),
.Y(n_1170)
);

AOI31xp67_ASAP7_75t_L g1171 ( 
.A1(n_988),
.A2(n_892),
.A3(n_871),
.B(n_825),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_SL g1174 ( 
.A1(n_999),
.A2(n_819),
.B(n_1079),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1082),
.A2(n_1083),
.A3(n_989),
.B(n_1016),
.Y(n_1175)
);

CKINVDCx11_ASAP7_75t_R g1176 ( 
.A(n_1075),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1082),
.A2(n_1083),
.A3(n_989),
.B(n_1016),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1082),
.A2(n_1083),
.A3(n_989),
.B(n_1016),
.Y(n_1178)
);

AOI221x1_ASAP7_75t_L g1179 ( 
.A1(n_989),
.A2(n_855),
.B1(n_1083),
.B2(n_1082),
.C(n_1017),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1092),
.B(n_806),
.C(n_855),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1064),
.B(n_553),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_989),
.A2(n_806),
.B(n_855),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_989),
.A2(n_806),
.B(n_855),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_972),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_1074),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_989),
.A2(n_1083),
.B(n_1082),
.C(n_1002),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_965),
.B(n_1069),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_971),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1079),
.A2(n_855),
.B(n_806),
.C(n_1002),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_SL g1191 ( 
.A1(n_989),
.A2(n_1083),
.B(n_1082),
.C(n_1002),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1092),
.A2(n_855),
.B1(n_806),
.B2(n_608),
.Y(n_1192)
);

NAND2xp33_ASAP7_75t_SL g1193 ( 
.A(n_1044),
.B(n_669),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1082),
.A2(n_1083),
.A3(n_989),
.B(n_1016),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1195)
);

AO32x2_ASAP7_75t_L g1196 ( 
.A1(n_1086),
.A2(n_1091),
.A3(n_1090),
.B1(n_964),
.B2(n_1048),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_SL g1197 ( 
.A1(n_995),
.A2(n_874),
.B1(n_937),
.B2(n_477),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_995),
.A2(n_855),
.B1(n_806),
.B2(n_724),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_SL g1200 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1090),
.C(n_717),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_954),
.A2(n_553),
.B1(n_806),
.B2(n_426),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_965),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1079),
.A2(n_855),
.B(n_806),
.C(n_1002),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1002),
.A2(n_855),
.B(n_874),
.C(n_1017),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_989),
.A2(n_1083),
.B(n_1082),
.C(n_1002),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1211)
);

NOR2x1_ASAP7_75t_R g1212 ( 
.A(n_1052),
.B(n_589),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1078),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1079),
.A2(n_855),
.B(n_806),
.C(n_1002),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_965),
.B(n_1069),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_1086),
.A2(n_1091),
.A3(n_1090),
.B1(n_964),
.B2(n_1048),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1082),
.A2(n_1083),
.A3(n_989),
.B(n_1016),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_969),
.A2(n_1023),
.B(n_1026),
.Y(n_1219)
);

AOI221xp5_ASAP7_75t_SL g1220 ( 
.A1(n_991),
.A2(n_617),
.B1(n_632),
.B2(n_650),
.C(n_855),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1092),
.A2(n_855),
.B1(n_806),
.B2(n_608),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1016),
.A2(n_1089),
.B(n_1067),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_971),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_972),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_965),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1213),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1176),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1109),
.A2(n_1095),
.B1(n_1180),
.B2(n_1183),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1129),
.Y(n_1233)
);

BUFx4_ASAP7_75t_R g1234 ( 
.A(n_1185),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1136),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1197),
.A2(n_1133),
.B1(n_1111),
.B2(n_1098),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1113),
.Y(n_1237)
);

INVx6_ASAP7_75t_L g1238 ( 
.A(n_1164),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1164),
.Y(n_1239)
);

INVx6_ASAP7_75t_L g1240 ( 
.A(n_1134),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_1112),
.Y(n_1241)
);

BUFx8_ASAP7_75t_L g1242 ( 
.A(n_1160),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1180),
.A2(n_1182),
.B1(n_1198),
.B2(n_1202),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1110),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1120),
.Y(n_1245)
);

BUFx4_ASAP7_75t_SL g1246 ( 
.A(n_1099),
.Y(n_1246)
);

CKINVDCx8_ASAP7_75t_R g1247 ( 
.A(n_1160),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1116),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1134),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1157),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1198),
.A2(n_1192),
.B1(n_1224),
.B2(n_1131),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1135),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1110),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1160),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1175),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1185),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1131),
.A2(n_1161),
.B1(n_1103),
.B2(n_1174),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1119),
.A2(n_1197),
.B1(n_1124),
.B2(n_1108),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1189),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1226),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1121),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1121),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1135),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1102),
.A2(n_1124),
.B1(n_1126),
.B2(n_1108),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1142),
.Y(n_1265)
);

NAND2x1p5_ASAP7_75t_L g1266 ( 
.A(n_1205),
.B(n_1228),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1102),
.A2(n_1181),
.B1(n_1141),
.B2(n_1123),
.Y(n_1267)
);

BUFx8_ASAP7_75t_SL g1268 ( 
.A(n_1147),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1105),
.A2(n_1229),
.B1(n_1096),
.B2(n_1223),
.Y(n_1269)
);

INVx3_ASAP7_75t_SL g1270 ( 
.A(n_1143),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1127),
.Y(n_1271)
);

CKINVDCx8_ASAP7_75t_R g1272 ( 
.A(n_1143),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1188),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1220),
.A2(n_1107),
.B1(n_1193),
.B2(n_1122),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_1188),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1215),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1195),
.A2(n_1221),
.B1(n_1211),
.B2(n_1204),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1117),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1215),
.Y(n_1279)
);

BUFx8_ASAP7_75t_L g1280 ( 
.A(n_1094),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1187),
.A2(n_1208),
.B1(n_1191),
.B2(n_1179),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1155),
.Y(n_1283)
);

CKINVDCx11_ASAP7_75t_R g1284 ( 
.A(n_1212),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1201),
.A2(n_1115),
.B1(n_1149),
.B2(n_1170),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1144),
.A2(n_1140),
.B1(n_1138),
.B2(n_1148),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1227),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1190),
.A2(n_1206),
.B1(n_1214),
.B2(n_1100),
.Y(n_1289)
);

CKINVDCx11_ASAP7_75t_R g1290 ( 
.A(n_1212),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1228),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1128),
.A2(n_1184),
.B1(n_1130),
.B2(n_1207),
.Y(n_1292)
);

INVx6_ASAP7_75t_L g1293 ( 
.A(n_1153),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_1152),
.B2(n_1145),
.Y(n_1294)
);

BUFx4f_ASAP7_75t_L g1295 ( 
.A(n_1114),
.Y(n_1295)
);

BUFx8_ASAP7_75t_L g1296 ( 
.A(n_1196),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1137),
.A2(n_1196),
.B1(n_1216),
.B2(n_1114),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1125),
.A2(n_1097),
.B1(n_1104),
.B2(n_1101),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1169),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1146),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1156),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1163),
.A2(n_1167),
.B1(n_1225),
.B2(n_1222),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1156),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1165),
.A2(n_1166),
.B1(n_1172),
.B2(n_1203),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1156),
.B(n_1162),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1137),
.A2(n_1216),
.B1(n_1196),
.B2(n_1199),
.Y(n_1307)
);

AOI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1151),
.A2(n_1186),
.B(n_1106),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1178),
.B(n_1217),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1194),
.Y(n_1310)
);

CKINVDCx16_ASAP7_75t_R g1311 ( 
.A(n_1171),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1194),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1217),
.A2(n_1200),
.B1(n_1150),
.B2(n_1132),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1132),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1139),
.A2(n_1118),
.B1(n_1168),
.B2(n_1173),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1209),
.A2(n_1210),
.B1(n_1218),
.B2(n_1219),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1119),
.A2(n_995),
.B1(n_1197),
.B2(n_1124),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1176),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1109),
.A2(n_995),
.B1(n_855),
.B2(n_806),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1176),
.Y(n_1320)
);

BUFx8_ASAP7_75t_SL g1321 ( 
.A(n_1099),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1197),
.A2(n_995),
.B1(n_426),
.B2(n_1095),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1129),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1119),
.A2(n_995),
.B1(n_1197),
.B2(n_1124),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1113),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1176),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1176),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1129),
.Y(n_1328)
);

BUFx8_ASAP7_75t_L g1329 ( 
.A(n_1160),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1213),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1176),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1176),
.Y(n_1332)
);

CKINVDCx11_ASAP7_75t_R g1333 ( 
.A(n_1176),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_1176),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1095),
.A2(n_1191),
.B(n_1187),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1190),
.A2(n_806),
.B(n_855),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1176),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1113),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1113),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1198),
.A2(n_855),
.B1(n_314),
.B2(n_364),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1096),
.B(n_1195),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1278),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1308),
.A2(n_1313),
.B(n_1307),
.Y(n_1343)
);

NOR2x1_ASAP7_75t_R g1344 ( 
.A(n_1326),
.B(n_1333),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1296),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1315),
.A2(n_1316),
.B(n_1299),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1287),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1321),
.Y(n_1348)
);

AOI21xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1258),
.A2(n_1324),
.B(n_1317),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1310),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1312),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1246),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1296),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1309),
.B(n_1236),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1297),
.B(n_1255),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1232),
.B(n_1236),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1250),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1302),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1287),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1257),
.B(n_1232),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1250),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1245),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1293),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1233),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1269),
.B(n_1277),
.Y(n_1365)
);

AOI222xp33_ASAP7_75t_L g1366 ( 
.A1(n_1289),
.A2(n_1264),
.B1(n_1319),
.B2(n_1336),
.C1(n_1251),
.C2(n_1243),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1280),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1314),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1295),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1295),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1293),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1323),
.B(n_1328),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1306),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1311),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1237),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1293),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1230),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1257),
.B(n_1251),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1341),
.B(n_1340),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1313),
.A2(n_1307),
.B(n_1294),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1260),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1325),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1338),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1280),
.A2(n_1335),
.B1(n_1301),
.B2(n_1322),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1339),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1241),
.B(n_1285),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1303),
.A2(n_1305),
.B(n_1299),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1259),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1298),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1298),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1322),
.A2(n_1319),
.B1(n_1264),
.B2(n_1243),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1286),
.B(n_1267),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1269),
.B(n_1285),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1305),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1254),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1286),
.A2(n_1267),
.B(n_1292),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_R g1397 ( 
.A(n_1248),
.B(n_1337),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1271),
.B(n_1265),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1281),
.B(n_1288),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1281),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1330),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1304),
.Y(n_1402)
);

INVxp33_ASAP7_75t_L g1403 ( 
.A(n_1256),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1274),
.A2(n_1266),
.B(n_1252),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1300),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1234),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1291),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1262),
.A2(n_1273),
.B1(n_1276),
.B2(n_1283),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1365),
.B(n_1276),
.Y(n_1409)
);

AOI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1349),
.A2(n_1279),
.B1(n_1275),
.B2(n_1282),
.C(n_1270),
.Y(n_1410)
);

OAI211xp5_ASAP7_75t_L g1411 ( 
.A1(n_1366),
.A2(n_1272),
.B(n_1247),
.C(n_1283),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1366),
.A2(n_1349),
.B(n_1379),
.Y(n_1412)
);

AND2x2_ASAP7_75t_SL g1413 ( 
.A(n_1387),
.B(n_1234),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1391),
.A2(n_1384),
.B1(n_1356),
.B2(n_1406),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1356),
.A2(n_1261),
.B(n_1332),
.C(n_1318),
.Y(n_1415)
);

AO21x1_ASAP7_75t_L g1416 ( 
.A1(n_1386),
.A2(n_1282),
.B(n_1253),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1375),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1396),
.A2(n_1393),
.B(n_1365),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1346),
.A2(n_1244),
.B(n_1263),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1357),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1378),
.A2(n_1240),
.B1(n_1263),
.B2(n_1249),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1357),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1393),
.A2(n_1378),
.B(n_1360),
.C(n_1392),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1346),
.A2(n_1249),
.B(n_1238),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1396),
.A2(n_1268),
.B(n_1290),
.C(n_1284),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1369),
.B(n_1334),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1345),
.B(n_1353),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1246),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1342),
.B(n_1329),
.Y(n_1429)
);

AO32x2_ASAP7_75t_L g1430 ( 
.A1(n_1347),
.A2(n_1239),
.A3(n_1329),
.B1(n_1242),
.B2(n_1235),
.Y(n_1430)
);

AO32x2_ASAP7_75t_L g1431 ( 
.A1(n_1347),
.A2(n_1239),
.A3(n_1242),
.B1(n_1231),
.B2(n_1320),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1360),
.A2(n_1327),
.B1(n_1331),
.B2(n_1392),
.C(n_1354),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1350),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1406),
.A2(n_1408),
.B1(n_1402),
.B2(n_1401),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1400),
.A2(n_1406),
.B1(n_1364),
.B2(n_1372),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1361),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1377),
.B(n_1406),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1404),
.A2(n_1394),
.B(n_1363),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_SL g1440 ( 
.A(n_1359),
.B(n_1355),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1362),
.B(n_1398),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1388),
.B(n_1407),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1404),
.B(n_1363),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1355),
.B(n_1394),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1446)
);

AO32x2_ASAP7_75t_L g1447 ( 
.A1(n_1363),
.A2(n_1371),
.A3(n_1390),
.B1(n_1389),
.B2(n_1380),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1344),
.A2(n_1367),
.B(n_1387),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1405),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1447),
.B(n_1424),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1433),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1447),
.B(n_1380),
.Y(n_1454)
);

OR2x6_ASAP7_75t_SL g1455 ( 
.A(n_1414),
.B(n_1445),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1436),
.B(n_1373),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1447),
.B(n_1343),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1419),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1447),
.B(n_1343),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1420),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1436),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1420),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_L g1463 ( 
.A(n_1412),
.B(n_1400),
.C(n_1399),
.Y(n_1463)
);

NOR2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1428),
.B(n_1367),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1417),
.Y(n_1465)
);

OAI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1423),
.A2(n_1367),
.B1(n_1371),
.B2(n_1405),
.C(n_1376),
.Y(n_1466)
);

AND2x2_ASAP7_75t_SL g1467 ( 
.A(n_1413),
.B(n_1358),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1451),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1418),
.B(n_1368),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1446),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1449),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1351),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1437),
.B(n_1368),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1457),
.A2(n_1444),
.B(n_1439),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1462),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1468),
.B(n_1422),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1462),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1467),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1466),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1453),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1468),
.B(n_1469),
.Y(n_1481)
);

OAI321xp33_ASAP7_75t_L g1482 ( 
.A1(n_1463),
.A2(n_1466),
.A3(n_1411),
.B1(n_1423),
.B2(n_1454),
.C(n_1457),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1461),
.B(n_1440),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1473),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1465),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1461),
.B(n_1413),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1467),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1467),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1472),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1463),
.A2(n_1435),
.B1(n_1395),
.B2(n_1434),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1456),
.B(n_1427),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1470),
.B(n_1422),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1467),
.B(n_1425),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1460),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1466),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1458),
.B(n_1443),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1463),
.A2(n_1432),
.B1(n_1444),
.B2(n_1435),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1467),
.A2(n_1425),
.B(n_1448),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1468),
.B(n_1469),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1455),
.A2(n_1409),
.B1(n_1421),
.B2(n_1410),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1489),
.B(n_1452),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1475),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1475),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1476),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1478),
.B(n_1458),
.Y(n_1506)
);

NAND4xp25_ASAP7_75t_L g1507 ( 
.A(n_1497),
.B(n_1415),
.C(n_1457),
.D(n_1459),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1477),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1458),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1478),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1498),
.B(n_1426),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

BUFx2_ASAP7_75t_SL g1513 ( 
.A(n_1478),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1498),
.B(n_1426),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1479),
.Y(n_1515)
);

NOR2x1_ASAP7_75t_L g1516 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1496),
.B(n_1454),
.Y(n_1518)
);

NOR2x1_ASAP7_75t_L g1519 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1477),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1458),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1480),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1492),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1485),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1496),
.B(n_1454),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1499),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1484),
.B(n_1479),
.Y(n_1529)
);

INVxp67_ASAP7_75t_SL g1530 ( 
.A(n_1495),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1485),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1484),
.B(n_1471),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1480),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1529),
.B(n_1474),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

AOI32xp33_ASAP7_75t_L g1536 ( 
.A1(n_1515),
.A2(n_1482),
.A3(n_1488),
.B1(n_1493),
.B2(n_1459),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1515),
.B(n_1495),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1512),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1521),
.B(n_1524),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1502),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1507),
.A2(n_1482),
.B(n_1415),
.C(n_1459),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1502),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1520),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1523),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1503),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1507),
.B(n_1474),
.Y(n_1550)
);

AOI21xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1511),
.A2(n_1490),
.B(n_1403),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1508),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1503),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1521),
.B(n_1474),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1525),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1514),
.A2(n_1455),
.B1(n_1490),
.B2(n_1488),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1510),
.B(n_1344),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1491),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1517),
.B(n_1483),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1528),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1504),
.B(n_1481),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1528),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1532),
.B(n_1491),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1517),
.B(n_1483),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1532),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1523),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1522),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1504),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1523),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1510),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1538),
.B(n_1542),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1505),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1566),
.B(n_1505),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1535),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1555),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1552),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1572),
.B(n_1519),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1564),
.B(n_1501),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1559),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1572),
.B(n_1513),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1564),
.B(n_1527),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1559),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1572),
.B(n_1513),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1537),
.B(n_1506),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1562),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1569),
.B(n_1501),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1569),
.B(n_1527),
.Y(n_1594)
);

NOR2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1550),
.B(n_1395),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1537),
.B(n_1560),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1506),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1541),
.B(n_1508),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1562),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1535),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1539),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1563),
.Y(n_1602)
);

NAND4xp75_ASAP7_75t_L g1603 ( 
.A(n_1557),
.B(n_1457),
.C(n_1459),
.D(n_1416),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1561),
.B(n_1568),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1575),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_L g1606 ( 
.A(n_1545),
.B(n_1405),
.C(n_1500),
.Y(n_1606)
);

AOI221x1_ASAP7_75t_L g1607 ( 
.A1(n_1551),
.A2(n_1500),
.B1(n_1405),
.B2(n_1450),
.C(n_1506),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1506),
.Y(n_1608)
);

INVxp67_ASAP7_75t_SL g1609 ( 
.A(n_1534),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1536),
.B(n_1509),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1604),
.B(n_1571),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1606),
.A2(n_1556),
.B(n_1534),
.Y(n_1612)
);

OAI322xp33_ASAP7_75t_L g1613 ( 
.A1(n_1605),
.A2(n_1554),
.A3(n_1573),
.B1(n_1549),
.B2(n_1544),
.C1(n_1546),
.C2(n_1553),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1604),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1606),
.A2(n_1607),
.B(n_1610),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1582),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1582),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1587),
.Y(n_1618)
);

NAND2x1_ASAP7_75t_SL g1619 ( 
.A(n_1584),
.B(n_1571),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1576),
.A2(n_1571),
.B1(n_1573),
.B2(n_1546),
.C(n_1544),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1587),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1603),
.A2(n_1455),
.B1(n_1567),
.B2(n_1509),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1577),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1395),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1577),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1596),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1603),
.A2(n_1455),
.B1(n_1509),
.B2(n_1522),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1590),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1590),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1576),
.B(n_1352),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1607),
.B(n_1596),
.C(n_1578),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1578),
.B(n_1549),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1581),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1558),
.Y(n_1634)
);

OAI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1584),
.A2(n_1543),
.B1(n_1565),
.B2(n_1563),
.C(n_1441),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1619),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1616),
.Y(n_1637)
);

NOR2xp67_ASAP7_75t_SL g1638 ( 
.A(n_1615),
.B(n_1348),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1619),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1617),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1623),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1625),
.Y(n_1642)
);

AOI311xp33_ASAP7_75t_L g1643 ( 
.A1(n_1622),
.A2(n_1609),
.A3(n_1599),
.B(n_1589),
.C(n_1602),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1633),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1618),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1612),
.A2(n_1598),
.B(n_1579),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1618),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1624),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1627),
.A2(n_1595),
.B(n_1609),
.C(n_1598),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1626),
.B(n_1591),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1628),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1621),
.B(n_1608),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1621),
.B(n_1628),
.Y(n_1653)
);

AOI22x1_ASAP7_75t_L g1654 ( 
.A1(n_1629),
.A2(n_1595),
.B1(n_1614),
.B2(n_1631),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1624),
.B(n_1608),
.C(n_1597),
.D(n_1583),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1638),
.A2(n_1629),
.B1(n_1597),
.B2(n_1634),
.Y(n_1656)
);

OAI31xp33_ASAP7_75t_L g1657 ( 
.A1(n_1639),
.A2(n_1620),
.A3(n_1635),
.B(n_1630),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1648),
.B(n_1630),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1655),
.B(n_1632),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1654),
.A2(n_1579),
.B1(n_1583),
.B2(n_1611),
.C(n_1593),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1637),
.Y(n_1661)
);

AO22x2_ASAP7_75t_L g1662 ( 
.A1(n_1637),
.A2(n_1599),
.B1(n_1589),
.B2(n_1602),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1649),
.B(n_1613),
.C(n_1611),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1647),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1657),
.B(n_1643),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1664),
.B(n_1651),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1662),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1662),
.A2(n_1646),
.B(n_1654),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1659),
.A2(n_1636),
.B1(n_1652),
.B2(n_1653),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1658),
.B(n_1640),
.Y(n_1671)
);

NOR3x1_ASAP7_75t_L g1672 ( 
.A(n_1663),
.B(n_1642),
.C(n_1641),
.Y(n_1672)
);

AND3x1_ASAP7_75t_L g1673 ( 
.A(n_1656),
.B(n_1636),
.C(n_1644),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_L g1674 ( 
.A(n_1661),
.B(n_1638),
.C(n_1586),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1669),
.A2(n_1660),
.B1(n_1665),
.B2(n_1592),
.C(n_1586),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1666),
.A2(n_1667),
.B1(n_1673),
.B2(n_1674),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_L g1677 ( 
.A1(n_1670),
.A2(n_1593),
.B(n_1585),
.Y(n_1677)
);

AOI31xp33_ASAP7_75t_L g1678 ( 
.A1(n_1668),
.A2(n_1397),
.A3(n_1594),
.B(n_1588),
.Y(n_1678)
);

NAND5xp2_ASAP7_75t_L g1679 ( 
.A(n_1671),
.B(n_1581),
.C(n_1592),
.D(n_1585),
.E(n_1438),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1678),
.Y(n_1680)
);

AOI221x1_ASAP7_75t_L g1681 ( 
.A1(n_1677),
.A2(n_1672),
.B1(n_1601),
.B2(n_1600),
.C(n_1580),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_R g1682 ( 
.A(n_1676),
.B(n_1429),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1675),
.A2(n_1601),
.B1(n_1600),
.B2(n_1580),
.C(n_1588),
.Y(n_1683)
);

OAI211xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1679),
.A2(n_1601),
.B(n_1600),
.C(n_1580),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1678),
.A2(n_1594),
.B(n_1543),
.C(n_1522),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1680),
.B(n_1565),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1681),
.B(n_1509),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1682),
.Y(n_1688)
);

XOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1685),
.B(n_1426),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1684),
.A2(n_1522),
.B1(n_1570),
.B2(n_1548),
.Y(n_1690)
);

OAI22x1_ASAP7_75t_L g1691 ( 
.A1(n_1688),
.A2(n_1683),
.B1(n_1522),
.B2(n_1570),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1686),
.B(n_1539),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1689),
.A2(n_1574),
.B1(n_1548),
.B2(n_1540),
.Y(n_1693)
);

XNOR2xp5_ASAP7_75t_L g1694 ( 
.A(n_1691),
.B(n_1687),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1690),
.B1(n_1693),
.B2(n_1692),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1695),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1574),
.C(n_1540),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_L g1698 ( 
.A(n_1696),
.B(n_1533),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1697),
.A2(n_1431),
.B1(n_1430),
.B2(n_1438),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1698),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1699),
.A2(n_1526),
.B(n_1518),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1700),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1701),
.B(n_1494),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1703),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1533),
.B1(n_1494),
.B2(n_1518),
.C(n_1526),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1705),
.A2(n_1431),
.B(n_1430),
.C(n_1533),
.Y(n_1706)
);


endmodule