module fake_jpeg_18149_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_46),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_58),
.B1(n_41),
.B2(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_19),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_60),
.C(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_34),
.B1(n_25),
.B2(n_23),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_64),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_34),
.C(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_0),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_34),
.B1(n_40),
.B2(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_36),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_33),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_27),
.B(n_28),
.C(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_76),
.A2(n_78),
.B1(n_85),
.B2(n_88),
.Y(n_143)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_37),
.B1(n_45),
.B2(n_21),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_87),
.B1(n_90),
.B2(n_94),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_83),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_37),
.B1(n_45),
.B2(n_21),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_23),
.B1(n_26),
.B2(n_35),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_26),
.B1(n_35),
.B2(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_97),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_92),
.B(n_100),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_45),
.B1(n_37),
.B2(n_25),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_35),
.B1(n_42),
.B2(n_18),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_107),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_108),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_106),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_109),
.Y(n_141)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_47),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_63),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_30),
.B1(n_27),
.B2(n_22),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_8),
.B1(n_14),
.B2(n_3),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_0),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_65),
.B1(n_57),
.B2(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_124),
.B1(n_138),
.B2(n_140),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_46),
.B(n_1),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_118),
.B(n_120),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_29),
.B1(n_19),
.B2(n_22),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_29),
.B1(n_19),
.B2(n_22),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_29),
.B1(n_22),
.B2(n_16),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_91),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_22),
.B1(n_16),
.B2(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_86),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_139),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_0),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_12),
.B(n_13),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_9),
.B1(n_14),
.B2(n_3),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_137),
.B1(n_10),
.B2(n_12),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_1),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_2),
.B1(n_7),
.B2(n_10),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_79),
.B1(n_106),
.B2(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_80),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_111),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_151),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_178),
.B1(n_179),
.B2(n_132),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_93),
.C(n_108),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_93),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_160),
.B(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_109),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_163),
.B(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_75),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_77),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_177),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_98),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_98),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_138),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_10),
.B(n_12),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_120),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_115),
.B1(n_116),
.B2(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_176),
.B1(n_124),
.B2(n_142),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_140),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_115),
.A2(n_119),
.B1(n_145),
.B2(n_137),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_73),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_73),
.B1(n_13),
.B2(n_15),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_122),
.A2(n_133),
.B1(n_125),
.B2(n_114),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_181),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_144),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_190),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_195),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_204),
.B1(n_209),
.B2(n_181),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_121),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_121),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_198),
.B(n_155),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_118),
.B1(n_120),
.B2(n_132),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_153),
.B1(n_152),
.B2(n_161),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_120),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_118),
.B1(n_117),
.B2(n_123),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_155),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_117),
.B1(n_13),
.B2(n_15),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_172),
.B(n_175),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_162),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_222),
.B(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_226),
.B1(n_227),
.B2(n_193),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_177),
.C(n_149),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_220),
.C(n_223),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_214),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_223),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_191),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_225),
.B1(n_198),
.B2(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_150),
.C(n_164),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_229),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_152),
.B(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_150),
.C(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_224),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_165),
.B(n_154),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_154),
.B1(n_192),
.B2(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_204),
.B1(n_202),
.B2(n_206),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_201),
.B(n_199),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_199),
.B(n_209),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_185),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_234),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_246),
.B1(n_252),
.B2(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_190),
.C(n_203),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_242),
.C(n_243),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_185),
.C(n_180),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_217),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_205),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_215),
.C(n_218),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_246),
.C(n_252),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_191),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_196),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_254),
.B(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_230),
.B1(n_214),
.B2(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_216),
.B1(n_225),
.B2(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_231),
.B(n_224),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_270),
.B(n_253),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_207),
.B1(n_239),
.B2(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_258),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_275),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_282),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_258),
.C(n_268),
.Y(n_285)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_289),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_265),
.C(n_267),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_253),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_262),
.B1(n_274),
.B2(n_283),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_263),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_283),
.Y(n_302)
);

AOI31xp67_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_287),
.A3(n_278),
.B(n_292),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_304),
.B(n_299),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_293),
.C(n_286),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_295),
.B(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_305),
.B(n_281),
.C(n_293),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_309),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_264),
.Y(n_313)
);


endmodule