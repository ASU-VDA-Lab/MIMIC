module fake_netlist_1_156_n_1232 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1232, n_1233);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1232;
output n_1233;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_1159;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_677;
wire n_756;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_536;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1195;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g326 ( .A(n_57), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_107), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_178), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_80), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_29), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_67), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_78), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_12), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_98), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_272), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_300), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_316), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_237), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_81), .Y(n_339) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_150), .Y(n_340) );
CKINVDCx14_ASAP7_75t_R g341 ( .A(n_164), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_33), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_0), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_123), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_313), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_24), .B(n_251), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_230), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_86), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_17), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_199), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_288), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_2), .Y(n_354) );
CKINVDCx14_ASAP7_75t_R g355 ( .A(n_122), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_179), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_312), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_259), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_32), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_80), .B(n_181), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_276), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_98), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_256), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_266), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_242), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_0), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_138), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_17), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_115), .Y(n_370) );
INVxp33_ASAP7_75t_L g371 ( .A(n_13), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_271), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_129), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_92), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_119), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_45), .Y(n_377) );
INVxp33_ASAP7_75t_SL g378 ( .A(n_70), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_183), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_166), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_167), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_307), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_264), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_297), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_169), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_320), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_283), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_111), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_130), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_137), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_68), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_114), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_285), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_258), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_103), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_318), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_279), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_311), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_155), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_195), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_184), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_16), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_25), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_177), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_27), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_111), .Y(n_407) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_189), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_92), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_244), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_239), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_262), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_205), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_149), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_59), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_20), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_234), .Y(n_417) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_173), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_116), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_107), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_115), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_144), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_231), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_193), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_41), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_61), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_249), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_203), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_42), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_156), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_296), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_278), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_267), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_51), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_196), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_188), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_25), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_141), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_51), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_229), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_72), .Y(n_441) );
INVxp33_ASAP7_75t_SL g442 ( .A(n_65), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_147), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_54), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_250), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_163), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_133), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_37), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_10), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_15), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_30), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_84), .Y(n_452) );
NOR2xp67_ASAP7_75t_L g453 ( .A(n_268), .B(n_53), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_182), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_93), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_26), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_299), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_95), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_99), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_226), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_135), .B(n_11), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_131), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_54), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_134), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_41), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_145), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_227), .Y(n_467) );
BUFx10_ASAP7_75t_L g468 ( .A(n_281), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_286), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_165), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_200), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_274), .Y(n_472) );
INVxp33_ASAP7_75t_SL g473 ( .A(n_43), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_32), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_260), .Y(n_475) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_254), .B(n_15), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_255), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_303), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_67), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_247), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_222), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_378), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_373), .B(n_1), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_344), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_399), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_346), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_363), .B(n_4), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_371), .B(n_5), .Y(n_488) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_388), .A2(n_121), .B(n_120), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_339), .B(n_6), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_354), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_371), .B(n_6), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_399), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_399), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_354), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_399), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_366), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_328), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_429), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_341), .B(n_7), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_370), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_352), .B(n_7), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_388), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_378), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_391), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_339), .B(n_8), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_341), .B(n_9), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_391), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_362), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_328), .Y(n_510) );
BUFx2_ASAP7_75t_L g511 ( .A(n_362), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_370), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_410), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_442), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_442), .A2(n_19), .B1(n_16), .B2(n_18), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_410), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_396), .B(n_18), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_374), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_462), .B(n_19), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_355), .B(n_21), .Y(n_520) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_413), .A2(n_125), .B(n_124), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_497), .B(n_383), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_503), .Y(n_524) );
OR2x6_ASAP7_75t_L g525 ( .A(n_484), .B(n_441), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_496), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_509), .B(n_469), .Y(n_527) );
AND2x6_ASAP7_75t_L g528 ( .A(n_490), .B(n_374), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_503), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_486), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_509), .B(n_475), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_496), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_496), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_484), .B(n_441), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_496), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_505), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_499), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_511), .B(n_396), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_496), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_498), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_521), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_511), .B(n_364), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_505), .Y(n_545) );
CKINVDCx6p67_ASAP7_75t_R g546 ( .A(n_500), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_500), .Y(n_547) );
AND2x6_ASAP7_75t_L g548 ( .A(n_490), .B(n_394), .Y(n_548) );
INVxp33_ASAP7_75t_L g549 ( .A(n_488), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_498), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_505), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_522), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_508), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_508), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_498), .Y(n_555) );
INVx4_ASAP7_75t_L g556 ( .A(n_490), .Y(n_556) );
INVx4_ASAP7_75t_L g557 ( .A(n_490), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_488), .B(n_327), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_492), .B(n_355), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_507), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_507), .B(n_468), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_517), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_498), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_517), .A2(n_330), .B1(n_332), .B2(n_326), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_508), .Y(n_565) );
AND3x1_ASAP7_75t_L g566 ( .A(n_523), .B(n_504), .C(n_482), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_556), .B(n_517), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_556), .B(n_517), .Y(n_568) );
NOR2x2_ASAP7_75t_L g569 ( .A(n_525), .B(n_375), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_559), .B(n_520), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_547), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_528), .A2(n_513), .B1(n_516), .B2(n_520), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_559), .B(n_487), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_530), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_549), .A2(n_487), .B1(n_502), .B2(n_483), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_524), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_556), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_547), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_546), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_546), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_540), .B(n_502), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_561), .B(n_519), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_543), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_527), .B(n_522), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_531), .B(n_522), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_560), .A2(n_473), .B1(n_357), .B2(n_386), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_528), .A2(n_516), .B1(n_513), .B2(n_495), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_560), .A2(n_375), .B1(n_404), .B2(n_393), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_540), .B(n_335), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_556), .B(n_522), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_529), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_557), .B(n_522), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_540), .B(n_335), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_558), .B(n_337), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_544), .B(n_557), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
OAI22x1_ASAP7_75t_SL g599 ( .A1(n_525), .A2(n_404), .B1(n_425), .B2(n_393), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_525), .B(n_327), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_525), .B(n_482), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_564), .B(n_351), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_562), .B(n_336), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_525), .B(n_504), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_534), .A2(n_386), .B1(n_401), .B2(n_345), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_562), .A2(n_521), .B(n_489), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_537), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_528), .B(n_356), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_562), .B(n_491), .Y(n_609) );
INVxp33_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_528), .A2(n_401), .B1(n_405), .B2(n_345), .Y(n_611) );
OR2x6_ASAP7_75t_L g612 ( .A(n_534), .B(n_514), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_545), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_545), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_528), .B(n_356), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_551), .B(n_514), .C(n_515), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_551), .Y(n_617) );
NOR2xp67_ASAP7_75t_L g618 ( .A(n_553), .B(n_515), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_528), .A2(n_495), .B1(n_501), .B2(n_491), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_528), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_553), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_548), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_554), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_554), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_548), .A2(n_427), .B1(n_440), .B2(n_405), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_565), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_534), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_548), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_543), .B(n_338), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_534), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_534), .B(n_506), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_548), .B(n_501), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_548), .A2(n_440), .B1(n_446), .B2(n_427), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_548), .A2(n_512), .B1(n_343), .B2(n_349), .Y(n_635) );
NOR2x2_ASAP7_75t_L g636 ( .A(n_542), .B(n_425), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_543), .B(n_342), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_543), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_543), .A2(n_512), .B1(n_350), .B2(n_359), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_543), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_552), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_535), .A2(n_446), .B1(n_334), .B2(n_409), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_552), .B(n_417), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_573), .B(n_331), .Y(n_644) );
NOR3xp33_ASAP7_75t_SL g645 ( .A(n_574), .B(n_409), .C(n_334), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_585), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_582), .B(n_415), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_585), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_606), .A2(n_489), .B(n_555), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_616), .A2(n_474), .B(n_403), .C(n_377), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_571), .A2(n_389), .B(n_392), .C(n_369), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_570), .B(n_415), .Y(n_652) );
NOR3xp33_ASAP7_75t_SL g653 ( .A(n_605), .B(n_439), .C(n_421), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_575), .B(n_597), .Y(n_654) );
AND2x6_ASAP7_75t_L g655 ( .A(n_628), .B(n_394), .Y(n_655) );
NOR2xp67_ASAP7_75t_L g656 ( .A(n_588), .B(n_421), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_598), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_630), .A2(n_563), .B(n_555), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_579), .B(n_439), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_613), .Y(n_660) );
OR2x6_ASAP7_75t_SL g661 ( .A(n_580), .B(n_448), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_632), .B(n_448), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_611), .A2(n_451), .B(n_449), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_630), .A2(n_563), .B(n_550), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_637), .A2(n_563), .B(n_550), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_577), .Y(n_666) );
INVx5_ASAP7_75t_L g667 ( .A(n_620), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_601), .A2(n_426), .B1(n_406), .B2(n_407), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_637), .A2(n_380), .B(n_340), .Y(n_669) );
BUFx4f_ASAP7_75t_L g670 ( .A(n_612), .Y(n_670) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_585), .Y(n_671) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_585), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_566), .A2(n_451), .B1(n_449), .B2(n_329), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_600), .B(n_426), .Y(n_674) );
AO32x1_ASAP7_75t_L g675 ( .A1(n_638), .A2(n_494), .A3(n_493), .B1(n_485), .B2(n_353), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_636), .Y(n_676) );
OR2x6_ASAP7_75t_L g677 ( .A(n_612), .B(n_465), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_602), .B(n_333), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_622), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_591), .B(n_424), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_572), .B(n_428), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_572), .B(n_428), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_619), .B(n_635), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_567), .A2(n_418), .B(n_408), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_625), .Y(n_685) );
BUFx2_ASAP7_75t_SL g686 ( .A(n_634), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_569), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_631), .A2(n_635), .B1(n_619), .B2(n_612), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_596), .B(n_416), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_599), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_629), .B(n_430), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_640), .A2(n_358), .B(n_348), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_609), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_595), .B(n_419), .Y(n_694) );
OR2x6_ASAP7_75t_L g695 ( .A(n_601), .B(n_465), .Y(n_695) );
BUFx4f_ASAP7_75t_L g696 ( .A(n_604), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_589), .B(n_433), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_583), .B(n_420), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_583), .B(n_433), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_607), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_609), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_614), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_639), .A2(n_589), .B1(n_618), .B2(n_568), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_568), .A2(n_365), .B(n_361), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_633), .A2(n_437), .B(n_444), .C(n_434), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_633), .B(n_457), .Y(n_706) );
INVxp67_ASAP7_75t_L g707 ( .A(n_642), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_603), .A2(n_452), .B1(n_455), .B2(n_450), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_639), .A2(n_578), .B1(n_584), .B2(n_576), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_593), .A2(n_456), .B(n_459), .C(n_458), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_592), .A2(n_368), .B(n_367), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_603), .A2(n_376), .B(n_372), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_590), .B(n_463), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_624), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_627), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_617), .A2(n_479), .B1(n_347), .B2(n_360), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_621), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_623), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_626), .A2(n_461), .B1(n_379), .B2(n_385), .C(n_384), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_608), .B(n_615), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_594), .A2(n_398), .B(n_395), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_586), .A2(n_476), .B1(n_453), .B2(n_400), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_586), .A2(n_411), .B(n_402), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_641), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_643), .Y(n_725) );
BUFx3_ASAP7_75t_L g726 ( .A(n_587), .Y(n_726) );
CKINVDCx11_ASAP7_75t_R g727 ( .A(n_587), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_574), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_606), .A2(n_414), .B(n_412), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_571), .B(n_468), .Y(n_730) );
AOI21x1_ASAP7_75t_L g731 ( .A1(n_606), .A2(n_536), .B(n_526), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_574), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_606), .A2(n_423), .B(n_422), .Y(n_733) );
INVx6_ASAP7_75t_L g734 ( .A(n_579), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_574), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_606), .A2(n_432), .B(n_431), .Y(n_736) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_581), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_598), .Y(n_738) );
OR2x6_ASAP7_75t_L g739 ( .A(n_605), .B(n_435), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_606), .A2(n_443), .B(n_436), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_574), .B(n_22), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_598), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_612), .A2(n_454), .B1(n_460), .B2(n_445), .Y(n_743) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_574), .B(n_397), .C(n_382), .Y(n_744) );
BUFx3_ASAP7_75t_L g745 ( .A(n_574), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_612), .A2(n_466), .B1(n_467), .B2(n_464), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_573), .B(n_381), .Y(n_747) );
AOI21x1_ASAP7_75t_L g748 ( .A1(n_606), .A2(n_541), .B(n_539), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g749 ( .A(n_620), .B(n_387), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_572), .B(n_390), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_606), .A2(n_477), .B(n_471), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_573), .B(n_470), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_572), .B(n_478), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_573), .B(n_480), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_610), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_606), .A2(n_541), .B(n_539), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_601), .A2(n_510), .B1(n_518), .B2(n_498), .Y(n_757) );
BUFx3_ASAP7_75t_L g758 ( .A(n_574), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_718), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_745), .Y(n_760) );
OAI221xp5_ASAP7_75t_L g761 ( .A1(n_668), .A2(n_413), .B1(n_438), .B2(n_447), .C(n_481), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_756), .A2(n_447), .B(n_438), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_729), .A2(n_541), .B(n_539), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_733), .A2(n_481), .B(n_472), .Y(n_764) );
AO31x2_ASAP7_75t_L g765 ( .A1(n_736), .A2(n_485), .A3(n_494), .B(n_493), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_707), .B(n_22), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_674), .A2(n_510), .B1(n_518), .B2(n_494), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_758), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_695), .B(n_23), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g770 ( .A1(n_739), .A2(n_518), .B1(n_510), .B2(n_26), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_740), .A2(n_518), .B(n_510), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_714), .A2(n_518), .B1(n_510), .B2(n_27), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_654), .B(n_23), .Y(n_773) );
AO22x1_ASAP7_75t_L g774 ( .A1(n_676), .A2(n_29), .B1(n_24), .B2(n_28), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_739), .A2(n_533), .B1(n_532), .B2(n_31), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_728), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_645), .B(n_533), .C(n_532), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_751), .A2(n_127), .B(n_126), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_714), .A2(n_33), .B1(n_30), .B2(n_31), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_700), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_673), .A2(n_34), .B1(n_35), .B2(n_36), .C(n_38), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_698), .B(n_34), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_649), .A2(n_533), .B(n_532), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_715), .Y(n_784) );
AO31x2_ASAP7_75t_L g785 ( .A1(n_722), .A2(n_533), .A3(n_532), .B(n_39), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_720), .A2(n_533), .B(n_532), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_739), .A2(n_39), .B1(n_35), .B2(n_38), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_734), .B(n_40), .Y(n_788) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_646), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_646), .Y(n_790) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_731), .A2(n_132), .B(n_128), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_755), .Y(n_792) );
A2O1A1Ixp33_ASAP7_75t_L g793 ( .A1(n_689), .A2(n_46), .B(n_44), .C(n_45), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_694), .B(n_644), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_717), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g796 ( .A(n_661), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_702), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_666), .Y(n_798) );
INVx4_ASAP7_75t_L g799 ( .A(n_737), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_735), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_686), .A2(n_48), .B1(n_46), .B2(n_47), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_657), .Y(n_802) );
O2A1O1Ixp33_ASAP7_75t_L g803 ( .A1(n_705), .A2(n_49), .B(n_47), .C(n_48), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_660), .B(n_49), .Y(n_804) );
AO32x2_ASAP7_75t_L g805 ( .A1(n_722), .A2(n_50), .A3(n_52), .B1(n_53), .B2(n_55), .Y(n_805) );
AO32x2_ASAP7_75t_L g806 ( .A1(n_743), .A2(n_50), .A3(n_52), .B1(n_55), .B2(n_56), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_693), .B(n_56), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_738), .Y(n_808) );
O2A1O1Ixp33_ASAP7_75t_SL g809 ( .A1(n_701), .A2(n_139), .B(n_140), .C(n_136), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_647), .B(n_57), .Y(n_810) );
O2A1O1Ixp33_ASAP7_75t_SL g811 ( .A1(n_709), .A2(n_208), .B(n_322), .C(n_321), .Y(n_811) );
AO31x2_ASAP7_75t_L g812 ( .A1(n_709), .A2(n_58), .A3(n_60), .B(n_61), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_646), .A2(n_143), .B(n_142), .Y(n_813) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_732), .Y(n_814) );
INVx4_ASAP7_75t_L g815 ( .A(n_677), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_662), .B(n_652), .Y(n_816) );
AO31x2_ASAP7_75t_L g817 ( .A1(n_703), .A2(n_60), .A3(n_62), .B(n_63), .Y(n_817) );
AO32x2_ASAP7_75t_L g818 ( .A1(n_743), .A2(n_62), .A3(n_63), .B1(n_64), .B2(n_65), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_648), .A2(n_148), .B(n_146), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_742), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_748), .A2(n_152), .B(n_151), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_695), .B(n_64), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_685), .B(n_66), .Y(n_823) );
CKINVDCx9p33_ASAP7_75t_R g824 ( .A(n_690), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_L g825 ( .A1(n_710), .A2(n_66), .B(n_69), .C(n_70), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_692), .A2(n_154), .B(n_153), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_648), .A2(n_158), .B(n_157), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_692), .A2(n_160), .B(n_159), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_754), .Y(n_829) );
BUFx3_ASAP7_75t_L g830 ( .A(n_687), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_650), .A2(n_69), .B(n_71), .C(n_72), .Y(n_831) );
O2A1O1Ixp33_ASAP7_75t_L g832 ( .A1(n_651), .A2(n_71), .B(n_73), .C(n_74), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_648), .A2(n_162), .B(n_161), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_696), .B(n_73), .Y(n_834) );
INVx3_ASAP7_75t_L g835 ( .A(n_666), .Y(n_835) );
NOR2xp67_ASAP7_75t_L g836 ( .A(n_744), .B(n_74), .Y(n_836) );
O2A1O1Ixp33_ASAP7_75t_SL g837 ( .A1(n_683), .A2(n_221), .B(n_319), .C(n_317), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_713), .A2(n_75), .B1(n_76), .B2(n_77), .C(n_78), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_746), .B(n_76), .Y(n_839) );
AO31x2_ASAP7_75t_L g840 ( .A1(n_703), .A2(n_79), .A3(n_81), .B(n_82), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_677), .Y(n_841) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_671), .Y(n_842) );
BUFx2_ASAP7_75t_L g843 ( .A(n_677), .Y(n_843) );
BUFx2_ASAP7_75t_L g844 ( .A(n_696), .Y(n_844) );
BUFx8_ASAP7_75t_L g845 ( .A(n_741), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_746), .B(n_79), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_663), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_847) );
AOI21xp5_ASAP7_75t_L g848 ( .A1(n_671), .A2(n_170), .B(n_168), .Y(n_848) );
AO31x2_ASAP7_75t_L g849 ( .A1(n_688), .A2(n_85), .A3(n_87), .B(n_88), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_747), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_704), .A2(n_172), .B(n_171), .Y(n_851) );
BUFx10_ASAP7_75t_L g852 ( .A(n_659), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_727), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_656), .B(n_85), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g855 ( .A1(n_671), .A2(n_175), .B(n_174), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_653), .B(n_87), .Y(n_856) );
AO31x2_ASAP7_75t_L g857 ( .A1(n_716), .A2(n_88), .A3(n_89), .B(n_90), .Y(n_857) );
OAI211xp5_ASAP7_75t_L g858 ( .A1(n_719), .A2(n_89), .B(n_91), .C(n_93), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_672), .A2(n_240), .B(n_315), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_752), .Y(n_860) );
AO21x2_ASAP7_75t_L g861 ( .A1(n_723), .A2(n_238), .B(n_314), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_670), .A2(n_94), .B1(n_96), .B2(n_97), .Y(n_862) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_672), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_678), .A2(n_97), .B(n_99), .C(n_100), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_757), .B(n_100), .C(n_101), .Y(n_865) );
AO31x2_ASAP7_75t_L g866 ( .A1(n_716), .A2(n_102), .A3(n_103), .B(n_104), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_726), .A2(n_102), .B1(n_105), .B2(n_106), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_753), .A2(n_105), .B1(n_108), .B2(n_109), .Y(n_868) );
O2A1O1Ixp33_ASAP7_75t_SL g869 ( .A1(n_750), .A2(n_245), .B(n_310), .C(n_309), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_699), .B(n_108), .Y(n_870) );
O2A1O1Ixp5_ASAP7_75t_SL g871 ( .A1(n_681), .A2(n_243), .B(n_306), .C(n_305), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_725), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_682), .A2(n_110), .B1(n_112), .B2(n_113), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_730), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_667), .Y(n_875) );
AO31x2_ASAP7_75t_L g876 ( .A1(n_658), .A2(n_112), .A3(n_113), .B(n_114), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_706), .A2(n_117), .B1(n_118), .B2(n_176), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_679), .A2(n_117), .B1(n_118), .B2(n_180), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_680), .B(n_185), .Y(n_879) );
OR2x2_ASAP7_75t_L g880 ( .A(n_708), .B(n_186), .Y(n_880) );
AO31x2_ASAP7_75t_L g881 ( .A1(n_664), .A2(n_187), .A3(n_190), .B(n_191), .Y(n_881) );
A2O1A1Ixp33_ASAP7_75t_L g882 ( .A1(n_711), .A2(n_192), .B(n_194), .C(n_197), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_667), .B(n_198), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_712), .B(n_201), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_712), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_SL g886 ( .A1(n_697), .A2(n_202), .B(n_204), .C(n_206), .Y(n_886) );
A2O1A1Ixp33_ASAP7_75t_L g887 ( .A1(n_721), .A2(n_207), .B(n_209), .C(n_210), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_679), .A2(n_211), .B1(n_212), .B2(n_213), .Y(n_888) );
BUFx12f_ASAP7_75t_L g889 ( .A(n_655), .Y(n_889) );
AO31x2_ASAP7_75t_L g890 ( .A1(n_665), .A2(n_214), .A3(n_215), .B(n_216), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_667), .A2(n_217), .B1(n_218), .B2(n_219), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_724), .Y(n_892) );
O2A1O1Ixp33_ASAP7_75t_SL g893 ( .A1(n_691), .A2(n_220), .B(n_223), .C(n_224), .Y(n_893) );
OAI21xp5_ASAP7_75t_L g894 ( .A1(n_684), .A2(n_225), .B(n_228), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_749), .A2(n_232), .B1(n_233), .B2(n_235), .Y(n_895) );
NAND3xp33_ASAP7_75t_SL g896 ( .A(n_760), .B(n_669), .C(n_749), .Y(n_896) );
AOI21xp33_ASAP7_75t_SL g897 ( .A1(n_853), .A2(n_236), .B(n_241), .Y(n_897) );
AOI32xp33_ASAP7_75t_L g898 ( .A1(n_769), .A2(n_655), .A3(n_246), .B1(n_248), .B2(n_252), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_766), .A2(n_655), .B1(n_675), .B2(n_253), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_795), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_783), .A2(n_675), .B(n_655), .Y(n_901) );
BUFx6f_ASAP7_75t_L g902 ( .A(n_789), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_797), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_788), .A2(n_257), .B1(n_261), .B2(n_263), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_759), .Y(n_905) );
INVx1_ASAP7_75t_SL g906 ( .A(n_800), .Y(n_906) );
OAI21xp33_ASAP7_75t_L g907 ( .A1(n_794), .A2(n_265), .B(n_269), .Y(n_907) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_850), .A2(n_270), .B(n_273), .C(n_275), .Y(n_908) );
OA21x2_ASAP7_75t_L g909 ( .A1(n_791), .A2(n_277), .B(n_280), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_829), .B(n_282), .Y(n_910) );
OR2x6_ASAP7_75t_L g911 ( .A(n_799), .B(n_284), .Y(n_911) );
OA21x2_ASAP7_75t_L g912 ( .A1(n_821), .A2(n_287), .B(n_289), .Y(n_912) );
OAI21xp5_ASAP7_75t_L g913 ( .A1(n_885), .A2(n_290), .B(n_291), .Y(n_913) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_788), .A2(n_292), .B1(n_293), .B2(n_294), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_792), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_844), .B(n_295), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_804), .Y(n_917) );
CKINVDCx11_ASAP7_75t_R g918 ( .A(n_796), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_773), .A2(n_301), .B(n_302), .Y(n_919) );
A2O1A1Ixp33_ASAP7_75t_L g920 ( .A1(n_832), .A2(n_324), .B(n_803), .C(n_831), .Y(n_920) );
INVx1_ASAP7_75t_SL g921 ( .A(n_776), .Y(n_921) );
BUFx2_ASAP7_75t_L g922 ( .A(n_768), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_814), .B(n_843), .Y(n_923) );
OR2x6_ASAP7_75t_L g924 ( .A(n_799), .B(n_815), .Y(n_924) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_822), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_872), .B(n_816), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_780), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_856), .B(n_834), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_807), .Y(n_929) );
A2O1A1Ixp33_ASAP7_75t_L g930 ( .A1(n_825), .A2(n_854), .B(n_870), .C(n_782), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_784), .B(n_810), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_823), .A2(n_846), .B1(n_839), .B2(n_841), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_771), .A2(n_763), .B(n_811), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_857), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_802), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_808), .Y(n_936) );
BUFx2_ASAP7_75t_L g937 ( .A(n_889), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_820), .B(n_879), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_857), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_775), .A2(n_787), .B1(n_801), .B2(n_770), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_892), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_765), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_857), .Y(n_943) );
INVx3_ASAP7_75t_L g944 ( .A(n_883), .Y(n_944) );
OAI211xp5_ASAP7_75t_L g945 ( .A1(n_862), .A2(n_838), .B(n_858), .C(n_781), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_866), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_761), .A2(n_867), .B1(n_779), .B2(n_864), .C(n_793), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_765), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_798), .B(n_835), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_866), .Y(n_950) );
A2O1A1Ixp33_ASAP7_75t_L g951 ( .A1(n_836), .A2(n_826), .B(n_828), .C(n_865), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_852), .A2(n_845), .B1(n_874), .B2(n_830), .Y(n_952) );
AO31x2_ASAP7_75t_L g953 ( .A1(n_772), .A2(n_877), .A3(n_882), .B(n_887), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_852), .A2(n_845), .B1(n_880), .B2(n_884), .Y(n_954) );
NAND2xp5_ASAP7_75t_SL g955 ( .A(n_883), .B(n_842), .Y(n_955) );
OA21x2_ASAP7_75t_L g956 ( .A1(n_778), .A2(n_894), .B(n_851), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_866), .Y(n_957) );
NAND2x1p5_ASAP7_75t_L g958 ( .A(n_790), .B(n_863), .Y(n_958) );
BUFx6f_ASAP7_75t_L g959 ( .A(n_790), .Y(n_959) );
INVx3_ASAP7_75t_L g960 ( .A(n_842), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_847), .A2(n_873), .B1(n_767), .B2(n_895), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_824), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_878), .A2(n_868), .B1(n_888), .B2(n_875), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_806), .B(n_818), .Y(n_964) );
INVxp67_ASAP7_75t_L g965 ( .A(n_774), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_806), .Y(n_966) );
OR2x2_ASAP7_75t_L g967 ( .A(n_798), .B(n_835), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_806), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_891), .A2(n_863), .B1(n_764), .B2(n_777), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_818), .Y(n_970) );
OAI211xp5_ASAP7_75t_L g971 ( .A1(n_809), .A2(n_819), .B(n_859), .C(n_848), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_849), .B(n_840), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_849), .B(n_840), .Y(n_973) );
AO21x2_ASAP7_75t_L g974 ( .A1(n_837), .A2(n_886), .B(n_861), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_813), .A2(n_827), .B1(n_855), .B2(n_833), .Y(n_975) );
NOR2xp67_ASAP7_75t_SL g976 ( .A(n_818), .B(n_805), .Y(n_976) );
OA21x2_ASAP7_75t_L g977 ( .A1(n_871), .A2(n_890), .B(n_881), .Y(n_977) );
INVx3_ASAP7_75t_L g978 ( .A(n_817), .Y(n_978) );
BUFx2_ASAP7_75t_L g979 ( .A(n_805), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_869), .A2(n_893), .B(n_890), .Y(n_980) );
AO21x2_ASAP7_75t_L g981 ( .A1(n_785), .A2(n_881), .B(n_817), .Y(n_981) );
OA21x2_ASAP7_75t_L g982 ( .A1(n_785), .A2(n_765), .B(n_812), .Y(n_982) );
NOR3xp33_ASAP7_75t_L g983 ( .A(n_876), .B(n_538), .C(n_574), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_876), .B(n_785), .Y(n_984) );
BUFx4f_ASAP7_75t_L g985 ( .A(n_876), .Y(n_985) );
INVxp67_ASAP7_75t_SL g986 ( .A(n_776), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_760), .Y(n_987) );
OAI21x1_ASAP7_75t_L g988 ( .A1(n_762), .A2(n_783), .B(n_756), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_829), .B(n_654), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_788), .A2(n_605), .B1(n_625), .B2(n_611), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_769), .B(n_601), .Y(n_991) );
O2A1O1Ixp33_ASAP7_75t_L g992 ( .A1(n_794), .A2(n_743), .B(n_746), .C(n_823), .Y(n_992) );
A2O1A1Ixp33_ASAP7_75t_L g993 ( .A1(n_794), .A2(n_860), .B(n_850), .C(n_829), .Y(n_993) );
BUFx3_ASAP7_75t_L g994 ( .A(n_760), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_800), .B(n_605), .Y(n_995) );
A2O1A1Ixp33_ASAP7_75t_L g996 ( .A1(n_794), .A2(n_860), .B(n_850), .C(n_829), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g997 ( .A1(n_766), .A2(n_605), .B1(n_574), .B2(n_612), .Y(n_997) );
A2O1A1Ixp33_ASAP7_75t_L g998 ( .A1(n_794), .A2(n_860), .B(n_850), .C(n_829), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_795), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_794), .A2(n_566), .B1(n_616), .B2(n_650), .C(n_829), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_795), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_795), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_760), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_800), .B(n_605), .Y(n_1004) );
INVx4_ASAP7_75t_L g1005 ( .A(n_799), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_769), .B(n_601), .Y(n_1006) );
AOI222xp33_ASAP7_75t_L g1007 ( .A1(n_796), .A2(n_599), .B1(n_601), .B2(n_604), .C1(n_690), .C2(n_670), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_769), .B(n_601), .Y(n_1008) );
AOI21xp5_ASAP7_75t_L g1009 ( .A1(n_783), .A2(n_786), .B(n_733), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_783), .A2(n_786), .B(n_733), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g1011 ( .A(n_789), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_783), .A2(n_786), .B(n_733), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_769), .B(n_601), .Y(n_1013) );
BUFx6f_ASAP7_75t_L g1014 ( .A(n_789), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_769), .B(n_601), .Y(n_1015) );
OAI21xp5_ASAP7_75t_L g1016 ( .A1(n_885), .A2(n_733), .B(n_729), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_905), .B(n_900), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_903), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_990), .A2(n_1007), .B1(n_1000), .B2(n_928), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_999), .B(n_1001), .Y(n_1020) );
NAND2xp33_ASAP7_75t_SL g1021 ( .A(n_944), .B(n_955), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1000), .B(n_926), .Y(n_1022) );
INVx3_ASAP7_75t_SL g1023 ( .A(n_962), .Y(n_1023) );
BUFx3_ASAP7_75t_L g1024 ( .A(n_922), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_942), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_915), .Y(n_1026) );
OR2x6_ASAP7_75t_L g1027 ( .A(n_911), .B(n_924), .Y(n_1027) );
OAI21xp5_ASAP7_75t_L g1028 ( .A1(n_992), .A2(n_920), .B(n_930), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_993), .B(n_996), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1030 ( .A1(n_997), .A2(n_932), .B1(n_998), .B2(n_954), .C(n_1004), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1002), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_906), .B(n_921), .Y(n_1032) );
OR2x6_ASAP7_75t_L g1033 ( .A(n_911), .B(n_924), .Y(n_1033) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_1005), .Y(n_1034) );
OA21x2_ASAP7_75t_L g1035 ( .A1(n_984), .A2(n_973), .B(n_972), .Y(n_1035) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_986), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_989), .B(n_995), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_906), .B(n_921), .Y(n_1038) );
OR2x6_ASAP7_75t_L g1039 ( .A(n_911), .B(n_924), .Y(n_1039) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_948), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_927), .B(n_935), .Y(n_1041) );
NAND3xp33_ASAP7_75t_L g1042 ( .A(n_983), .B(n_957), .C(n_950), .Y(n_1042) );
OAI21xp5_ASAP7_75t_L g1043 ( .A1(n_945), .A2(n_951), .B(n_940), .Y(n_1043) );
INVx2_ASAP7_75t_L g1044 ( .A(n_988), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_1007), .A2(n_965), .B1(n_947), .B2(n_940), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_936), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_941), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_989), .B(n_929), .Y(n_1048) );
OAI21xp33_ASAP7_75t_L g1049 ( .A1(n_972), .A2(n_973), .B(n_943), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_991), .B(n_1006), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_947), .A2(n_1015), .B1(n_1013), .B2(n_1008), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_994), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_925), .B(n_923), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_902), .Y(n_1054) );
AO21x2_ASAP7_75t_L g1055 ( .A1(n_980), .A2(n_901), .B(n_933), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_987), .B(n_1003), .Y(n_1056) );
BUFx8_ASAP7_75t_SL g1057 ( .A(n_937), .Y(n_1057) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_916), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_960), .Y(n_1059) );
OA21x2_ASAP7_75t_L g1060 ( .A1(n_934), .A2(n_939), .B(n_946), .Y(n_1060) );
AO31x2_ASAP7_75t_L g1061 ( .A1(n_979), .A2(n_970), .A3(n_968), .B(n_966), .Y(n_1061) );
NAND2x1_ASAP7_75t_L g1062 ( .A(n_902), .B(n_959), .Y(n_1062) );
INVx3_ASAP7_75t_L g1063 ( .A(n_959), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_931), .Y(n_1064) );
OR2x6_ASAP7_75t_L g1065 ( .A(n_958), .B(n_913), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1011), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_917), .B(n_964), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_931), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_952), .B(n_910), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1011), .Y(n_1070) );
INVx6_ASAP7_75t_L g1071 ( .A(n_1014), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1014), .Y(n_1072) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_967), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_982), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_982), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_976), .Y(n_1076) );
OA21x2_ASAP7_75t_L g1077 ( .A1(n_1012), .A2(n_1010), .B(n_1009), .Y(n_1077) );
INVx3_ASAP7_75t_L g1078 ( .A(n_985), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_981), .B(n_978), .Y(n_1079) );
OR2x6_ASAP7_75t_L g1080 ( .A(n_949), .B(n_938), .Y(n_1080) );
OR2x6_ASAP7_75t_L g1081 ( .A(n_949), .B(n_938), .Y(n_1081) );
AO221x2_ASAP7_75t_L g1082 ( .A1(n_963), .A2(n_919), .B1(n_969), .B2(n_961), .C(n_985), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_909), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_896), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_904), .B(n_914), .Y(n_1085) );
INVx2_ASAP7_75t_L g1086 ( .A(n_909), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_918), .B(n_1016), .Y(n_1087) );
AOI21xp5_ASAP7_75t_SL g1088 ( .A1(n_956), .A2(n_907), .B(n_912), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_912), .Y(n_1089) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_898), .A2(n_897), .B1(n_969), .B2(n_899), .C(n_908), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_953), .B(n_977), .Y(n_1091) );
OAI21x1_ASAP7_75t_L g1092 ( .A1(n_975), .A2(n_977), .B(n_974), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_953), .B(n_971), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1094 ( .A1(n_953), .A2(n_1000), .B1(n_566), .B2(n_650), .C(n_651), .Y(n_1094) );
NAND4xp25_ASAP7_75t_L g1095 ( .A(n_1007), .B(n_1000), .C(n_504), .D(n_515), .Y(n_1095) );
AO21x2_ASAP7_75t_L g1096 ( .A1(n_983), .A2(n_984), .B(n_980), .Y(n_1096) );
INVxp33_ASAP7_75t_SL g1097 ( .A(n_918), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_905), .B(n_900), .Y(n_1098) );
AO21x2_ASAP7_75t_L g1099 ( .A1(n_983), .A2(n_984), .B(n_980), .Y(n_1099) );
OAI31xp33_ASAP7_75t_L g1100 ( .A1(n_1095), .A2(n_1045), .A3(n_1030), .B(n_1019), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1067), .B(n_1076), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_1027), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1067), .B(n_1079), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_1025), .Y(n_1104) );
INVx3_ASAP7_75t_L g1105 ( .A(n_1078), .Y(n_1105) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_1078), .B(n_1079), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1060), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1060), .Y(n_1108) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_1024), .Y(n_1109) );
OAI31xp33_ASAP7_75t_L g1110 ( .A1(n_1045), .A2(n_1019), .A3(n_1051), .B(n_1085), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1022), .B(n_1053), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1061), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1061), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1020), .B(n_1048), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_1074), .B(n_1075), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1048), .B(n_1017), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1017), .B(n_1098), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1098), .B(n_1082), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1082), .B(n_1041), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1061), .Y(n_1120) );
AND2x4_ASAP7_75t_SL g1121 ( .A(n_1027), .B(n_1033), .Y(n_1121) );
OR2x6_ASAP7_75t_L g1122 ( .A(n_1033), .B(n_1039), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1082), .B(n_1041), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1037), .B(n_1064), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_1094), .A2(n_1043), .B1(n_1051), .B2(n_1028), .C(n_1029), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1025), .B(n_1040), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1061), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_1032), .B(n_1038), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1036), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1040), .B(n_1035), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1068), .B(n_1050), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1049), .Y(n_1132) );
INVx3_ASAP7_75t_SL g1133 ( .A(n_1039), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1077), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_1093), .B(n_1065), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1042), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1137 ( .A(n_1093), .B(n_1065), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1050), .B(n_1018), .Y(n_1138) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_1087), .A2(n_1058), .B1(n_1081), .B2(n_1080), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1073), .B(n_1080), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1026), .B(n_1031), .Y(n_1141) );
BUFx3_ASAP7_75t_L g1142 ( .A(n_1062), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1091), .Y(n_1143) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_1071), .Y(n_1144) );
INVx1_ASAP7_75t_SL g1145 ( .A(n_1057), .Y(n_1145) );
AO21x2_ASAP7_75t_L g1146 ( .A1(n_1088), .A2(n_1083), .B(n_1089), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1046), .B(n_1047), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1103), .B(n_1101), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1107), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1107), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1103), .B(n_1101), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1128), .B(n_1099), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1118), .B(n_1084), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1128), .B(n_1099), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1119), .B(n_1096), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1108), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1123), .B(n_1055), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1114), .B(n_1092), .Y(n_1158) );
INVx3_ASAP7_75t_L g1159 ( .A(n_1146), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1116), .B(n_1143), .Y(n_1160) );
NOR4xp25_ASAP7_75t_SL g1161 ( .A(n_1102), .B(n_1021), .C(n_1090), .D(n_1059), .Y(n_1161) );
INVx3_ASAP7_75t_L g1162 ( .A(n_1146), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1106), .B(n_1044), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1104), .B(n_1069), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1106), .B(n_1072), .Y(n_1165) );
AND2x4_ASAP7_75t_L g1166 ( .A(n_1135), .B(n_1083), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1135), .B(n_1089), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1126), .B(n_1054), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1126), .B(n_1117), .Y(n_1169) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_1122), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1129), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1130), .B(n_1070), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1138), .B(n_1066), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1138), .B(n_1072), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1137), .B(n_1086), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1171), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1149), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1160), .B(n_1141), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1149), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1169), .B(n_1132), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1148), .B(n_1132), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1148), .B(n_1131), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1158), .B(n_1112), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1150), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_1153), .A2(n_1100), .B1(n_1110), .B2(n_1125), .Y(n_1185) );
NAND3xp33_ASAP7_75t_SL g1186 ( .A(n_1161), .B(n_1145), .C(n_1100), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1151), .B(n_1097), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1173), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_1152), .B(n_1113), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1157), .B(n_1120), .Y(n_1190) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1156), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1152), .B(n_1127), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1155), .B(n_1115), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1156), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1154), .B(n_1140), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1181), .B(n_1164), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1180), .B(n_1168), .Y(n_1197) );
NAND3xp33_ASAP7_75t_L g1198 ( .A(n_1185), .B(n_1110), .C(n_1136), .Y(n_1198) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_1187), .A2(n_1139), .B1(n_1122), .B2(n_1133), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1177), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1195), .B(n_1172), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1183), .B(n_1175), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1183), .B(n_1175), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1191), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1193), .B(n_1163), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1190), .B(n_1174), .Y(n_1206) );
NOR2xp33_ASAP7_75t_L g1207 ( .A(n_1176), .B(n_1097), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1193), .B(n_1165), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1190), .B(n_1174), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1196), .B(n_1182), .Y(n_1210) );
XNOR2x1_ASAP7_75t_L g1211 ( .A(n_1198), .B(n_1056), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_1207), .A2(n_1186), .B1(n_1121), .B2(n_1102), .Y(n_1212) );
AOI211xp5_ASAP7_75t_L g1213 ( .A1(n_1199), .A2(n_1133), .B(n_1023), .C(n_1170), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1197), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1201), .B(n_1178), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1214), .Y(n_1216) );
O2A1O1Ixp33_ASAP7_75t_L g1217 ( .A1(n_1212), .A2(n_1052), .B(n_1034), .C(n_1124), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1210), .B(n_1206), .Y(n_1218) );
OAI322xp33_ASAP7_75t_L g1219 ( .A1(n_1211), .A2(n_1209), .A3(n_1189), .B1(n_1192), .B2(n_1188), .C1(n_1111), .C2(n_1184), .Y(n_1219) );
OAI221xp5_ASAP7_75t_SL g1220 ( .A1(n_1213), .A2(n_1189), .B1(n_1192), .B2(n_1202), .C(n_1203), .Y(n_1220) );
A2O1A1Ixp33_ASAP7_75t_L g1221 ( .A1(n_1217), .A2(n_1215), .B(n_1109), .C(n_1205), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1216), .B(n_1208), .Y(n_1222) );
NAND4xp25_ASAP7_75t_SL g1223 ( .A(n_1221), .B(n_1220), .C(n_1219), .D(n_1218), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1222), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1224), .Y(n_1225) );
NOR4xp25_ASAP7_75t_L g1226 ( .A(n_1223), .B(n_1147), .C(n_1144), .D(n_1162), .Y(n_1226) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_1225), .Y(n_1227) );
XNOR2xp5_ASAP7_75t_L g1228 ( .A(n_1227), .B(n_1226), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1228), .Y(n_1229) );
AOI222xp33_ASAP7_75t_SL g1230 ( .A1(n_1229), .A2(n_1105), .B1(n_1159), .B2(n_1162), .C1(n_1063), .C2(n_1179), .Y(n_1230) );
AOI222xp33_ASAP7_75t_L g1231 ( .A1(n_1230), .A2(n_1194), .B1(n_1142), .B2(n_1134), .C1(n_1204), .C2(n_1200), .Y(n_1231) );
UNKNOWN g1232 ( );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_1232), .A2(n_1204), .B1(n_1167), .B2(n_1166), .Y(n_1233) );
endmodule