module fake_jpeg_24958_n_109 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_12),
.B1(n_13),
.B2(n_22),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_22),
.B1(n_17),
.B2(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_53),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_58),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_20),
.B(n_19),
.C(n_31),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_59),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_14),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_0),
.B2(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_21),
.B1(n_20),
.B2(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_24),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_20),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_32),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_24),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_51),
.B(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_73),
.B1(n_55),
.B2(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_46),
.B1(n_52),
.B2(n_49),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_59),
.C(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_80),
.C(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_83),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_81),
.C(n_80),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_94),
.B(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_66),
.B1(n_68),
.B2(n_74),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_85),
.B(n_68),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_99),
.B(n_3),
.Y(n_102)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_72),
.B(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_103),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_93),
.A3(n_65),
.B1(n_83),
.B2(n_66),
.C1(n_11),
.C2(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_5),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_106),
.B(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_9),
.Y(n_109)
);


endmodule