module fake_netlist_1_7228_n_35 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_7;
wire n_27;
INVx2_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
BUFx6f_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_4), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_12), .B(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
NAND3xp33_ASAP7_75t_SL g15 ( .A(n_9), .B(n_0), .C(n_1), .Y(n_15) );
OA21x2_ASAP7_75t_L g16 ( .A1(n_7), .A2(n_2), .B(n_5), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_10), .B(n_6), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_7), .A2(n_2), .B1(n_5), .B2(n_6), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_13), .B(n_8), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_17), .B(n_8), .Y(n_20) );
AOI22xp33_ASAP7_75t_SL g21 ( .A1(n_18), .A2(n_8), .B1(n_11), .B2(n_16), .Y(n_21) );
INVxp33_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_16), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
OAI22xp33_ASAP7_75t_SL g26 ( .A1(n_23), .A2(n_20), .B1(n_19), .B2(n_21), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AOI321xp33_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_19), .A3(n_20), .B1(n_25), .B2(n_24), .C(n_14), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx5_ASAP7_75t_L g32 ( .A(n_28), .Y(n_32) );
NAND2x1p5_ASAP7_75t_L g33 ( .A(n_29), .B(n_24), .Y(n_33) );
AO22x2_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B1(n_30), .B2(n_20), .Y(n_34) );
AOI222xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_31), .B1(n_32), .B2(n_33), .C1(n_29), .C2(n_18), .Y(n_35) );
endmodule