module fake_jpeg_21850_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_48),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_33),
.Y(n_75)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_26),
.B1(n_34),
.B2(n_23),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_61),
.B1(n_65),
.B2(n_31),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_78),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_66),
.B1(n_77),
.B2(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_26),
.B1(n_34),
.B2(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_16),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_75),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_31),
.B(n_18),
.C(n_35),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_30),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_47),
.B(n_1),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_39),
.A2(n_27),
.B1(n_33),
.B2(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_18),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_91),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_40),
.B(n_27),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_58),
.B(n_59),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_53),
.B1(n_58),
.B2(n_68),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_93),
.B(n_100),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2x1_ASAP7_75t_R g149 ( 
.A(n_97),
.B(n_120),
.Y(n_149)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_20),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_20),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_113),
.B(n_119),
.Y(n_141)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_117),
.B1(n_58),
.B2(n_68),
.Y(n_123)
);

AO22x2_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_40),
.B1(n_52),
.B2(n_79),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_117),
.B1(n_105),
.B2(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_62),
.B(n_40),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_110),
.B(n_112),
.Y(n_148)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_47),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_35),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_38),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_127),
.B1(n_137),
.B2(n_144),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_131),
.B(n_118),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_59),
.C(n_72),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_147),
.C(n_41),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_92),
.B1(n_106),
.B2(n_121),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_88),
.B1(n_50),
.B2(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_38),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_38),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_31),
.B1(n_67),
.B2(n_18),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_36),
.C(n_50),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_18),
.B1(n_31),
.B2(n_50),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_103),
.B1(n_99),
.B2(n_108),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_105),
.B1(n_110),
.B2(n_98),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_155),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_154),
.B(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_166),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_87),
.B1(n_104),
.B2(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_102),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_84),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_94),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_88),
.B1(n_111),
.B2(n_119),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_174),
.B1(n_180),
.B2(n_150),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_124),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_171),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_80),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_150),
.C(n_130),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_41),
.B1(n_45),
.B2(n_36),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_45),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_35),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_133),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_182),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_141),
.B1(n_123),
.B2(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_141),
.A2(n_36),
.B1(n_82),
.B2(n_35),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_22),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_82),
.B1(n_85),
.B2(n_116),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_187),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_9),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_22),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_145),
.Y(n_186)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_145),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g246 ( 
.A(n_190),
.B(n_218),
.C(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_130),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_210),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_204),
.C(n_160),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_201),
.B1(n_202),
.B2(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_198),
.B(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_146),
.B1(n_134),
.B2(n_128),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_146),
.B1(n_134),
.B2(n_128),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_154),
.C(n_167),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_215),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_132),
.B(n_22),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_213),
.B(n_215),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_4),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_0),
.B(n_2),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_156),
.A2(n_0),
.B(n_2),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_217),
.A2(n_179),
.B1(n_153),
.B2(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_205),
.C(n_208),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_228),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_214),
.Y(n_229)
);

NOR2x1_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_239),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_243),
.B1(n_248),
.B2(n_217),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_196),
.A2(n_199),
.B1(n_212),
.B2(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_162),
.A3(n_174),
.B1(n_168),
.B2(n_164),
.C1(n_178),
.C2(n_187),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_193),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_176),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_194),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_238)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_3),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_6),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_13),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_249),
.B1(n_248),
.B2(n_241),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_207),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_10),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_190),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_261),
.C(n_264),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_226),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_231),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_216),
.B1(n_191),
.B2(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_213),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_260),
.B(n_272),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_255),
.B1(n_266),
.B2(n_240),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_276),
.B(n_282),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_230),
.B(n_245),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_250),
.B(n_220),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_246),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_225),
.C(n_228),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_288),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_216),
.B1(n_221),
.B2(n_202),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_279),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_224),
.B1(n_201),
.B2(n_239),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_242),
.B1(n_227),
.B2(n_195),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_262),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_300),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_288),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_300)
);

AO221x1_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_244),
.B1(n_227),
.B2(n_252),
.C(n_257),
.Y(n_301)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_278),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_277),
.B1(n_284),
.B2(n_291),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_273),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_281),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_237),
.Y(n_305)
);

HAxp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_237),
.CON(n_314),
.SN(n_314)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_223),
.B1(n_238),
.B2(n_283),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_274),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_316),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_314),
.B1(n_318),
.B2(n_320),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_296),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_285),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_304),
.C(n_303),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_259),
.C(n_273),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_298),
.C(n_293),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_258),
.B1(n_7),
.B2(n_8),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_300),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_310),
.A2(n_307),
.B(n_295),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_308),
.B(n_305),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_327),
.C(n_328),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_319),
.C(n_309),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_302),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_309),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_307),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_334),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_314),
.B(n_313),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_332),
.A2(n_333),
.B1(n_327),
.B2(n_326),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_311),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_11),
.Y(n_340)
);

NOR2x1_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_326),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_336),
.B(n_11),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_339),
.B(n_340),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_12),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_342),
.B(n_338),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_336),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_337),
.B1(n_206),
.B2(n_12),
.Y(n_346)
);

OAI321xp33_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_6),
.A3(n_7),
.B1(n_206),
.B2(n_341),
.C(n_275),
.Y(n_347)
);


endmodule