module fake_jpeg_30948_n_152 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_16),
.B1(n_24),
.B2(n_23),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_30),
.B1(n_38),
.B2(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_22),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_15),
.B(n_18),
.C(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_70),
.Y(n_86)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_69),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_15),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_11),
.B(n_14),
.C(n_10),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_74),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_61),
.B(n_11),
.C(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_5),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_53),
.B1(n_60),
.B2(n_48),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_60),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_81),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_41),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_75),
.C(n_69),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_50),
.B(n_33),
.C(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_9),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_7),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_77),
.B1(n_64),
.B2(n_72),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_73),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_75),
.C(n_83),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_90),
.C(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_70),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_80),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_82),
.B(n_67),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_46),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_98),
.B1(n_101),
.B2(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_85),
.C(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_94),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_125),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_109),
.Y(n_130)
);

OA21x2_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_115),
.B(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_132),
.Y(n_135)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_109),
.A3(n_113),
.B1(n_53),
.B2(n_95),
.C(n_34),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_34),
.C(n_95),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_113),
.C(n_62),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_121),
.B(n_125),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_136),
.A2(n_0),
.B(n_2),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_137),
.A2(n_130),
.B1(n_131),
.B2(n_39),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_9),
.B(n_1),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_0),
.B(n_2),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_141),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_144),
.B1(n_3),
.B2(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_135),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_143),
.A2(n_3),
.B(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_143),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_148),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_76),
.Y(n_152)
);


endmodule