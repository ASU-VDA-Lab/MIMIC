module fake_jpeg_2444_n_571 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_571);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_571;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_31),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_65),
.B(n_69),
.Y(n_160)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_67),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_71),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_74),
.Y(n_188)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_75),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_80),
.B(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

HAxp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_1),
.CON(n_84),
.SN(n_84)
);

INVx2_ASAP7_75t_R g185 ( 
.A(n_84),
.Y(n_185)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_85),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_104),
.B1(n_48),
.B2(n_30),
.Y(n_144)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_96),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_103),
.B(n_109),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_27),
.B1(n_48),
.B2(n_42),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_105),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_110),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

CKINVDCx9p33_ASAP7_75t_R g181 ( 
.A(n_111),
.Y(n_181)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_112),
.B(n_114),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_19),
.B(n_28),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_124),
.Y(n_154)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_118),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_2),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_120),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_34),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_125),
.Y(n_204)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_24),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_123),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_126),
.B(n_8),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_21),
.B(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_127),
.B(n_14),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_58),
.A2(n_49),
.B1(n_51),
.B2(n_27),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_129),
.A2(n_181),
.B1(n_151),
.B2(n_199),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_49),
.B1(n_24),
.B2(n_28),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_139),
.A2(n_140),
.B1(n_152),
.B2(n_196),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_49),
.B1(n_21),
.B2(n_29),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_69),
.B(n_42),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_141),
.B(n_147),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_144),
.A2(n_147),
.B1(n_141),
.B2(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_40),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_150),
.B(n_151),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_59),
.B(n_29),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_106),
.A2(n_34),
.B1(n_38),
.B2(n_36),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_61),
.B(n_4),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_175),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_46),
.B1(n_38),
.B2(n_6),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_157),
.A2(n_194),
.B1(n_205),
.B2(n_202),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_4),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_165),
.B(n_171),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_4),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_90),
.A2(n_46),
.B(n_38),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_173),
.A2(n_184),
.B(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_68),
.B(n_5),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_5),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_176),
.B(n_186),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_71),
.B(n_46),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_179),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_117),
.A2(n_5),
.B(n_7),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_123),
.B(n_16),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_190),
.B(n_195),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_76),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_7),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_79),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_105),
.B(n_16),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_198),
.B(n_200),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_86),
.B(n_16),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_98),
.B(n_16),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_203),
.B(n_217),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_87),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_97),
.B(n_14),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_220),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_92),
.A2(n_14),
.B1(n_93),
.B2(n_94),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_169),
.B1(n_158),
.B2(n_170),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_95),
.B(n_14),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_69),
.B(n_65),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_222),
.A2(n_223),
.B1(n_254),
.B2(n_255),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_155),
.A2(n_209),
.B1(n_175),
.B2(n_154),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_149),
.B1(n_129),
.B2(n_214),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_224),
.A2(n_247),
.B1(n_259),
.B2(n_260),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_225),
.B(n_238),
.Y(n_308)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_246),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_227),
.A2(n_235),
.B(n_225),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_153),
.B1(n_204),
.B2(n_168),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_228),
.A2(n_237),
.B1(n_229),
.B2(n_274),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_202),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g328 ( 
.A1(n_229),
.A2(n_230),
.B(n_240),
.Y(n_328)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_160),
.B(n_132),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_179),
.A2(n_162),
.B1(n_174),
.B2(n_206),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_234),
.A2(n_243),
.B1(n_276),
.B2(n_280),
.Y(n_337)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_145),
.Y(n_236)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_236),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

BUFx4f_ASAP7_75t_SL g321 ( 
.A(n_239),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_131),
.B(n_161),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_241),
.Y(n_350)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_133),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_245),
.B(n_256),
.Y(n_312)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_212),
.B1(n_161),
.B2(n_131),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_248),
.B(n_249),
.Y(n_314)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_250),
.B(n_266),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_169),
.A2(n_188),
.B1(n_213),
.B2(n_143),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_179),
.A2(n_213),
.B(n_177),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_253),
.A2(n_229),
.B(n_273),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_138),
.A2(n_166),
.B1(n_182),
.B2(n_187),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_206),
.B1(n_168),
.B2(n_172),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_133),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_166),
.A2(n_182),
.B1(n_187),
.B2(n_143),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_130),
.A2(n_191),
.B1(n_135),
.B2(n_136),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_135),
.A2(n_136),
.B1(n_191),
.B2(n_167),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_261),
.A2(n_291),
.B1(n_298),
.B2(n_260),
.Y(n_326)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_145),
.Y(n_264)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_148),
.A2(n_172),
.B1(n_189),
.B2(n_180),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_265),
.A2(n_274),
.B1(n_281),
.B2(n_287),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_148),
.Y(n_267)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_180),
.B(n_189),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_297),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_134),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_159),
.Y(n_272)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_128),
.B(n_170),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_275),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_134),
.A2(n_218),
.B1(n_167),
.B2(n_183),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_156),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_218),
.A2(n_216),
.B1(n_193),
.B2(n_208),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_279),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_145),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_193),
.A2(n_216),
.B1(n_128),
.B2(n_164),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_193),
.A2(n_216),
.B1(n_164),
.B2(n_183),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_289),
.Y(n_342)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_193),
.A2(n_216),
.B1(n_146),
.B2(n_183),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_164),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_286),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_192),
.A2(n_140),
.B1(n_210),
.B2(n_139),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_192),
.A2(n_220),
.B(n_163),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_294),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_144),
.A2(n_151),
.B1(n_175),
.B2(n_155),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_130),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_292),
.Y(n_311)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_197),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_295),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_296),
.Y(n_318)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_144),
.A2(n_104),
.B1(n_181),
.B2(n_151),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_302),
.A2(n_330),
.B(n_304),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_253),
.B1(n_222),
.B2(n_269),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_304),
.A2(n_320),
.B1(n_344),
.B2(n_345),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_257),
.B(n_233),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_313),
.B(n_322),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_234),
.B1(n_296),
.B2(n_267),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_225),
.B(n_257),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_330),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_339),
.B1(n_341),
.B2(n_347),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_268),
.B(n_282),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_329),
.B(n_333),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_271),
.B(n_284),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_233),
.B(n_223),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_343),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_263),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_335),
.B(n_318),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_234),
.B(n_247),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

AOI32xp33_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_244),
.A3(n_227),
.B1(n_231),
.B2(n_221),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_342),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_234),
.A2(n_261),
.B1(n_231),
.B2(n_240),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_240),
.A2(n_292),
.B1(n_252),
.B2(n_258),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_272),
.B(n_297),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_255),
.A2(n_281),
.B1(n_294),
.B2(n_242),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_285),
.A2(n_295),
.B1(n_239),
.B2(n_241),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_285),
.A2(n_262),
.B1(n_278),
.B2(n_270),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_285),
.A2(n_266),
.B1(n_278),
.B2(n_286),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_309),
.B1(n_299),
.B2(n_327),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g349 ( 
.A(n_290),
.B(n_264),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_349),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_351),
.B(n_379),
.Y(n_415)
);

O2A1O1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_336),
.A2(n_275),
.B(n_283),
.C(n_236),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_353),
.A2(n_370),
.B(n_347),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_350),
.Y(n_355)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_362),
.Y(n_403)
);

AO22x1_ASAP7_75t_L g363 ( 
.A1(n_339),
.A2(n_309),
.B1(n_348),
.B2(n_336),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_371),
.Y(n_402)
);

XNOR2x2_ASAP7_75t_SL g364 ( 
.A(n_334),
.B(n_302),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_309),
.A2(n_320),
.B(n_319),
.Y(n_370)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_335),
.C(n_322),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_375),
.C(n_385),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_342),
.C(n_302),
.Y(n_375)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_376),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_306),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_377),
.B(n_383),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_329),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_SL g381 ( 
.A(n_319),
.B(n_338),
.C(n_309),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_381),
.Y(n_409)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_382),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_308),
.B(n_306),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_384),
.B(n_387),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_324),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_312),
.Y(n_386)
);

INVx13_ASAP7_75t_L g398 ( 
.A(n_386),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_326),
.A2(n_310),
.B1(n_327),
.B2(n_299),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_389),
.A2(n_310),
.B1(n_344),
.B2(n_341),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_314),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_390),
.B(n_391),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_312),
.B(n_316),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_314),
.B(n_346),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_392),
.B(n_332),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_396),
.A2(n_399),
.B1(n_360),
.B2(n_345),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_397),
.A2(n_370),
.B(n_399),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_366),
.A2(n_311),
.B1(n_337),
.B2(n_300),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_390),
.Y(n_400)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_346),
.C(n_303),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_417),
.C(n_375),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_332),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_355),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_422),
.Y(n_435)
);

INVx13_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_352),
.B(n_315),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_424),
.B(n_425),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_355),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_356),
.B(n_374),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_427),
.A2(n_423),
.B(n_416),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_428),
.B(n_434),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_430),
.A2(n_415),
.B(n_418),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_389),
.B1(n_363),
.B2(n_354),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_431),
.A2(n_436),
.B1(n_438),
.B2(n_440),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_364),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_433),
.B(n_451),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_356),
.C(n_365),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_402),
.A2(n_363),
.B1(n_407),
.B2(n_403),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_386),
.Y(n_437)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_371),
.B1(n_361),
.B2(n_354),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_383),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_439),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_402),
.A2(n_366),
.B1(n_361),
.B2(n_362),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_426),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_445),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_367),
.C(n_364),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_444),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_367),
.C(n_357),
.Y(n_444)
);

OAI32xp33_ASAP7_75t_L g445 ( 
.A1(n_395),
.A2(n_387),
.A3(n_377),
.B1(n_392),
.B2(n_351),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_446),
.A2(n_457),
.B1(n_393),
.B2(n_415),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_368),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_414),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_402),
.A2(n_360),
.B1(n_353),
.B2(n_337),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_448),
.A2(n_453),
.B1(n_397),
.B2(n_401),
.Y(n_467)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_369),
.Y(n_450)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_382),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_384),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_454),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_409),
.A2(n_337),
.B1(n_311),
.B2(n_305),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_398),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_414),
.B(n_305),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_418),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_398),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_425),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_337),
.B1(n_388),
.B2(n_340),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_458),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_464),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_440),
.A2(n_409),
.B1(n_406),
.B2(n_408),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_466),
.A2(n_432),
.B1(n_435),
.B2(n_442),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_467),
.A2(n_436),
.B1(n_427),
.B2(n_457),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_468),
.A2(n_470),
.B1(n_477),
.B2(n_478),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_424),
.Y(n_471)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_474),
.A2(n_481),
.B(n_486),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_422),
.Y(n_475)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_475),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_441),
.Y(n_476)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_476),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_438),
.A2(n_419),
.B1(n_398),
.B2(n_411),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_416),
.B1(n_423),
.B2(n_420),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_433),
.B(n_337),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_480),
.B(n_431),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_307),
.Y(n_483)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_483),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_450),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_455),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_453),
.A2(n_413),
.B1(n_412),
.B2(n_404),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_434),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_503),
.Y(n_514)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_489),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_490),
.B(n_497),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_496),
.B1(n_501),
.B2(n_507),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_462),
.B1(n_474),
.B2(n_477),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_432),
.B1(n_435),
.B2(n_442),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_482),
.B(n_443),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_482),
.B(n_451),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_499),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_428),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_471),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_476),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_466),
.A2(n_430),
.B1(n_445),
.B2(n_452),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_449),
.C(n_317),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_461),
.C(n_479),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_480),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_470),
.A2(n_429),
.B1(n_413),
.B2(n_412),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_429),
.Y(n_508)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_508),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_522),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_459),
.Y(n_510)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_510),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_512),
.A2(n_517),
.B1(n_524),
.B2(n_486),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_459),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_518),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_492),
.A2(n_469),
.B1(n_479),
.B2(n_467),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_488),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_487),
.B(n_481),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_521),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_508),
.C(n_504),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_501),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_478),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_461),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_515),
.A2(n_491),
.B(n_505),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_530),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_516),
.A2(n_495),
.B1(n_505),
.B2(n_494),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_528),
.A2(n_534),
.B1(n_473),
.B2(n_523),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_521),
.A2(n_520),
.B(n_519),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_513),
.A2(n_504),
.B(n_494),
.Y(n_531)
);

XOR2x2_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_404),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_522),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_533),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_511),
.A2(n_469),
.B1(n_490),
.B2(n_491),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_532),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_525),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_539),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_497),
.C(n_503),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_548),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_537),
.B(n_517),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_542),
.B(n_536),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_536),
.A2(n_464),
.B(n_525),
.Y(n_544)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_544),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_550),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_528),
.A2(n_523),
.B(n_473),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_546),
.A2(n_531),
.B(n_421),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_533),
.B(n_465),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_549),
.B(n_529),
.Y(n_552)
);

XOR2x2_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_498),
.Y(n_550)
);

OAI21xp33_ASAP7_75t_L g560 ( 
.A1(n_551),
.A2(n_552),
.B(n_547),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_538),
.C(n_539),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_553),
.B(n_555),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_527),
.Y(n_555)
);

AOI21x1_ASAP7_75t_SL g561 ( 
.A1(n_558),
.A2(n_546),
.B(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_562),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_557),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_548),
.C(n_545),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_556),
.B(n_550),
.C(n_465),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_557),
.C(n_554),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_388),
.C(n_340),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_559),
.B(n_465),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_567),
.A2(n_568),
.B(n_564),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_565),
.B(n_421),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_349),
.Y(n_571)
);


endmodule