module real_aes_7080_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g729 ( .A(n_0), .B(n_84), .C(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g489 ( .A(n_1), .Y(n_489) );
INVx1_ASAP7_75t_L g142 ( .A(n_2), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_3), .A2(n_37), .B1(n_167), .B2(n_445), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g186 ( .A1(n_4), .A2(n_158), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_5), .B(n_156), .Y(n_500) );
AND2x6_ASAP7_75t_L g135 ( .A(n_6), .B(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_38), .Y(n_112) );
INVx1_ASAP7_75t_L g192 ( .A(n_9), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_10), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g127 ( .A(n_11), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_12), .B(n_148), .Y(n_453) );
INVx1_ASAP7_75t_L g246 ( .A(n_13), .Y(n_246) );
INVx1_ASAP7_75t_L g483 ( .A(n_14), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_15), .B(n_123), .Y(n_505) );
AO32x2_ASAP7_75t_L g472 ( .A1(n_16), .A2(n_122), .A3(n_156), .B1(n_447), .B2(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_17), .B(n_167), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_18), .B(n_163), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_19), .B(n_123), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_20), .A2(n_49), .B1(n_167), .B2(n_445), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_21), .B(n_158), .Y(n_203) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_22), .A2(n_75), .B1(n_148), .B2(n_167), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_23), .B(n_167), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_24), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_25), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_26), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_27), .B(n_153), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_28), .B(n_146), .Y(n_145) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_29), .A2(n_100), .B1(n_725), .B2(n_733), .Y(n_99) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_30), .A2(n_115), .B1(n_714), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_30), .Y(n_723) );
INVx1_ASAP7_75t_L g181 ( .A(n_31), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_32), .B(n_153), .Y(n_470) );
INVx2_ASAP7_75t_L g133 ( .A(n_33), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_34), .B(n_167), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_35), .B(n_153), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_36), .A2(n_135), .B(n_138), .C(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g179 ( .A(n_39), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_40), .B(n_146), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_41), .B(n_167), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_42), .Y(n_106) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_43), .A2(n_85), .B1(n_210), .B2(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_44), .B(n_167), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_45), .B(n_167), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_46), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_47), .B(n_488), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_48), .B(n_158), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_50), .A2(n_59), .B1(n_148), .B2(n_167), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_51), .A2(n_138), .B1(n_148), .B2(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_52), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_53), .B(n_167), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_54), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_55), .B(n_167), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_56), .A2(n_166), .B(n_190), .C(n_191), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_57), .Y(n_237) );
INVx1_ASAP7_75t_L g188 ( .A(n_58), .Y(n_188) );
INVx1_ASAP7_75t_L g136 ( .A(n_60), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_61), .B(n_167), .Y(n_490) );
INVx1_ASAP7_75t_L g126 ( .A(n_62), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_63), .Y(n_104) );
AO32x2_ASAP7_75t_L g442 ( .A1(n_64), .A2(n_156), .A3(n_215), .B1(n_443), .B2(n_447), .Y(n_442) );
INVx1_ASAP7_75t_L g522 ( .A(n_65), .Y(n_522) );
INVx1_ASAP7_75t_L g465 ( .A(n_66), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g113 ( .A1(n_67), .A2(n_68), .B1(n_114), .B2(n_713), .C1(n_717), .C2(n_718), .Y(n_113) );
INVx1_ASAP7_75t_L g717 ( .A(n_68), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_SL g162 ( .A1(n_69), .A2(n_163), .B(n_164), .C(n_166), .Y(n_162) );
INVxp67_ASAP7_75t_L g165 ( .A(n_70), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_71), .B(n_148), .Y(n_466) );
INVx1_ASAP7_75t_L g732 ( .A(n_72), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_73), .Y(n_184) );
INVx1_ASAP7_75t_L g230 ( .A(n_74), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_76), .A2(n_135), .B(n_138), .C(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_77), .B(n_445), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_78), .B(n_148), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_79), .B(n_143), .Y(n_206) );
INVx2_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_81), .B(n_163), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_82), .B(n_148), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_83), .A2(n_135), .B(n_138), .C(n_141), .Y(n_137) );
OR2x2_ASAP7_75t_L g108 ( .A(n_84), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g434 ( .A(n_84), .B(n_110), .Y(n_434) );
INVx2_ASAP7_75t_L g712 ( .A(n_84), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_86), .A2(n_98), .B1(n_148), .B2(n_149), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_87), .B(n_153), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_88), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_89), .A2(n_135), .B(n_138), .C(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_90), .Y(n_225) );
INVx1_ASAP7_75t_L g161 ( .A(n_91), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_92), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_93), .B(n_143), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_94), .B(n_148), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_95), .B(n_156), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_96), .A2(n_158), .B(n_159), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_97), .B(n_732), .Y(n_731) );
AOI22x1_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_113), .B1(n_719), .B2(n_721), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g720 ( .A(n_103), .Y(n_720) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_105), .A2(n_722), .B(n_724), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_108), .Y(n_724) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_109), .B(n_712), .Y(n_718) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g711 ( .A(n_110), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x2_ASAP7_75t_L g727 ( .A(n_112), .B(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_432), .B1(n_435), .B2(n_709), .Y(n_114) );
INVx2_ASAP7_75t_L g714 ( .A(n_115), .Y(n_714) );
OR4x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_321), .C(n_381), .D(n_408), .Y(n_115) );
NAND4xp25_ASAP7_75t_SL g116 ( .A(n_117), .B(n_269), .C(n_300), .D(n_317), .Y(n_116) );
O2A1O1Ixp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_194), .B(n_196), .C(n_249), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_172), .Y(n_118) );
INVx1_ASAP7_75t_L g311 ( .A(n_119), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_119), .A2(n_352), .B1(n_400), .B2(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_154), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_120), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g262 ( .A(n_120), .B(n_174), .Y(n_262) );
AND2x2_ASAP7_75t_L g304 ( .A(n_120), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_120), .B(n_195), .Y(n_316) );
INVx1_ASAP7_75t_L g356 ( .A(n_120), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_120), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g284 ( .A(n_121), .B(n_174), .Y(n_284) );
INVx3_ASAP7_75t_L g288 ( .A(n_121), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_121), .B(n_346), .Y(n_345) );
AO21x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_128), .B(n_150), .Y(n_121) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_122), .A2(n_175), .B(n_183), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_122), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g211 ( .A(n_122), .Y(n_211) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_123), .Y(n_156) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_124), .B(n_125), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_137), .Y(n_128) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_130), .A2(n_168), .B1(n_176), .B2(n_182), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_130), .A2(n_230), .B(n_231), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
AND2x4_ASAP7_75t_L g158 ( .A(n_131), .B(n_135), .Y(n_158) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g488 ( .A(n_132), .Y(n_488) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx3_ASAP7_75t_L g144 ( .A(n_134), .Y(n_144) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_134), .Y(n_146) );
INVx1_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVx4_ASAP7_75t_SL g168 ( .A(n_135), .Y(n_168) );
BUFx3_ASAP7_75t_L g447 ( .A(n_135), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_135), .A2(n_451), .B(n_455), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_135), .A2(n_464), .B(n_467), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_135), .A2(n_482), .B(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_135), .A2(n_494), .B(n_497), .Y(n_493) );
INVx5_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
BUFx3_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
INVx1_ASAP7_75t_L g445 ( .A(n_139), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_145), .C(n_147), .Y(n_141) );
O2A1O1Ixp5_ASAP7_75t_SL g464 ( .A1(n_143), .A2(n_166), .B(n_465), .C(n_466), .Y(n_464) );
INVx2_ASAP7_75t_L g475 ( .A(n_143), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_143), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_143), .A2(n_519), .B(n_520), .Y(n_518) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_144), .B(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_144), .B(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_144), .A2(n_146), .B1(n_444), .B2(n_446), .Y(n_443) );
INVx2_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
INVx4_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_146), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_146), .A2(n_475), .B1(n_508), .B2(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_147), .A2(n_483), .B(n_484), .C(n_485), .Y(n_482) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_152), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_152), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_153), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_153), .A2(n_450), .B(n_458), .Y(n_449) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_153), .A2(n_463), .B(n_470), .Y(n_462) );
AND2x2_ASAP7_75t_L g375 ( .A(n_154), .B(n_185), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_154), .B(n_288), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_154), .B(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g195 ( .A(n_155), .B(n_174), .Y(n_195) );
INVx1_ASAP7_75t_L g257 ( .A(n_155), .Y(n_257) );
BUFx2_ASAP7_75t_L g261 ( .A(n_155), .Y(n_261) );
AND2x2_ASAP7_75t_L g305 ( .A(n_155), .B(n_173), .Y(n_305) );
OR2x2_ASAP7_75t_L g344 ( .A(n_155), .B(n_173), .Y(n_344) );
AND2x2_ASAP7_75t_L g369 ( .A(n_155), .B(n_185), .Y(n_369) );
AND2x2_ASAP7_75t_L g428 ( .A(n_155), .B(n_258), .Y(n_428) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_169), .Y(n_155) );
INVx4_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_156), .A2(n_493), .B(n_500), .Y(n_492) );
BUFx2_ASAP7_75t_L g240 ( .A(n_158), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_162), .C(n_168), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_160), .A2(n_168), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_160), .A2(n_168), .B(n_242), .C(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g454 ( .A(n_163), .Y(n_454) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_167), .Y(n_222) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_170), .A2(n_186), .B(n_193), .Y(n_185) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_171), .B(n_213), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_171), .B(n_447), .C(n_507), .Y(n_506) );
AO21x1_ASAP7_75t_L g553 ( .A1(n_171), .A2(n_507), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g403 ( .A(n_172), .Y(n_403) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_185), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_173), .B(n_185), .Y(n_289) );
AND2x2_ASAP7_75t_L g299 ( .A(n_173), .B(n_288), .Y(n_299) );
BUFx2_ASAP7_75t_L g310 ( .A(n_173), .Y(n_310) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g332 ( .A(n_174), .B(n_185), .Y(n_332) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_174), .Y(n_387) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_177) );
INVx2_ASAP7_75t_L g180 ( .A(n_178), .Y(n_180) );
INVx4_ASAP7_75t_L g244 ( .A(n_178), .Y(n_244) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_185), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_SL g258 ( .A(n_185), .Y(n_258) );
BUFx2_ASAP7_75t_L g283 ( .A(n_185), .Y(n_283) );
INVx2_ASAP7_75t_L g302 ( .A(n_185), .Y(n_302) );
AND2x2_ASAP7_75t_L g364 ( .A(n_185), .B(n_288), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_190), .A2(n_456), .B(n_457), .Y(n_455) );
O2A1O1Ixp5_ASAP7_75t_L g521 ( .A1(n_190), .A2(n_487), .B(n_522), .C(n_523), .Y(n_521) );
AOI321xp33_ASAP7_75t_L g383 ( .A1(n_194), .A2(n_384), .A3(n_385), .B1(n_386), .B2(n_388), .C(n_389), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_195), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_195), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g377 ( .A(n_195), .B(n_356), .Y(n_377) );
AND2x2_ASAP7_75t_L g410 ( .A(n_195), .B(n_302), .Y(n_410) );
INVx1_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_226), .Y(n_197) );
OR2x2_ASAP7_75t_L g312 ( .A(n_198), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g264 ( .A(n_201), .Y(n_264) );
AND2x2_ASAP7_75t_L g274 ( .A(n_201), .B(n_228), .Y(n_274) );
AND2x2_ASAP7_75t_L g279 ( .A(n_201), .B(n_254), .Y(n_279) );
INVx1_ASAP7_75t_L g296 ( .A(n_201), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_201), .B(n_277), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_201), .B(n_253), .Y(n_320) );
OR2x2_ASAP7_75t_L g352 ( .A(n_201), .B(n_341), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_201), .B(n_265), .Y(n_391) );
AND2x2_ASAP7_75t_L g425 ( .A(n_201), .B(n_251), .Y(n_425) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
AOI21xp5_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_204), .B(n_211), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_208), .A2(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g247 ( .A(n_210), .Y(n_247) );
INVx1_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_211), .A2(n_481), .B(n_491), .Y(n_480) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_211), .A2(n_517), .B(n_524), .Y(n_516) );
INVx1_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
INVx2_ASAP7_75t_L g267 ( .A(n_214), .Y(n_267) );
AND2x2_ASAP7_75t_L g307 ( .A(n_214), .B(n_278), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_214), .B(n_254), .Y(n_329) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_222), .Y(n_218) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g413 ( .A(n_227), .B(n_264), .Y(n_413) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_238), .Y(n_227) );
INVx2_ASAP7_75t_L g254 ( .A(n_228), .Y(n_254) );
AND2x2_ASAP7_75t_L g407 ( .A(n_228), .B(n_267), .Y(n_407) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_235), .B(n_236), .Y(n_228) );
AND2x2_ASAP7_75t_L g253 ( .A(n_238), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g268 ( .A(n_238), .Y(n_268) );
INVx1_ASAP7_75t_L g278 ( .A(n_238), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_244), .A2(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g485 ( .A(n_244), .Y(n_485) );
OAI22xp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_255), .B1(n_259), .B2(n_263), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_250), .A2(n_368), .B1(n_405), .B2(n_406), .Y(n_404) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_253), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g314 ( .A(n_254), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_254), .B(n_267), .Y(n_341) );
INVx1_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
AND2x2_ASAP7_75t_L g298 ( .A(n_256), .B(n_299), .Y(n_298) );
INVx3_ASAP7_75t_SL g337 ( .A(n_256), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_256), .B(n_262), .Y(n_414) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g423 ( .A(n_259), .Y(n_423) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_260), .B(n_356), .Y(n_398) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_SL g303 ( .A(n_262), .Y(n_303) );
NAND2x1_ASAP7_75t_SL g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x2_ASAP7_75t_L g324 ( .A(n_264), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g331 ( .A(n_264), .B(n_268), .Y(n_331) );
AND2x2_ASAP7_75t_L g336 ( .A(n_264), .B(n_277), .Y(n_336) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_264), .Y(n_385) );
OAI311xp33_ASAP7_75t_L g408 ( .A1(n_265), .A2(n_409), .A3(n_411), .B1(n_412), .C1(n_422), .Y(n_408) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g421 ( .A(n_266), .B(n_294), .Y(n_421) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g277 ( .A(n_267), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g325 ( .A(n_267), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g380 ( .A(n_267), .Y(n_380) );
INVx1_ASAP7_75t_L g273 ( .A(n_268), .Y(n_273) );
INVx1_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_268), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g326 ( .A(n_268), .Y(n_326) );
AOI221xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_272), .B1(n_280), .B2(n_285), .C(n_290), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx4_ASAP7_75t_L g294 ( .A(n_274), .Y(n_294) );
AND2x2_ASAP7_75t_L g388 ( .A(n_274), .B(n_307), .Y(n_388) );
AND2x2_ASAP7_75t_L g395 ( .A(n_274), .B(n_277), .Y(n_395) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_277), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g306 ( .A(n_279), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_282), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g431 ( .A(n_284), .B(n_375), .Y(n_431) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g416 ( .A(n_288), .B(n_344), .Y(n_416) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_289), .A2(n_382), .B(n_383), .C(n_396), .Y(n_381) );
AOI21xp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_295), .B(n_297), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_295), .A2(n_390), .B1(n_391), .B2(n_392), .C(n_393), .Y(n_389) );
AND2x2_ASAP7_75t_L g366 ( .A(n_296), .B(n_307), .Y(n_366) );
AND2x2_ASAP7_75t_L g419 ( .A(n_296), .B(n_314), .Y(n_419) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_299), .B(n_337), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B(n_306), .C(n_308), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g347 ( .A(n_302), .B(n_305), .Y(n_347) );
OR2x2_ASAP7_75t_L g390 ( .A(n_302), .B(n_344), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_303), .B(n_369), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_303), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g334 ( .A(n_304), .Y(n_334) );
INVx1_ASAP7_75t_L g400 ( .A(n_307), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_312), .B1(n_315), .B2(n_316), .Y(n_308) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_310), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g386 ( .A(n_311), .B(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g372 ( .A(n_313), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_314), .B(n_400), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_374), .B1(n_376), .B2(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g382 ( .A(n_318), .Y(n_382) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g424 ( .A(n_319), .B(n_419), .Y(n_424) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_320), .A2(n_354), .B1(n_357), .B2(n_358), .C1(n_361), .C2(n_362), .Y(n_353) );
NAND4xp25_ASAP7_75t_SL g321 ( .A(n_322), .B(n_342), .C(n_353), .D(n_365), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_327), .B2(n_332), .C(n_333), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_325), .B(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g351 ( .A(n_326), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_327), .A2(n_397), .B1(n_399), .B2(n_401), .C(n_404), .Y(n_396) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g339 ( .A(n_331), .B(n_340), .Y(n_339) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_332), .A2(n_394), .B(n_395), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_337), .B2(n_338), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B(n_348), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_356), .B(n_375), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_356), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_360), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g392 ( .A(n_364), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_370), .B2(n_372), .C(n_373), .Y(n_365) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI222xp33_ASAP7_75t_L g412 ( .A1(n_375), .A2(n_413), .B1(n_414), .B2(n_415), .C1(n_417), .C2(n_420), .Y(n_412) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_379), .B(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp33_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_425), .B2(n_426), .C(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_432), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g716 ( .A(n_435), .Y(n_716) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND3x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_629), .C(n_677), .Y(n_436) );
NOR4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_557), .C(n_602), .D(n_616), .Y(n_437) );
OAI311xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_477), .A3(n_501), .B1(n_510), .C1(n_525), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_448), .Y(n_439) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_440), .A2(n_511), .B(n_513), .Y(n_510) );
AND2x2_ASAP7_75t_L g618 ( .A(n_440), .B(n_545), .Y(n_618) );
AND2x2_ASAP7_75t_L g675 ( .A(n_440), .B(n_561), .Y(n_675) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g568 ( .A(n_441), .B(n_471), .Y(n_568) );
AND2x2_ASAP7_75t_L g625 ( .A(n_441), .B(n_573), .Y(n_625) );
INVx1_ASAP7_75t_L g666 ( .A(n_441), .Y(n_666) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_442), .Y(n_534) );
AND2x2_ASAP7_75t_L g575 ( .A(n_442), .B(n_471), .Y(n_575) );
AND2x2_ASAP7_75t_L g579 ( .A(n_442), .B(n_472), .Y(n_579) );
INVx1_ASAP7_75t_L g591 ( .A(n_442), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_447), .A2(n_518), .B(n_521), .Y(n_517) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_459), .Y(n_448) );
AND2x2_ASAP7_75t_L g512 ( .A(n_449), .B(n_471), .Y(n_512) );
INVx2_ASAP7_75t_L g546 ( .A(n_449), .Y(n_546) );
AND2x2_ASAP7_75t_L g561 ( .A(n_449), .B(n_472), .Y(n_561) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_449), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_449), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g581 ( .A(n_449), .B(n_544), .Y(n_581) );
INVx1_ASAP7_75t_L g593 ( .A(n_449), .Y(n_593) );
INVx1_ASAP7_75t_L g634 ( .A(n_449), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_449), .B(n_534), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_454), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g511 ( .A(n_461), .B(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_461), .B(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g596 ( .A(n_461), .B(n_471), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_461), .B(n_591), .Y(n_654) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g544 ( .A(n_462), .Y(n_544) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_462), .Y(n_560) );
OR2x2_ASAP7_75t_L g633 ( .A(n_462), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
AND2x2_ASAP7_75t_L g545 ( .A(n_472), .B(n_546), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_475), .A2(n_487), .B(n_489), .C(n_490), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_475), .A2(n_498), .B(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_477), .B(n_528), .Y(n_691) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g661 ( .A(n_478), .B(n_503), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_492), .Y(n_478) );
AND2x2_ASAP7_75t_L g537 ( .A(n_479), .B(n_528), .Y(n_537) );
INVx2_ASAP7_75t_L g549 ( .A(n_479), .Y(n_549) );
AND2x2_ASAP7_75t_L g583 ( .A(n_479), .B(n_531), .Y(n_583) );
AND2x2_ASAP7_75t_L g650 ( .A(n_479), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_480), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g530 ( .A(n_480), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g570 ( .A(n_480), .B(n_492), .Y(n_570) );
AND2x2_ASAP7_75t_L g587 ( .A(n_480), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g513 ( .A(n_492), .B(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g531 ( .A(n_492), .Y(n_531) );
AND2x2_ASAP7_75t_L g536 ( .A(n_492), .B(n_516), .Y(n_536) );
AND2x2_ASAP7_75t_L g609 ( .A(n_492), .B(n_588), .Y(n_609) );
AND2x2_ASAP7_75t_L g674 ( .A(n_492), .B(n_664), .Y(n_674) );
OAI311xp33_ASAP7_75t_L g557 ( .A1(n_501), .A2(n_558), .A3(n_562), .B1(n_564), .C1(n_584), .Y(n_557) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g628 ( .A(n_502), .B(n_536), .Y(n_628) );
AND2x2_ASAP7_75t_L g702 ( .A(n_502), .B(n_583), .Y(n_702) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_503), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g637 ( .A(n_503), .Y(n_637) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g528 ( .A(n_504), .Y(n_528) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_504), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g657 ( .A(n_504), .B(n_531), .Y(n_657) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
AND2x2_ASAP7_75t_L g532 ( .A(n_512), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g585 ( .A(n_512), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g665 ( .A(n_512), .B(n_666), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_513), .A2(n_545), .B1(n_565), .B2(n_569), .C(n_571), .Y(n_564) );
INVx1_ASAP7_75t_L g689 ( .A(n_514), .Y(n_689) );
OR2x2_ASAP7_75t_L g655 ( .A(n_515), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g550 ( .A(n_516), .B(n_531), .Y(n_550) );
OR2x2_ASAP7_75t_L g552 ( .A(n_516), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
INVx2_ASAP7_75t_L g588 ( .A(n_516), .Y(n_588) );
AND2x2_ASAP7_75t_L g615 ( .A(n_516), .B(n_553), .Y(n_615) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_516), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_532), .B1(n_535), .B2(n_538), .C(n_541), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g626 ( .A(n_528), .B(n_536), .Y(n_626) );
AND2x2_ASAP7_75t_L g676 ( .A(n_528), .B(n_530), .Y(n_676) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g563 ( .A(n_530), .B(n_534), .Y(n_563) );
AND2x2_ASAP7_75t_L g642 ( .A(n_530), .B(n_615), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_531), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g601 ( .A(n_531), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_532), .A2(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g555 ( .A(n_533), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g621 ( .A(n_533), .B(n_581), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_533), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g598 ( .A(n_534), .B(n_567), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_534), .B(n_681), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_535), .B(n_561), .Y(n_671) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_L g594 ( .A(n_536), .B(n_549), .Y(n_594) );
INVx1_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_547), .B1(n_551), .B2(n_555), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g573 ( .A(n_544), .Y(n_573) );
INVx1_ASAP7_75t_L g586 ( .A(n_544), .Y(n_586) );
INVx1_ASAP7_75t_L g556 ( .A(n_545), .Y(n_556) );
AND2x2_ASAP7_75t_L g627 ( .A(n_545), .B(n_573), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_545), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
OR2x2_ASAP7_75t_L g551 ( .A(n_548), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_548), .B(n_664), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g695 ( .A(n_548), .B(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g698 ( .A(n_550), .B(n_650), .Y(n_698) );
INVx1_ASAP7_75t_SL g664 ( .A(n_552), .Y(n_664) );
AND2x2_ASAP7_75t_L g604 ( .A(n_553), .B(n_588), .Y(n_604) );
INVx1_ASAP7_75t_L g651 ( .A(n_553), .Y(n_651) );
OAI222xp33_ASAP7_75t_L g692 ( .A1(n_558), .A2(n_648), .B1(n_693), .B2(n_694), .C1(n_697), .C2(n_699), .Y(n_692) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g613 ( .A(n_560), .Y(n_613) );
AND2x2_ASAP7_75t_L g624 ( .A(n_561), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_561), .B(n_666), .Y(n_693) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_563), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g668 ( .A(n_565), .Y(n_668) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_SL g606 ( .A(n_568), .Y(n_606) );
AND2x2_ASAP7_75t_L g685 ( .A(n_568), .B(n_646), .Y(n_685) );
AND2x2_ASAP7_75t_L g708 ( .A(n_568), .B(n_592), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_570), .B(n_604), .Y(n_603) );
OAI32xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .A3(n_576), .B1(n_578), .B2(n_582), .Y(n_571) );
BUFx2_ASAP7_75t_L g646 ( .A(n_573), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_574), .B(n_592), .Y(n_673) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g612 ( .A(n_575), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g680 ( .A(n_575), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g669 ( .A(n_576), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x2_ASAP7_75t_L g640 ( .A(n_579), .B(n_613), .Y(n_640) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OAI221xp5_ASAP7_75t_SL g602 ( .A1(n_581), .A2(n_603), .B1(n_605), .B2(n_607), .C(n_611), .Y(n_602) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g614 ( .A(n_583), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_583), .B(n_604), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B1(n_589), .B2(n_594), .C(n_595), .Y(n_584) );
INVx1_ASAP7_75t_L g703 ( .A(n_585), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_586), .B(n_680), .Y(n_679) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_587), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_592), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g658 ( .A(n_592), .Y(n_658) );
BUFx3_ASAP7_75t_L g681 ( .A(n_593), .Y(n_681) );
INVx1_ASAP7_75t_SL g622 ( .A(n_594), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_594), .B(n_636), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B(n_599), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_596), .A2(n_697), .B1(n_701), .B2(n_703), .C(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g643 ( .A(n_601), .B(n_604), .Y(n_643) );
INVx1_ASAP7_75t_L g707 ( .A(n_601), .Y(n_707) );
INVx2_ASAP7_75t_L g696 ( .A(n_604), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_604), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g649 ( .A(n_609), .B(n_650), .Y(n_649) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_619), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_625), .A2(n_687), .B1(n_688), .B2(n_690), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_628), .A2(n_705), .B(n_708), .Y(n_704) );
NOR4xp25_ASAP7_75t_SL g629 ( .A(n_630), .B(n_638), .C(n_647), .D(n_667), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_644), .B2(n_645), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g683 ( .A(n_643), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_652), .B1(n_655), .B2(n_658), .C(n_659), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g670 ( .A(n_650), .Y(n_670) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_662), .B(n_665), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_671), .C(n_672), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_672) );
CKINVDCx14_ASAP7_75t_R g682 ( .A(n_676), .Y(n_682) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_692), .C(n_700), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B1(n_683), .B2(n_684), .C(n_686), .Y(n_678) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx16_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g715 ( .A(n_710), .Y(n_715) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx12_ASAP7_75t_R g735 ( .A(n_727), .Y(n_735) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
endmodule