module fake_jpeg_12523_n_563 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_563);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_563;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_62),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_75),
.Y(n_129)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_69),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_74),
.B(n_76),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_27),
.B(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_13),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_79),
.Y(n_183)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_84),
.Y(n_135)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_87),
.Y(n_181)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_51),
.Y(n_90)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_26),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_94),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_39),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_96),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_19),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_22),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_118),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_114),
.Y(n_145)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_31),
.B(n_1),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_120),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_121),
.Y(n_173)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_41),
.B(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_123),
.B(n_125),
.Y(n_191)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_58),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_22),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_57),
.B1(n_46),
.B2(n_55),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_127),
.A2(n_134),
.B1(n_139),
.B2(n_152),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_25),
.B1(n_55),
.B2(n_46),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_131),
.A2(n_154),
.B1(n_158),
.B2(n_161),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_42),
.B1(n_51),
.B2(n_40),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_25),
.B1(n_55),
.B2(n_40),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_137),
.B(n_177),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_67),
.A2(n_42),
.B1(n_32),
.B2(n_57),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_49),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_146),
.B(n_128),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_64),
.B(n_37),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_148),
.B(n_151),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_31),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_65),
.A2(n_57),
.B1(n_37),
.B2(n_54),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_73),
.B(n_54),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_153),
.B(n_159),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_66),
.A2(n_50),
.B1(n_44),
.B2(n_32),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_68),
.A2(n_59),
.B1(n_53),
.B2(n_41),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_50),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_71),
.A2(n_44),
.B1(n_53),
.B2(n_59),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_67),
.A2(n_49),
.B1(n_58),
.B2(n_6),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_169),
.A2(n_187),
.B1(n_117),
.B2(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_174),
.B(n_193),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_79),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_176),
.A2(n_128),
.B1(n_141),
.B2(n_126),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_62),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_62),
.A2(n_3),
.B(n_8),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_179),
.B(n_192),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_94),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_182),
.A2(n_197),
.B1(n_187),
.B2(n_134),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_117),
.A2(n_11),
.B1(n_12),
.B2(n_124),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_86),
.B(n_12),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_89),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_101),
.A2(n_12),
.B1(n_122),
.B2(n_106),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_78),
.B(n_81),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_198),
.B(n_199),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_205),
.A2(n_222),
.B1(n_249),
.B2(n_239),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_100),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_206),
.B(n_215),
.Y(n_282)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_147),
.A2(n_104),
.B1(n_97),
.B2(n_115),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_208),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_245),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_212),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_108),
.B1(n_97),
.B2(n_110),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_213),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_214),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_132),
.B(n_102),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_129),
.B(n_108),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_217),
.B(n_235),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_103),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_219),
.B(n_224),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_139),
.A2(n_69),
.B1(n_109),
.B2(n_110),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_220),
.A2(n_252),
.B1(n_253),
.B2(n_238),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_149),
.B(n_115),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_221),
.B(n_272),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_168),
.B1(n_162),
.B2(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

BUFx12_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_145),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_229),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_146),
.B(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_136),
.B(n_155),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_230),
.B(n_237),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_231),
.B(n_234),
.Y(n_284)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_233),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_166),
.B(n_171),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_142),
.B(n_140),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_272),
.B1(n_209),
.B2(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_172),
.B(n_135),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_238),
.A2(n_234),
.B1(n_273),
.B2(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_168),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_266),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_202),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_240),
.B(n_243),
.Y(n_309)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_170),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_246),
.B(n_257),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_262),
.Y(n_299)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_190),
.A2(n_170),
.B1(n_178),
.B2(n_138),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_126),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_255),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_127),
.A2(n_169),
.B1(n_197),
.B2(n_195),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_133),
.B(n_175),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_138),
.B(n_178),
.Y(n_257)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_144),
.Y(n_260)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_181),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_144),
.B(n_195),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_269),
.Y(n_328)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_180),
.Y(n_264)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_130),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_265),
.B(n_270),
.Y(n_324)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_164),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_271),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_221),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_167),
.B(n_175),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_167),
.B(n_183),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_183),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_186),
.B(n_188),
.Y(n_272)
);

OR2x4_ASAP7_75t_L g273 ( 
.A(n_186),
.B(n_188),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.Y(n_289)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_185),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_275),
.A2(n_285),
.B1(n_295),
.B2(n_271),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_206),
.C(n_231),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_288),
.C(n_292),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_231),
.A2(n_209),
.B(n_229),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_326),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_218),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_283),
.B(n_313),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_258),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_241),
.C(n_210),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_225),
.C(n_234),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_293),
.A2(n_301),
.B1(n_254),
.B2(n_267),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_226),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_310),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_269),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_304),
.Y(n_370)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_227),
.A2(n_274),
.A3(n_223),
.B1(n_237),
.B2(n_216),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_211),
.B(n_262),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_207),
.B(n_261),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_314),
.B(n_299),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_242),
.A2(n_244),
.B1(n_248),
.B2(n_232),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_321),
.A2(n_322),
.B(n_278),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_233),
.B(n_268),
.C(n_247),
.Y(n_326)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_331),
.A2(n_336),
.B1(n_349),
.B2(n_358),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_266),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_339),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_334),
.B(n_354),
.Y(n_379)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_293),
.A2(n_260),
.B1(n_251),
.B2(n_256),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_327),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_347),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_212),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_289),
.A2(n_226),
.B(n_212),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_363),
.B(n_322),
.Y(n_375)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_343),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_212),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_344),
.B(n_348),
.Y(n_382)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_327),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_316),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_301),
.A2(n_323),
.B1(n_285),
.B2(n_289),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_312),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_352),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_295),
.A2(n_323),
.B1(n_291),
.B2(n_328),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_351),
.A2(n_307),
.B1(n_287),
.B2(n_311),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_327),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_290),
.A2(n_329),
.B1(n_284),
.B2(n_324),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_353),
.A2(n_367),
.B(n_325),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_291),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_277),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_356),
.B(n_357),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_310),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_286),
.A2(n_298),
.B1(n_288),
.B2(n_283),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_364),
.Y(n_395)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_284),
.A2(n_290),
.B1(n_329),
.B2(n_312),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_361),
.Y(n_381)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

AO22x2_ASAP7_75t_L g365 ( 
.A1(n_284),
.A2(n_292),
.B1(n_300),
.B2(n_303),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_366),
.Y(n_388)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_298),
.A2(n_279),
.B1(n_326),
.B2(n_306),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_305),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_368),
.Y(n_373)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_281),
.A2(n_318),
.B1(n_305),
.B2(n_307),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_371),
.A2(n_315),
.B1(n_320),
.B2(n_306),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_294),
.C(n_318),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_383),
.C(n_385),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_375),
.A2(n_400),
.B(n_350),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_391),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_311),
.C(n_287),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_356),
.B(n_280),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_385),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_308),
.C(n_315),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_280),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_407),
.C(n_347),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_371),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_345),
.B(n_320),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_396),
.B(n_397),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_280),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_332),
.A2(n_325),
.B(n_280),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_398),
.A2(n_362),
.B(n_330),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_349),
.A2(n_336),
.B1(n_357),
.B2(n_333),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_365),
.B1(n_364),
.B2(n_360),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_353),
.A2(n_367),
.B(n_340),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_363),
.B(n_365),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_351),
.B(n_334),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_382),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_409),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_395),
.Y(n_409)
);

INVx3_ASAP7_75t_SL g410 ( 
.A(n_388),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_414),
.Y(n_451)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_382),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_411),
.A2(n_420),
.B1(n_429),
.B2(n_432),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_339),
.Y(n_413)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_374),
.B(n_404),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_394),
.Y(n_416)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_422),
.Y(n_458)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_394),
.Y(n_418)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_340),
.B1(n_370),
.B2(n_337),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_342),
.C(n_346),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_343),
.Y(n_423)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_430),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_425),
.B(n_435),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_372),
.B(n_365),
.C(n_369),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_431),
.C(n_437),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_428),
.A2(n_434),
.B1(n_388),
.B2(n_376),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_365),
.C(n_366),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_407),
.A2(n_335),
.B1(n_368),
.B2(n_388),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_390),
.A2(n_379),
.B1(n_374),
.B2(n_381),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_383),
.B(n_384),
.C(n_407),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_438),
.A2(n_457),
.B1(n_459),
.B2(n_417),
.Y(n_482)
);

OA22x2_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_381),
.B1(n_390),
.B2(n_391),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_420),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_384),
.C(n_400),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_454),
.C(n_456),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_379),
.B1(n_387),
.B2(n_375),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_453),
.B1(n_414),
.B2(n_410),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_410),
.A2(n_387),
.B1(n_386),
.B2(n_398),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_405),
.C(n_386),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_377),
.C(n_389),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_434),
.A2(n_397),
.B1(n_396),
.B2(n_402),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_414),
.A2(n_402),
.B1(n_406),
.B2(n_373),
.Y(n_459)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_421),
.Y(n_461)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_406),
.C(n_378),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_429),
.C(n_423),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_435),
.B(n_425),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_464),
.B(n_431),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_468),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_409),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_466),
.B(n_487),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_428),
.Y(n_468)
);

XOR2x1_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_470),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_460),
.A2(n_419),
.B1(n_412),
.B2(n_413),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_438),
.B1(n_457),
.B2(n_459),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_436),
.Y(n_472)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_483),
.C(n_485),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_443),
.Y(n_474)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_450),
.B(n_423),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_480),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_458),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_481),
.Y(n_503)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_479),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_450),
.B(n_426),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_439),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_449),
.B1(n_447),
.B2(n_446),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_464),
.C(n_454),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_484),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_424),
.C(n_378),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_412),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_486),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_380),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_488),
.A2(n_486),
.B1(n_452),
.B2(n_433),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_485),
.A2(n_451),
.B(n_448),
.Y(n_491)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_465),
.C(n_480),
.Y(n_515)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_470),
.A2(n_451),
.B(n_442),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_494),
.A2(n_469),
.B(n_471),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_447),
.C(n_453),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_504),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_476),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_478),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_446),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_482),
.A2(n_446),
.B1(n_452),
.B2(n_455),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_505),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_521),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_503),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_512),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_510),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_472),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_474),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_514),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_501),
.B(n_467),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_517),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_493),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_467),
.C(n_473),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g531 ( 
.A(n_518),
.B(n_520),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_519),
.A2(n_505),
.B1(n_499),
.B2(n_495),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_475),
.C(n_418),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_497),
.Y(n_521)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_518),
.Y(n_525)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_504),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_526),
.B(n_528),
.Y(n_536)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_527),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_488),
.Y(n_528)
);

XNOR2x1_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_496),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_498),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_489),
.C(n_495),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_532),
.B(n_489),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_507),
.Y(n_535)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_535),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_524),
.A2(n_512),
.B(n_521),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_494),
.B(n_510),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_539),
.Y(n_547)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_523),
.A2(n_519),
.B(n_516),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_542),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_498),
.Y(n_542)
);

NAND2xp67_ASAP7_75t_SL g543 ( 
.A(n_529),
.B(n_533),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_543),
.B(n_524),
.Y(n_548)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_544),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_536),
.B(n_525),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_545),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_548),
.A2(n_539),
.B(n_531),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_493),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_527),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_535),
.C(n_540),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_551),
.A2(n_538),
.B(n_547),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_553),
.A2(n_555),
.B(n_537),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_556),
.B(n_557),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_552),
.B(n_546),
.C(n_549),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_558),
.B(n_554),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_560),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_559),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_562),
.A2(n_532),
.B(n_502),
.Y(n_563)
);


endmodule