module fake_jpeg_31070_n_412 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_412);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_46),
.Y(n_90)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_81),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_58),
.Y(n_108)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_19),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_70),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_11),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_75),
.Y(n_118)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_39),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_25),
.B(n_11),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_123),
.Y(n_145)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_30),
.B1(n_23),
.B2(n_41),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_96),
.B1(n_103),
.B2(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_38),
.B1(n_32),
.B2(n_43),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_43),
.B1(n_27),
.B2(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_99),
.B1(n_114),
.B2(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_43),
.B1(n_27),
.B2(n_39),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_27),
.B1(n_40),
.B2(n_28),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_42),
.B1(n_35),
.B2(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_113),
.B1(n_122),
.B2(n_52),
.Y(n_130)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_61),
.A2(n_22),
.B1(n_40),
.B2(n_28),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_54),
.A2(n_39),
.B1(n_24),
.B2(n_20),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_42),
.B1(n_35),
.B2(n_33),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_44),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_71),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_79),
.B1(n_65),
.B2(n_63),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_129),
.B(n_142),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_130),
.B(n_131),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_78),
.B1(n_80),
.B2(n_60),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_136),
.A2(n_139),
.B1(n_157),
.B2(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_82),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_146),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_80),
.B1(n_78),
.B2(n_70),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_47),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_46),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_55),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_155),
.Y(n_176)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_91),
.B(n_74),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_92),
.Y(n_205)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_66),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_124),
.B1(n_116),
.B2(n_119),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_1),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_167),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_53),
.B1(n_45),
.B2(n_51),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_69),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_161),
.Y(n_182)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_93),
.A2(n_69),
.B1(n_51),
.B2(n_74),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_164),
.Y(n_202)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_87),
.B(n_74),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_1),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_88),
.B(n_2),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_171),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_5),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_101),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_111),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_124),
.B1(n_116),
.B2(n_101),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_154),
.B1(n_157),
.B2(n_130),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_120),
.B(n_121),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_178),
.A2(n_135),
.B(n_137),
.Y(n_223)
);

BUFx16f_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_115),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_194),
.B(n_213),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_167),
.B1(n_144),
.B2(n_174),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_187),
.B(n_197),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_192),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_115),
.B(n_83),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_131),
.B(n_110),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_204),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_151),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_7),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_146),
.B(n_92),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_133),
.A2(n_126),
.B1(n_110),
.B2(n_119),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_8),
.B1(n_211),
.B2(n_195),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_141),
.A2(n_111),
.B1(n_105),
.B2(n_84),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_9),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_171),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_228),
.B1(n_243),
.B2(n_210),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_133),
.B1(n_163),
.B2(n_150),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_223),
.B(n_240),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_225),
.A2(n_237),
.B1(n_238),
.B2(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_227),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_149),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_159),
.B1(n_168),
.B2(n_152),
.Y(n_228)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_166),
.B(n_164),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_134),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_233),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_134),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_234),
.B(n_235),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_179),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_158),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_242),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_140),
.B1(n_161),
.B2(n_9),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_7),
.B1(n_8),
.B2(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_197),
.B(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_244),
.B(n_245),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_180),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_246),
.B(n_247),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_188),
.B(n_180),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_208),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_212),
.B1(n_194),
.B2(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_205),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_204),
.C(n_178),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_259),
.C(n_260),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_210),
.B(n_202),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_256),
.A2(n_263),
.B(n_264),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_257),
.A2(n_277),
.B1(n_285),
.B2(n_237),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_184),
.C(n_215),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_184),
.C(n_182),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_201),
.B(n_183),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_217),
.A2(n_201),
.B(n_179),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_212),
.C(n_176),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_284),
.C(n_222),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_218),
.A2(n_190),
.B(n_209),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_276),
.B(n_285),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_195),
.B1(n_181),
.B2(n_192),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_281),
.B1(n_219),
.B2(n_231),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_200),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_273),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_236),
.A2(n_181),
.B(n_200),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_221),
.A2(n_186),
.B1(n_181),
.B2(n_189),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_220),
.B(n_193),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_278),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_243),
.A2(n_186),
.B1(n_189),
.B2(n_193),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_233),
.C(n_248),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_219),
.A2(n_243),
.B1(n_245),
.B2(n_234),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_217),
.B1(n_252),
.B2(n_241),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_290),
.A2(n_295),
.B1(n_306),
.B2(n_277),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_220),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_244),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_299),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_242),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_243),
.B1(n_222),
.B2(n_230),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_262),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_267),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_300),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_301),
.A2(n_281),
.B1(n_274),
.B2(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_223),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_283),
.C(n_254),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_305),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_222),
.B1(n_230),
.B2(n_232),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_256),
.Y(n_316)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_311),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_313),
.B(n_264),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_310),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_224),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_238),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_280),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_255),
.B(n_230),
.C(n_249),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_329),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_324),
.C(n_330),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_320),
.A2(n_329),
.B(n_296),
.Y(n_349)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_295),
.A2(n_255),
.A3(n_258),
.B1(n_280),
.B2(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_284),
.C(n_260),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_301),
.B1(n_287),
.B2(n_290),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_293),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_263),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_265),
.C(n_276),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_271),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_334),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_271),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_335),
.A2(n_306),
.B1(n_298),
.B2(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_323),
.B(n_305),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_322),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_320),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

BUFx12f_ASAP7_75t_SL g342 ( 
.A(n_314),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_354),
.B1(n_335),
.B2(n_334),
.Y(n_362)
);

A2O1A1O1Ixp25_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_327),
.B(n_318),
.C(n_299),
.D(n_319),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_311),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_328),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_346),
.B(n_350),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_314),
.A2(n_298),
.B1(n_304),
.B2(n_287),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_347),
.A2(n_355),
.B1(n_332),
.B2(n_325),
.Y(n_361)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_351),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_319),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_296),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_317),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_352),
.B(n_336),
.Y(n_368)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_333),
.C(n_324),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_356),
.B(n_357),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_330),
.C(n_315),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_364),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_312),
.C(n_332),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_292),
.B1(n_294),
.B2(n_326),
.Y(n_366)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_355),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_310),
.C(n_304),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_342),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_373),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_369),
.B(n_341),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_382),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_359),
.A2(n_339),
.B(n_349),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_378),
.A2(n_358),
.B(n_338),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_343),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_340),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_359),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_384),
.B(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_380),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_387),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_365),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_379),
.A2(n_358),
.B(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_331),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_390),
.B(n_391),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_376),
.A2(n_367),
.B(n_364),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_282),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_373),
.C(n_376),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_395),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_372),
.C(n_378),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_388),
.A2(n_345),
.B1(n_351),
.B2(n_297),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_396),
.B(n_398),
.Y(n_402)
);

A2O1A1O1Ixp25_ASAP7_75t_L g397 ( 
.A1(n_384),
.A2(n_367),
.B(n_308),
.C(n_302),
.D(n_288),
.Y(n_397)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_397),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_403),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_269),
.C(n_250),
.Y(n_403)
);

AOI321xp33_ASAP7_75t_L g407 ( 
.A1(n_405),
.A2(n_400),
.A3(n_394),
.B1(n_395),
.B2(n_397),
.C(n_398),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_407),
.B(n_408),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_404),
.A2(n_229),
.B(n_225),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_406),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_409),
.B(n_402),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_410),
.Y(n_412)
);


endmodule