module real_aes_8263_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_0), .A2(n_145), .B(n_466), .C(n_469), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_1), .B(n_460), .Y(n_471) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g183 ( .A(n_3), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_4), .B(n_146), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_5), .A2(n_124), .B1(n_125), .B2(n_431), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_5), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_5), .A2(n_95), .B1(n_431), .B2(n_735), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_6), .A2(n_445), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_7), .A2(n_152), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_8), .A2(n_36), .B1(n_149), .B2(n_201), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_9), .B(n_152), .Y(n_169) );
AND2x6_ASAP7_75t_L g154 ( .A(n_10), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_11), .A2(n_154), .B(n_448), .C(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_12), .B(n_38), .Y(n_115) );
INVx1_ASAP7_75t_L g136 ( .A(n_13), .Y(n_136) );
INVx1_ASAP7_75t_L g175 ( .A(n_14), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_15), .B(n_142), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_16), .B(n_146), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_17), .B(n_132), .Y(n_131) );
AO32x2_ASAP7_75t_L g212 ( .A1(n_18), .A2(n_152), .A3(n_153), .B1(n_172), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_19), .B(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_20), .B(n_132), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_21), .A2(n_54), .B1(n_149), .B2(n_201), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g209 ( .A1(n_22), .A2(n_80), .B1(n_142), .B2(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_23), .B(n_149), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_24), .A2(n_153), .B(n_448), .C(n_450), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_25), .A2(n_153), .B(n_448), .C(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_27), .A2(n_96), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_27), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_28), .B(n_191), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_29), .A2(n_445), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_30), .B(n_191), .Y(n_228) );
INVx2_ASAP7_75t_L g144 ( .A(n_31), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_32), .A2(n_480), .B(n_481), .C(n_485), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_33), .B(n_149), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_34), .B(n_191), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_35), .B(n_197), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_37), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_39), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_40), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_41), .B(n_146), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_42), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_43), .B(n_445), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_44), .A2(n_480), .B(n_485), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_45), .B(n_149), .Y(n_162) );
INVx1_ASAP7_75t_L g467 ( .A(n_46), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_47), .A2(n_733), .B1(n_736), .B2(n_737), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_47), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_48), .A2(n_89), .B1(n_201), .B2(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g506 ( .A(n_49), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_50), .B(n_149), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_51), .B(n_149), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_52), .B(n_445), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_53), .B(n_167), .Y(n_166) );
AOI22xp33_ASAP7_75t_SL g148 ( .A1(n_55), .A2(n_59), .B1(n_142), .B2(n_149), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_56), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_57), .B(n_149), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_58), .B(n_149), .Y(n_248) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_61), .B(n_445), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_62), .B(n_460), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_63), .A2(n_167), .B(n_178), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_64), .B(n_149), .Y(n_184) );
INVx1_ASAP7_75t_L g135 ( .A(n_65), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_66), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_67), .B(n_146), .Y(n_483) );
AO32x2_ASAP7_75t_L g205 ( .A1(n_68), .A2(n_152), .A3(n_153), .B1(n_206), .B2(n_210), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_69), .B(n_147), .Y(n_517) );
INVx1_ASAP7_75t_L g247 ( .A(n_70), .Y(n_247) );
INVx1_ASAP7_75t_L g223 ( .A(n_71), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_72), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_73), .A2(n_103), .B1(n_116), .B2(n_744), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_74), .B(n_452), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_75), .A2(n_448), .B(n_485), .C(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_76), .B(n_142), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_77), .Y(n_493) );
INVx1_ASAP7_75t_L g108 ( .A(n_78), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_79), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_81), .B(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_82), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_83), .B(n_142), .Y(n_227) );
INVx2_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_85), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_86), .B(n_139), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_87), .B(n_142), .Y(n_163) );
INVx2_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
OR2x2_ASAP7_75t_L g434 ( .A(n_88), .B(n_113), .Y(n_434) );
OR2x2_ASAP7_75t_L g731 ( .A(n_88), .B(n_112), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_90), .A2(n_101), .B1(n_142), .B2(n_143), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_91), .B(n_445), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_92), .Y(n_482) );
INVxp67_ASAP7_75t_L g496 ( .A(n_93), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_94), .B(n_142), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_95), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_96), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_97), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g513 ( .A(n_98), .Y(n_513) );
INVx1_ASAP7_75t_L g542 ( .A(n_99), .Y(n_542) );
AND2x2_ASAP7_75t_L g508 ( .A(n_100), .B(n_191), .Y(n_508) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx12_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g745 ( .A(n_106), .Y(n_745) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g725 ( .A(n_110), .Y(n_725) );
NOR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g719 ( .A(n_111), .B(n_113), .Y(n_719) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AO221x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_726), .B1(n_729), .B2(n_738), .C(n_740), .Y(n_116) );
OAI222xp33_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_121), .B1(n_720), .B2(n_721), .C1(n_724), .C2(n_725), .Y(n_117) );
INVx1_ASAP7_75t_L g720 ( .A(n_118), .Y(n_720) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_432), .B1(n_435), .B2(n_717), .Y(n_122) );
INVx1_ASAP7_75t_L g723 ( .A(n_123), .Y(n_723) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g733 ( .A(n_125), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_365), .Y(n_125) );
NOR5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_278), .C(n_324), .D(n_337), .E(n_349), .Y(n_126) );
OAI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_186), .B(n_232), .C(n_259), .Y(n_127) );
INVx1_ASAP7_75t_SL g360 ( .A(n_128), .Y(n_360) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_156), .Y(n_128) );
AND2x2_ASAP7_75t_L g284 ( .A(n_129), .B(n_157), .Y(n_284) );
AND2x2_ASAP7_75t_L g312 ( .A(n_129), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_129), .B(n_263), .Y(n_320) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g250 ( .A(n_130), .B(n_158), .Y(n_250) );
INVx2_ASAP7_75t_L g262 ( .A(n_130), .Y(n_262) );
AND2x2_ASAP7_75t_L g387 ( .A(n_130), .B(n_329), .Y(n_387) );
OR2x2_ASAP7_75t_L g389 ( .A(n_130), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .Y(n_130) );
INVx1_ASAP7_75t_L g256 ( .A(n_131), .Y(n_256) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx1_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_133), .B(n_134), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
NAND3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_151), .C(n_153), .Y(n_137) );
AO21x1_ASAP7_75t_L g255 ( .A1(n_138), .A2(n_151), .B(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_141), .B1(n_145), .B2(n_148), .Y(n_138) );
INVx2_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g206 ( .A1(n_139), .A2(n_147), .B1(n_207), .B2(n_209), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_139), .A2(n_145), .B1(n_214), .B2(n_215), .Y(n_213) );
INVx4_ASAP7_75t_L g468 ( .A(n_139), .Y(n_468) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
INVx1_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
AND2x2_ASAP7_75t_L g446 ( .A(n_140), .B(n_168), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_140), .Y(n_449) );
INVx2_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx1_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_145), .A2(n_165), .B(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_145), .A2(n_182), .B(n_183), .C(n_184), .Y(n_181) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_146), .A2(n_162), .B(n_163), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_SL g221 ( .A1(n_146), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_146), .A2(n_244), .B(n_245), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_146), .B(n_496), .Y(n_495) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_149), .Y(n_544) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g201 ( .A(n_150), .Y(n_201) );
BUFx3_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
AND2x6_ASAP7_75t_L g448 ( .A(n_150), .B(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g460 ( .A(n_151), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_151), .B(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_151), .A2(n_512), .B(n_519), .Y(n_511) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_151), .A2(n_539), .B(n_546), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_151), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_152), .A2(n_160), .B(n_169), .Y(n_159) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_152), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_152), .A2(n_524), .B(n_525), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_153), .A2(n_243), .B(n_246), .Y(n_242) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_154), .A2(n_161), .B(n_164), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_154), .A2(n_174), .B(n_181), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_154), .A2(n_193), .B(n_198), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_154), .A2(n_221), .B(n_225), .Y(n_220) );
AND2x4_ASAP7_75t_L g445 ( .A(n_154), .B(n_446), .Y(n_445) );
INVx4_ASAP7_75t_SL g470 ( .A(n_154), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_154), .B(n_446), .Y(n_514) );
INVx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g300 ( .A(n_157), .B(n_272), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_157), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g414 ( .A(n_157), .B(n_254), .Y(n_414) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_170), .Y(n_157) );
AND2x2_ASAP7_75t_L g257 ( .A(n_158), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g304 ( .A(n_158), .Y(n_304) );
AND2x2_ASAP7_75t_L g329 ( .A(n_158), .B(n_241), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_158), .B(n_362), .Y(n_399) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g263 ( .A(n_159), .B(n_241), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_159), .B(n_240), .Y(n_277) );
AND2x2_ASAP7_75t_L g294 ( .A(n_159), .B(n_170), .Y(n_294) );
AND2x2_ASAP7_75t_L g351 ( .A(n_159), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_159), .B(n_258), .Y(n_364) );
AND2x2_ASAP7_75t_L g416 ( .A(n_159), .B(n_341), .Y(n_416) );
INVx2_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g239 ( .A(n_170), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g258 ( .A(n_170), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_170), .B(n_241), .Y(n_335) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_185), .Y(n_170) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_171), .A2(n_242), .B(n_249), .Y(n_241) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_172), .B(n_520), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_178), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_176), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_176), .A2(n_527), .B(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_178), .A2(n_542), .B(n_543), .C(n_544), .Y(n_541) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_179), .A2(n_226), .B(n_227), .Y(n_225) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g452 ( .A(n_180), .Y(n_452) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_182), .A2(n_202), .B(n_247), .C(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_182), .A2(n_451), .B(n_453), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_216), .B(n_229), .Y(n_186) );
INVx1_ASAP7_75t_SL g348 ( .A(n_187), .Y(n_348) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_204), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_189), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
INVx1_ASAP7_75t_L g268 ( .A(n_190), .Y(n_268) );
AND2x2_ASAP7_75t_L g289 ( .A(n_190), .B(n_211), .Y(n_289) );
AND2x2_ASAP7_75t_L g323 ( .A(n_190), .B(n_212), .Y(n_323) );
OR2x2_ASAP7_75t_L g342 ( .A(n_190), .B(n_218), .Y(n_342) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_190), .Y(n_356) );
AND2x2_ASAP7_75t_L g369 ( .A(n_190), .B(n_370), .Y(n_369) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_203), .Y(n_190) );
INVx2_ASAP7_75t_L g210 ( .A(n_191), .Y(n_210) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_191), .A2(n_220), .B(n_228), .Y(n_219) );
INVx1_ASAP7_75t_L g458 ( .A(n_191), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_191), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_191), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_202), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_204), .A2(n_291), .B1(n_292), .B2(n_301), .Y(n_290) );
AND2x2_ASAP7_75t_L g374 ( .A(n_204), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_211), .Y(n_204) );
INVx1_ASAP7_75t_L g235 ( .A(n_205), .Y(n_235) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_205), .Y(n_272) );
INVx1_ASAP7_75t_L g283 ( .A(n_205), .Y(n_283) );
AND2x2_ASAP7_75t_L g298 ( .A(n_205), .B(n_212), .Y(n_298) );
INVx2_ASAP7_75t_L g469 ( .A(n_208), .Y(n_469) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_208), .Y(n_484) );
INVx1_ASAP7_75t_L g455 ( .A(n_210), .Y(n_455) );
OR2x2_ASAP7_75t_L g252 ( .A(n_211), .B(n_237), .Y(n_252) );
AND2x2_ASAP7_75t_L g282 ( .A(n_211), .B(n_283), .Y(n_282) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_211), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g230 ( .A(n_212), .B(n_231), .Y(n_230) );
BUFx2_ASAP7_75t_L g339 ( .A(n_212), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_216), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g317 ( .A(n_217), .B(n_283), .Y(n_317) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g229 ( .A(n_218), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g237 ( .A(n_219), .Y(n_237) );
OR2x2_ASAP7_75t_L g267 ( .A(n_219), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_219), .Y(n_322) );
AOI32xp33_ASAP7_75t_L g359 ( .A1(n_229), .A2(n_289), .A3(n_360), .B1(n_361), .B2(n_363), .Y(n_359) );
AND2x2_ASAP7_75t_L g285 ( .A(n_230), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_230), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_230), .B(n_317), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_230), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_238), .B1(n_251), .B2(n_253), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g338 ( .A(n_234), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_235), .B(n_237), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_236), .A2(n_260), .B1(n_264), .B2(n_274), .Y(n_259) );
AND2x2_ASAP7_75t_L g281 ( .A(n_236), .B(n_282), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_236), .A2(n_250), .B(n_298), .C(n_333), .Y(n_332) );
OAI332xp33_ASAP7_75t_L g337 ( .A1(n_236), .A2(n_338), .A3(n_340), .B1(n_342), .B2(n_343), .B3(n_345), .C1(n_346), .C2(n_348), .Y(n_337) );
INVx2_ASAP7_75t_L g378 ( .A(n_236), .Y(n_378) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
INVx1_ASAP7_75t_L g371 ( .A(n_237), .Y(n_371) );
AND2x2_ASAP7_75t_L g425 ( .A(n_237), .B(n_289), .Y(n_425) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_250), .Y(n_238) );
AND2x2_ASAP7_75t_L g305 ( .A(n_240), .B(n_255), .Y(n_305) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g254 ( .A(n_241), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g353 ( .A(n_241), .B(n_255), .Y(n_353) );
INVx1_ASAP7_75t_L g362 ( .A(n_241), .Y(n_362) );
INVx1_ASAP7_75t_L g336 ( .A(n_250), .Y(n_336) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_272), .Y(n_420) );
INVx1_ASAP7_75t_SL g331 ( .A(n_253), .Y(n_331) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
AND2x2_ASAP7_75t_L g358 ( .A(n_254), .B(n_316), .Y(n_358) );
INVx1_ASAP7_75t_L g377 ( .A(n_254), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_254), .B(n_344), .Y(n_379) );
INVx1_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
AND2x2_ASAP7_75t_L g280 ( .A(n_257), .B(n_261), .Y(n_280) );
AND2x2_ASAP7_75t_L g347 ( .A(n_257), .B(n_305), .Y(n_347) );
INVx2_ASAP7_75t_L g390 ( .A(n_257), .Y(n_390) );
INVx2_ASAP7_75t_L g273 ( .A(n_258), .Y(n_273) );
AND2x2_ASAP7_75t_L g275 ( .A(n_258), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_262), .B(n_335), .Y(n_341) );
OR2x2_ASAP7_75t_L g405 ( .A(n_262), .B(n_364), .Y(n_405) );
INVx1_ASAP7_75t_L g429 ( .A(n_262), .Y(n_429) );
INVx1_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
AND2x2_ASAP7_75t_L g430 ( .A(n_263), .B(n_273), .Y(n_430) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_267), .A2(n_293), .B1(n_295), .B2(n_299), .Y(n_292) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI322xp33_ASAP7_75t_SL g376 ( .A1(n_270), .A2(n_377), .A3(n_378), .B1(n_379), .B2(n_380), .C1(n_383), .C2(n_385), .Y(n_376) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
AND2x2_ASAP7_75t_L g373 ( .A(n_271), .B(n_289), .Y(n_373) );
OR2x2_ASAP7_75t_L g407 ( .A(n_271), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g410 ( .A(n_271), .B(n_342), .Y(n_410) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g355 ( .A(n_272), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g411 ( .A(n_272), .B(n_342), .Y(n_411) );
INVx3_ASAP7_75t_L g344 ( .A(n_273), .Y(n_344) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g400 ( .A(n_275), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g279 ( .A1(n_277), .A2(n_280), .B1(n_281), .B2(n_284), .C1(n_285), .C2(n_287), .Y(n_279) );
INVx1_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_279), .B(n_290), .C(n_307), .Y(n_278) );
AND2x2_ASAP7_75t_L g395 ( .A(n_282), .B(n_296), .Y(n_395) );
BUFx2_ASAP7_75t_L g286 ( .A(n_283), .Y(n_286) );
INVx1_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_284), .A2(n_320), .B1(n_373), .B2(n_374), .C(n_376), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_286), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
AND2x2_ASAP7_75t_L g326 ( .A(n_289), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_294), .B(n_305), .Y(n_306) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OAI21xp33_ASAP7_75t_L g301 ( .A1(n_296), .A2(n_302), .B(n_306), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_296), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g393 ( .A(n_298), .B(n_375), .Y(n_393) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g316 ( .A(n_304), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_305), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g422 ( .A(n_305), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_313), .B1(n_314), .B2(n_317), .C(n_318), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_309), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g418 ( .A(n_317), .B(n_323), .Y(n_418) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OAI31xp33_ASAP7_75t_SL g386 ( .A1(n_321), .A2(n_360), .A3(n_387), .B(n_388), .Y(n_386) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g375 ( .A(n_322), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_323), .B(n_327), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_328), .B1(n_330), .B2(n_331), .C(n_332), .Y(n_324) );
INVx1_ASAP7_75t_L g330 ( .A(n_326), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_329), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g345 ( .A(n_338), .Y(n_345) );
INVx2_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g367 ( .A(n_344), .B(n_353), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_344), .A2(n_361), .B(n_418), .C(n_419), .Y(n_417) );
OAI221xp5_ASAP7_75t_SL g349 ( .A1(n_345), .A2(n_350), .B1(n_354), .B2(n_357), .C(n_359), .Y(n_349) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g412 ( .A1(n_348), .A2(n_413), .B(n_415), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_351), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_391), .C(n_412), .D(n_423), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B(n_372), .C(n_386), .Y(n_366) );
INVx1_ASAP7_75t_SL g421 ( .A(n_373), .Y(n_421) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_SL g384 ( .A(n_382), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_389), .A2(n_398), .B1(n_410), .B2(n_411), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_396), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI31xp33_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_424), .A3(n_426), .B(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_434), .A2(n_436), .B1(n_719), .B2(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_437), .B(n_653), .Y(n_436) );
NOR5xp2_ASAP7_75t_L g437 ( .A(n_438), .B(n_584), .C(n_613), .D(n_633), .E(n_640), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_472), .B(n_529), .C(n_571), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_440), .A2(n_656), .B1(n_658), .B2(n_659), .Y(n_655) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_459), .Y(n_440) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_441), .Y(n_532) );
AND2x4_ASAP7_75t_L g564 ( .A(n_441), .B(n_565), .Y(n_564) );
INVx5_ASAP7_75t_L g582 ( .A(n_441), .Y(n_582) );
AND2x2_ASAP7_75t_L g591 ( .A(n_441), .B(n_583), .Y(n_591) );
AND2x2_ASAP7_75t_L g603 ( .A(n_441), .B(n_476), .Y(n_603) );
AND2x2_ASAP7_75t_L g699 ( .A(n_441), .B(n_567), .Y(n_699) );
OR2x6_ASAP7_75t_L g441 ( .A(n_442), .B(n_456), .Y(n_441) );
AOI21xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_447), .B(n_455), .Y(n_442) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx5_ASAP7_75t_L g464 ( .A(n_448), .Y(n_464) );
INVx2_ASAP7_75t_L g454 ( .A(n_452), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_454), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_454), .A2(n_484), .B(n_506), .C(n_507), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx2_ASAP7_75t_L g565 ( .A(n_459), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_459), .B(n_538), .Y(n_583) );
AND2x2_ASAP7_75t_L g602 ( .A(n_459), .B(n_537), .Y(n_602) );
AND2x2_ASAP7_75t_L g642 ( .A(n_459), .B(n_582), .Y(n_642) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_471), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_464), .B(n_465), .C(n_470), .Y(n_462) );
INVx2_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_464), .A2(n_470), .B(n_493), .C(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g485 ( .A(n_470), .Y(n_485) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_498), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI322xp5_ASAP7_75t_L g701 ( .A1(n_475), .A2(n_509), .A3(n_556), .B1(n_564), .B2(n_618), .C1(n_702), .C2(n_705), .Y(n_701) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_488), .Y(n_475) );
INVx5_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
AND2x2_ASAP7_75t_L g550 ( .A(n_476), .B(n_536), .Y(n_550) );
BUFx2_ASAP7_75t_L g628 ( .A(n_476), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_476), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g705 ( .A(n_476), .B(n_612), .Y(n_705) );
OR2x6_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_488), .B(n_500), .Y(n_559) );
INVx1_ASAP7_75t_L g586 ( .A(n_488), .Y(n_586) );
AND2x2_ASAP7_75t_L g599 ( .A(n_488), .B(n_521), .Y(n_599) );
AND2x2_ASAP7_75t_L g700 ( .A(n_488), .B(n_618), .Y(n_700) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g554 ( .A(n_489), .B(n_500), .Y(n_554) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
OR2x2_ASAP7_75t_L g569 ( .A(n_489), .B(n_521), .Y(n_569) );
AND2x2_ASAP7_75t_L g579 ( .A(n_489), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_489), .B(n_511), .Y(n_608) );
INVxp67_ASAP7_75t_L g632 ( .A(n_489), .Y(n_632) );
AND2x2_ASAP7_75t_L g639 ( .A(n_489), .B(n_509), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_489), .B(n_521), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_489), .B(n_510), .Y(n_665) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_497), .Y(n_489) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_500), .B(n_522), .Y(n_609) );
OR2x2_ASAP7_75t_L g631 ( .A(n_500), .B(n_510), .Y(n_631) );
AND2x2_ASAP7_75t_L g644 ( .A(n_500), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_500), .B(n_599), .Y(n_650) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_500), .A2(n_655), .B(n_660), .C(n_669), .Y(n_654) );
AND2x2_ASAP7_75t_L g715 ( .A(n_500), .B(n_521), .Y(n_715) );
INVx5_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_501), .B(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_501), .B(n_563), .Y(n_575) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_501), .Y(n_577) );
OR2x2_ASAP7_75t_L g588 ( .A(n_501), .B(n_510), .Y(n_588) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_501), .B(n_579), .Y(n_593) );
AND2x2_ASAP7_75t_L g618 ( .A(n_501), .B(n_510), .Y(n_618) );
AND2x2_ASAP7_75t_L g638 ( .A(n_501), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g676 ( .A(n_501), .B(n_509), .Y(n_676) );
OR2x2_ASAP7_75t_L g679 ( .A(n_501), .B(n_665), .Y(n_679) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_510), .A2(n_623), .B(n_626), .C(n_632), .Y(n_622) );
INVx5_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_511), .B(n_521), .Y(n_553) );
AND2x2_ASAP7_75t_L g557 ( .A(n_511), .B(n_522), .Y(n_557) );
OR2x2_ASAP7_75t_L g563 ( .A(n_511), .B(n_521), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_SL g580 ( .A(n_521), .Y(n_580) );
OR2x2_ASAP7_75t_L g708 ( .A(n_521), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_548), .B(n_551), .C(n_560), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI31xp33_ASAP7_75t_L g633 ( .A1(n_531), .A2(n_634), .A3(n_636), .B(n_637), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_532), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_533), .B(n_564), .Y(n_570) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_534), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g590 ( .A(n_534), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g595 ( .A(n_534), .B(n_565), .Y(n_595) );
AND2x2_ASAP7_75t_L g605 ( .A(n_534), .B(n_564), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_534), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g625 ( .A(n_534), .B(n_582), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_534), .B(n_602), .Y(n_630) );
OR2x2_ASAP7_75t_L g649 ( .A(n_534), .B(n_536), .Y(n_649) );
OR2x2_ASAP7_75t_L g651 ( .A(n_534), .B(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_534), .Y(n_698) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g598 ( .A(n_536), .B(n_565), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_536), .B(n_582), .Y(n_621) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g567 ( .A(n_538), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_545), .Y(n_539) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g658 ( .A(n_550), .B(n_582), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g660 ( .A1(n_550), .A2(n_564), .A3(n_602), .B1(n_661), .B2(n_662), .C1(n_663), .C2(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g668 ( .A(n_550), .Y(n_668) );
NAND2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_SL g662 ( .A(n_552), .Y(n_662) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OR2x2_ASAP7_75t_L g614 ( .A(n_553), .B(n_559), .Y(n_614) );
INVx1_ASAP7_75t_L g645 ( .A(n_553), .Y(n_645) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI32xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .A3(n_566), .B1(n_568), .B2(n_570), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AOI21xp33_ASAP7_75t_SL g600 ( .A1(n_563), .A2(n_578), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_SL g615 ( .A(n_564), .Y(n_615) );
AND2x4_ASAP7_75t_L g612 ( .A(n_565), .B(n_582), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_565), .B(n_648), .Y(n_647) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_566), .A2(n_593), .A3(n_612), .B1(n_645), .B2(n_678), .C1(n_680), .C2(n_681), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_566), .A2(n_643), .B1(n_707), .B2(n_708), .C(n_710), .Y(n_706) );
AND2x2_ASAP7_75t_L g594 ( .A(n_567), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g574 ( .A(n_569), .Y(n_574) );
OR2x2_ASAP7_75t_L g646 ( .A(n_569), .B(n_631), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .A3(n_576), .B(n_581), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_572), .A2(n_605), .B1(n_606), .B2(n_610), .Y(n_604) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g617 ( .A(n_574), .B(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_576), .A2(n_617), .B1(n_670), .B2(n_673), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g659 ( .A(n_579), .B(n_628), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_579), .B(n_618), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_580), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g693 ( .A(n_580), .B(n_631), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_581), .A2(n_676), .B1(n_689), .B2(n_692), .Y(n_688) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g597 ( .A(n_582), .Y(n_597) );
AND2x2_ASAP7_75t_L g680 ( .A(n_582), .B(n_602), .Y(n_680) );
OR2x2_ASAP7_75t_L g682 ( .A(n_582), .B(n_649), .Y(n_682) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_582), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_583), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_583), .B(n_628), .Y(n_636) );
OAI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B(n_592), .C(n_604), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_596), .B2(n_599), .C(n_600), .Y(n_592) );
INVxp67_ASAP7_75t_L g704 ( .A(n_595), .Y(n_704) );
INVx1_ASAP7_75t_L g671 ( .A(n_596), .Y(n_671) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g635 ( .A(n_597), .B(n_602), .Y(n_635) );
INVx1_ASAP7_75t_L g652 ( .A(n_598), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_598), .B(n_625), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g667 ( .A(n_602), .Y(n_667) );
AND2x2_ASAP7_75t_L g673 ( .A(n_602), .B(n_628), .Y(n_673) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_SL g661 ( .A(n_609), .Y(n_661) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_612), .B(n_648), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_616), .B2(n_619), .C(n_622), .Y(n_613) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g709 ( .A(n_618), .Y(n_709) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g627 ( .A(n_621), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_625), .B(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_631), .Y(n_626) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_629), .A2(n_675), .B(n_677), .C(n_683), .Y(n_674) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g686 ( .A(n_631), .Y(n_686) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI222xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_646), .B2(n_647), .C1(n_650), .C2(n_651), .Y(n_640) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g716 ( .A(n_647), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_648), .B(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_648), .A2(n_695), .B1(n_697), .B2(n_700), .Y(n_694) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
NOR4xp25_ASAP7_75t_L g653 ( .A(n_654), .B(n_674), .C(n_687), .D(n_706), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_656), .B(n_686), .Y(n_696) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g663 ( .A(n_661), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_664), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_694), .C(n_701), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_L g703 ( .A(n_699), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_713), .B(n_716), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g739 ( .A(n_727), .Y(n_739) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g743 ( .A(n_731), .Y(n_743) );
INVx1_ASAP7_75t_L g736 ( .A(n_733), .Y(n_736) );
BUFx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
endmodule