module fake_jpeg_5542_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_53),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_21),
.B1(n_27),
.B2(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_1),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_65),
.Y(n_104)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_76),
.B1(n_8),
.B2(n_9),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_1),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_17),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_73),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_32),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_9),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_39),
.A2(n_28),
.B1(n_23),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_26),
.B1(n_24),
.B2(n_15),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_15),
.B1(n_27),
.B2(n_25),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_21),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_12),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_80),
.B1(n_57),
.B2(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_95),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_111),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_8),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_104),
.B(n_89),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_86),
.B1(n_59),
.B2(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_64),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_13),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_110),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_68),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_110),
.C(n_111),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_122),
.C(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_123),
.B1(n_109),
.B2(n_81),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_107),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_77),
.C(n_75),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_71),
.B1(n_67),
.B2(n_65),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_106),
.B(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_58),
.C(n_83),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_72),
.B(n_64),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_109),
.Y(n_144)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_91),
.CON(n_132),
.SN(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NOR4xp25_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_142),
.C(n_100),
.D(n_96),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_105),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_139),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_124),
.B(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_93),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_103),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_143),
.C(n_130),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_90),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_147),
.B(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_118),
.B1(n_125),
.B2(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_146),
.B1(n_149),
.B2(n_148),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_117),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_155),
.C(n_140),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_160),
.B(n_162),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_96),
.C(n_100),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_141),
.C(n_145),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_120),
.B1(n_96),
.B2(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_145),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_100),
.B(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_170),
.C(n_171),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_135),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_166),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_146),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_139),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_135),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_150),
.B1(n_153),
.B2(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_168),
.B1(n_165),
.B2(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_178),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_158),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_134),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_173),
.C(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_176),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_182),
.B(n_179),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_178),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_187),
.Y(n_188)
);


endmodule