module fake_jpeg_15990_n_223 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_223);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_36),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_0),
.CON(n_29),
.SN(n_29)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_16),
.CON(n_39),
.SN(n_39)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_6),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_27),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_44),
.B1(n_54),
.B2(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_20),
.B1(n_18),
.B2(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_25),
.B1(n_13),
.B2(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_31),
.A2(n_25),
.B1(n_26),
.B2(n_15),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_42),
.C(n_43),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_66),
.C(n_38),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_65),
.B1(n_73),
.B2(n_41),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_30),
.B1(n_42),
.B2(n_39),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_37),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_37),
.C(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_51),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_40),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_97),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_70),
.B1(n_68),
.B2(n_72),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_80),
.B1(n_51),
.B2(n_52),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_92),
.B(n_66),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_51),
.C(n_45),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_45),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_72),
.B(n_68),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_33),
.B(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_15),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_26),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_40),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_103),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_37),
.B(n_17),
.C(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_66),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_40),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_113),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_102),
.B(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_109),
.B(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_122),
.B(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_63),
.B1(n_73),
.B2(n_52),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_119),
.B1(n_80),
.B2(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_77),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_124),
.B1(n_89),
.B2(n_91),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_88),
.C(n_97),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_88),
.C(n_82),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_63),
.B(n_76),
.C(n_52),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_60),
.B1(n_66),
.B2(n_51),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_83),
.B(n_74),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_132),
.C(n_136),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_133),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_89),
.C(n_84),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_138),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_87),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_91),
.B1(n_85),
.B2(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_149),
.B1(n_111),
.B2(n_110),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_145),
.B1(n_134),
.B2(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_102),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_93),
.C(n_85),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_53),
.B1(n_51),
.B2(n_86),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_112),
.B1(n_118),
.B2(n_111),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_165),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_107),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_136),
.C(n_147),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_122),
.B1(n_124),
.B2(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_122),
.B1(n_109),
.B2(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_115),
.B1(n_119),
.B2(n_98),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_98),
.B(n_86),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_146),
.B(n_133),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_175),
.C(n_177),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_155),
.B(n_131),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_178),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_140),
.Y(n_173)
);

AOI321xp33_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_171),
.A3(n_172),
.B1(n_185),
.B2(n_157),
.C(n_184),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_129),
.B(n_143),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_128),
.C(n_149),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_129),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_139),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_98),
.B(n_1),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_79),
.C(n_34),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_183),
.C(n_150),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_79),
.C(n_34),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_53),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_183),
.CI(n_169),
.CON(n_200),
.SN(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_195),
.C(n_35),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_153),
.C(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_35),
.C(n_34),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_197),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_177),
.B(n_69),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_180),
.B(n_185),
.C(n_173),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_190),
.B(n_193),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_206),
.C(n_35),
.Y(n_211)
);

OAI31xp33_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_178),
.A3(n_181),
.B(n_2),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_203),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

OAI221xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_194),
.B1(n_192),
.B2(n_195),
.C(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_210),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_212),
.B(n_204),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_5),
.B(n_10),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_206),
.C(n_200),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_202),
.C(n_199),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_12),
.C(n_22),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

AOI21x1_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_216),
.B(n_3),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_220),
.B(n_12),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_22),
.Y(n_223)
);


endmodule