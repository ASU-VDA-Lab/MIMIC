module fake_jpeg_9969_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_21),
.B1(n_30),
.B2(n_20),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_58),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_50),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_74),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_78),
.B1(n_80),
.B2(n_85),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_44),
.B1(n_39),
.B2(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_75),
.B1(n_56),
.B2(n_63),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_41),
.C(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_62),
.B1(n_56),
.B2(n_46),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_27),
.B1(n_33),
.B2(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_34),
.B1(n_33),
.B2(n_25),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_19),
.B1(n_27),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_59),
.B1(n_64),
.B2(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_94),
.Y(n_116)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_46),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_109),
.B(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_77),
.B(n_81),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_115),
.B1(n_102),
.B2(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_103),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_76),
.C(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.C(n_31),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_83),
.C(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_58),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_53),
.B1(n_64),
.B2(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_129),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_92),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_32),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_100),
.B1(n_110),
.B2(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_125),
.B1(n_131),
.B2(n_109),
.Y(n_144)
);

BUFx16f_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_107),
.B1(n_101),
.B2(n_95),
.Y(n_125)
);

NOR2x1_ASAP7_75t_R g164 ( 
.A(n_128),
.B(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_79),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_82),
.B1(n_53),
.B2(n_81),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_137),
.C(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_2),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_69),
.C(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_99),
.B(n_112),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_32),
.B(n_24),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_113),
.B1(n_108),
.B2(n_92),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_148),
.B(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_115),
.B1(n_104),
.B2(n_92),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_29),
.B(n_28),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_119),
.C(n_132),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_60),
.C(n_32),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_133),
.C(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_125),
.B1(n_136),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_24),
.B1(n_60),
.B2(n_16),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_2),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_3),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_118),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_185),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_186),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_126),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_126),
.C(n_120),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_192),
.B1(n_148),
.B2(n_121),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_138),
.B1(n_131),
.B2(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NOR4xp25_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_160),
.C(n_164),
.D(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_201),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_149),
.B(n_157),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_207),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_149),
.B(n_150),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_161),
.B(n_155),
.C(n_139),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_206),
.B1(n_211),
.B2(n_212),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_147),
.B(n_155),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_210),
.B1(n_213),
.B2(n_179),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_153),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_185),
.C(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_220),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_176),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_222),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_180),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_206),
.C(n_196),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_225),
.B(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_175),
.C(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_175),
.C(n_173),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_228),
.B(n_213),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_183),
.B1(n_172),
.B2(n_182),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_4),
.B(n_7),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_200),
.C(n_202),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_209),
.B1(n_210),
.B2(n_156),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_142),
.B1(n_141),
.B2(n_6),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_223),
.B(n_216),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_241),
.B(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_217),
.C(n_225),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_9),
.B(n_10),
.Y(n_241)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_248),
.Y(n_255)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_251),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_252),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_232),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_238),
.B(n_218),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.C(n_233),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_261),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_239),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_254),
.B(n_12),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_11),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_244),
.A3(n_250),
.B1(n_236),
.B2(n_13),
.C1(n_10),
.C2(n_15),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_267),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_11),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_270),
.A2(n_271),
.B(n_264),
.Y(n_272)
);

OAI311xp33_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_262),
.A3(n_268),
.B1(n_15),
.C1(n_13),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_273),
.B(n_14),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_275),
.A2(n_15),
.B(n_13),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_14),
.Y(n_277)
);


endmodule