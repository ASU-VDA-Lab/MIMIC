module fake_netlist_1_2385_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_8), .B(n_1), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
OAI22xp5_ASAP7_75t_SL g19 ( .A1(n_11), .A2(n_0), .B1(n_3), .B2(n_5), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_14), .B(n_3), .C(n_5), .Y(n_20) );
OAI22xp33_ASAP7_75t_L g21 ( .A1(n_10), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_13), .Y(n_22) );
AND2x4_ASAP7_75t_SL g23 ( .A(n_20), .B(n_16), .Y(n_23) );
CKINVDCx16_ASAP7_75t_R g24 ( .A(n_19), .Y(n_24) );
AND2x2_ASAP7_75t_SL g25 ( .A(n_18), .B(n_16), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_18), .B(n_10), .Y(n_26) );
INVx3_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_23), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_25), .B1(n_23), .B2(n_17), .Y(n_30) );
AO22x1_ASAP7_75t_L g31 ( .A1(n_27), .A2(n_16), .B1(n_15), .B2(n_12), .Y(n_31) );
AOI221x1_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_22), .B1(n_12), .B2(n_29), .C(n_13), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_27), .B1(n_21), .B2(n_22), .C1(n_28), .C2(n_7), .Y(n_33) );
BUFx2_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
XNOR2xp5_ASAP7_75t_L g36 ( .A(n_34), .B(n_28), .Y(n_36) );
OAI22x1_ASAP7_75t_SL g37 ( .A1(n_35), .A2(n_27), .B1(n_33), .B2(n_34), .Y(n_37) );
AOI22xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_27), .B1(n_36), .B2(n_33), .Y(n_38) );
endmodule