module fake_jpeg_808_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_36),
.B(n_57),
.Y(n_73)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_1),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_44),
.B(n_23),
.C(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_2),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_16),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_65),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_83),
.B1(n_87),
.B2(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_30),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_15),
.B1(n_27),
.B2(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_90),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_40),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_34),
.B1(n_15),
.B2(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_97),
.B1(n_74),
.B2(n_85),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_46),
.B1(n_41),
.B2(n_37),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_78),
.B1(n_48),
.B2(n_85),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_49),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_21),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_109),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_77),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_63),
.B(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_51),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_3),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_78),
.B1(n_61),
.B2(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_119),
.B1(n_131),
.B2(n_97),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_135),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_3),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_133),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_3),
.B1(n_5),
.B2(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_5),
.B1(n_104),
.B2(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_94),
.B1(n_89),
.B2(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_103),
.B(n_109),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_145),
.B(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_89),
.B(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_114),
.B1(n_113),
.B2(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_153),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_115),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_121),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_120),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_144),
.C(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_163),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_127),
.B(n_120),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_145),
.B(n_143),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_117),
.B(n_119),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_165),
.B(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_144),
.B1(n_154),
.B2(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_177),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.C(n_164),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_134),
.C(n_111),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_157),
.B(n_155),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_160),
.B1(n_158),
.B2(n_166),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_169),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_185),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_166),
.B(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_167),
.B1(n_162),
.B2(n_129),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_187),
.B1(n_182),
.B2(n_186),
.Y(n_196)
);

AOI31xp67_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_175),
.A3(n_176),
.B(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_173),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_185),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_187),
.C(n_192),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_181),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_189),
.B(n_162),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_197),
.B(n_194),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_203),
.B(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_195),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_123),
.B(n_129),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_123),
.Y(n_206)
);


endmodule