module fake_netlist_6_4249_n_1063 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1063);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1063;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_875;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_427;
wire n_288;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_230),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_27),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_24),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_54),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_40),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_171),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_175),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_21),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_82),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_20),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_46),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_137),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_83),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_53),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_60),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_18),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_108),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_9),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_75),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_190),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_189),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_121),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_195),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_49),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_133),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_64),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_88),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_106),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_25),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_101),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_18),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_30),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_134),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_161),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_78),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_90),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_70),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_8),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_191),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_87),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_47),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_32),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_213),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_103),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_156),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_209),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_99),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_143),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_84),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_34),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_194),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_146),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_132),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_14),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_34),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_211),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_218),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_145),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_2),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_110),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_212),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_57),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_73),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_127),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_196),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_27),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_68),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_112),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_17),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_207),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_58),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_236),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_0),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_246),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_251),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_239),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_234),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_244),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_258),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_267),
.B(n_1),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_251),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_233),
.B(n_2),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_3),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_263),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_235),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_238),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_240),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_247),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_263),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_237),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_274),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_289),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_289),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_271),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_241),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_308),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_308),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_245),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_282),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_324),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_277),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_284),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_255),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_232),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_285),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_291),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_259),
.B(n_4),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_256),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_324),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_259),
.B(n_4),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_261),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_232),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_264),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_262),
.B(n_5),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_297),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_242),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_283),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_311),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_R g386 ( 
.A(n_243),
.B(n_41),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_315),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_262),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_349),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_312),
.B(n_281),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_383),
.B(n_340),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_333),
.B(n_281),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_382),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_312),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_276),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_279),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_354),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_334),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_370),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_346),
.B(n_290),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

NAND2x1p5_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_265),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_355),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_294),
.Y(n_415)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_298),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_378),
.B(n_257),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_339),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_358),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_301),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_350),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_367),
.B(n_303),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_356),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_387),
.B(n_367),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_386),
.A2(n_320),
.B(n_318),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_426),
.B(n_352),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_R g449 ( 
.A(n_404),
.B(n_385),
.Y(n_449)
);

AND2x4_ASAP7_75t_SL g450 ( 
.A(n_430),
.B(n_357),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_416),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_415),
.A2(n_327),
.B1(n_322),
.B2(n_385),
.Y(n_453)
);

BUFx8_ASAP7_75t_SL g454 ( 
.A(n_439),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_L g455 ( 
.A(n_415),
.B(n_248),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_416),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_249),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_415),
.A2(n_421),
.B1(n_422),
.B2(n_401),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_419),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_422),
.B(n_250),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_398),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_252),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_253),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_415),
.A2(n_257),
.B1(n_309),
.B2(n_283),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_257),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_413),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_361),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_425),
.B(n_362),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g475 ( 
.A1(n_424),
.A2(n_292),
.B1(n_304),
.B2(n_310),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_415),
.B(n_254),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_415),
.B(n_266),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_403),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_401),
.A2(n_309),
.B1(n_283),
.B2(n_326),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_309),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_403),
.B(n_42),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_442),
.B(n_268),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_292),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_443),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_404),
.B(n_365),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_412),
.B(n_375),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_439),
.A2(n_304),
.B1(n_310),
.B2(n_270),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_402),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_401),
.A2(n_328),
.B1(n_325),
.B2(n_321),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_403),
.A2(n_319),
.B1(n_317),
.B2(n_316),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_388),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_313),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_393),
.Y(n_507)
);

NOR2x1p5_ASAP7_75t_L g508 ( 
.A(n_408),
.B(n_269),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_388),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_272),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_443),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_395),
.A2(n_307),
.B1(n_305),
.B2(n_302),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_390),
.Y(n_514)
);

INVxp33_ASAP7_75t_SL g515 ( 
.A(n_433),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_396),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_428),
.A2(n_299),
.B1(n_296),
.B2(n_293),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_412),
.A2(n_288),
.B1(n_287),
.B2(n_278),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_438),
.B(n_275),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_397),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_409),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_483),
.B(n_392),
.Y(n_526)
);

INVx8_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_483),
.B(n_399),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_458),
.B(n_430),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_429),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_512),
.B(n_430),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_525),
.B(n_431),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_447),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_453),
.A2(n_436),
.B1(n_444),
.B2(n_445),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_525),
.B(n_430),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_459),
.B(n_434),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_514),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_500),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_457),
.B(n_432),
.Y(n_543)
);

BUFx5_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_458),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_454),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_497),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_463),
.B(n_441),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_488),
.A2(n_436),
.B1(n_444),
.B2(n_446),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_463),
.B(n_432),
.Y(n_550)
);

AOI221xp5_ASAP7_75t_L g551 ( 
.A1(n_475),
.A2(n_484),
.B1(n_496),
.B2(n_470),
.C(n_494),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_R g552 ( 
.A(n_524),
.B(n_405),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_458),
.B(n_432),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_488),
.B(n_432),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_436),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_497),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_465),
.B(n_388),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_469),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_457),
.B(n_397),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_499),
.A2(n_437),
.B1(n_117),
.B2(n_118),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_516),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_457),
.B(n_437),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_457),
.B(n_43),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_520),
.B(n_5),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_511),
.B(n_6),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_505),
.B(n_507),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_516),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_467),
.B(n_6),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_518),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_451),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_518),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_454),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_522),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_519),
.B(n_231),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_477),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_477),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_505),
.B(n_44),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_480),
.B(n_45),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_507),
.B(n_48),
.Y(n_583)
);

A2O1A1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_482),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_478),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_452),
.B(n_50),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_489),
.B(n_7),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_510),
.B(n_51),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_510),
.B(n_52),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_488),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_472),
.B(n_55),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_481),
.B(n_56),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_476),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_490),
.B(n_59),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_491),
.B(n_61),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_478),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_501),
.B(n_62),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_489),
.B(n_10),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_479),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_449),
.Y(n_602)
);

AO22x1_ASAP7_75t_L g603 ( 
.A1(n_488),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_462),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_460),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_524),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_449),
.A2(n_128),
.B1(n_228),
.B2(n_225),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_506),
.B(n_63),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_488),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_569),
.A2(n_455),
.B(n_456),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_515),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_580),
.A2(n_455),
.B(n_456),
.Y(n_613)
);

AOI21x1_ASAP7_75t_L g614 ( 
.A1(n_583),
.A2(n_464),
.B(n_460),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_528),
.B(n_456),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_587),
.A2(n_473),
.B(n_502),
.C(n_474),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_526),
.B(n_515),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_539),
.B(n_521),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_587),
.A2(n_466),
.B(n_508),
.C(n_452),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_566),
.Y(n_621)
);

AO21x1_ASAP7_75t_L g622 ( 
.A1(n_565),
.A2(n_448),
.B(n_450),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_599),
.A2(n_495),
.B(n_513),
.C(n_450),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_610),
.A2(n_492),
.B1(n_475),
.B2(n_471),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_585),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_590),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_533),
.B(n_488),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_585),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_533),
.B(n_471),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_531),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_542),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_529),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_547),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_555),
.B(n_492),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_605),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_471),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_550),
.B(n_487),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_588),
.A2(n_503),
.B(n_485),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_552),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_590),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_589),
.A2(n_503),
.B(n_485),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_531),
.B(n_492),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_558),
.A2(n_503),
.B(n_485),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_550),
.B(n_464),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_548),
.B(n_492),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_548),
.B(n_487),
.Y(n_648)
);

AO21x1_ASAP7_75t_L g649 ( 
.A1(n_565),
.A2(n_509),
.B(n_504),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_568),
.B(n_487),
.C(n_504),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_560),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_544),
.B(n_487),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_573),
.B(n_504),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_610),
.B(n_509),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_561),
.B(n_509),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_554),
.A2(n_475),
.B1(n_486),
.B2(n_131),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_599),
.A2(n_568),
.B(n_571),
.C(n_534),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_545),
.B(n_14),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_607),
.B(n_553),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_543),
.A2(n_486),
.B(n_130),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_591),
.B(n_65),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_486),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_543),
.A2(n_486),
.B(n_135),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_537),
.B(n_486),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_581),
.A2(n_129),
.B(n_224),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_581),
.A2(n_126),
.B(n_223),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_549),
.A2(n_535),
.B(n_593),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_593),
.A2(n_125),
.B(n_221),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_586),
.Y(n_672)
);

OAI321xp33_ASAP7_75t_L g673 ( 
.A1(n_551),
.A2(n_15),
.A3(n_16),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_544),
.B(n_66),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_654),
.A2(n_549),
.B(n_537),
.Y(n_675)
);

CKINVDCx14_ASAP7_75t_R g676 ( 
.A(n_624),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_616),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_618),
.B(n_561),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_630),
.B(n_571),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_611),
.A2(n_609),
.B(n_532),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_629),
.B(n_648),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_619),
.B(n_544),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_613),
.A2(n_627),
.B(n_639),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_642),
.A2(n_544),
.B(n_564),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_617),
.A2(n_567),
.B(n_564),
.C(n_562),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_612),
.B(n_594),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_624),
.A2(n_577),
.B1(n_604),
.B2(n_535),
.Y(n_687)
);

AOI22x1_ASAP7_75t_L g688 ( 
.A1(n_670),
.A2(n_582),
.B1(n_574),
.B2(n_572),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_621),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_659),
.A2(n_584),
.B(n_570),
.C(n_576),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_L g691 ( 
.A1(n_623),
.A2(n_643),
.B1(n_647),
.B2(n_658),
.C(n_637),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_625),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_626),
.B(n_586),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_646),
.A2(n_544),
.B(n_598),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_635),
.B(n_527),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_631),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_672),
.B(n_544),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_640),
.B(n_552),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_632),
.B(n_527),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_660),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_672),
.B(n_597),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_646),
.A2(n_674),
.B(n_615),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_672),
.B(n_600),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_674),
.A2(n_596),
.B(n_592),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_632),
.B(n_527),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_626),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_645),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_644),
.A2(n_595),
.B(n_557),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_638),
.B(n_636),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_633),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_664),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_651),
.Y(n_713)
);

O2A1O1Ixp5_ASAP7_75t_SL g714 ( 
.A1(n_670),
.A2(n_634),
.B(n_673),
.C(n_652),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_657),
.A2(n_556),
.B(n_530),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_652),
.A2(n_541),
.B(n_538),
.Y(n_716)
);

AND3x1_ASAP7_75t_SL g717 ( 
.A(n_673),
.B(n_603),
.C(n_546),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_SL g718 ( 
.A1(n_640),
.A2(n_575),
.B1(n_608),
.B2(n_601),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_641),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_650),
.A2(n_606),
.B1(n_536),
.B2(n_19),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_664),
.B(n_15),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_650),
.A2(n_16),
.B1(n_22),
.B2(n_23),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_641),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_622),
.B(n_22),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_SL g727 ( 
.A1(n_634),
.A2(n_23),
.B(n_24),
.C(n_26),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_655),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_653),
.B(n_28),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_628),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_662),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_686),
.B(n_679),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_692),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_699),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_683),
.A2(n_614),
.B(n_649),
.Y(n_735)
);

OAI221xp5_ASAP7_75t_L g736 ( 
.A1(n_687),
.A2(n_661),
.B1(n_669),
.B2(n_668),
.C(n_671),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_678),
.A2(n_666),
.B(n_663),
.C(n_667),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_677),
.Y(n_738)
);

CKINVDCx11_ASAP7_75t_R g739 ( 
.A(n_728),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_703),
.A2(n_653),
.B(n_656),
.Y(n_740)
);

BUFx4f_ASAP7_75t_L g741 ( 
.A(n_707),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_716),
.A2(n_665),
.B(n_656),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_685),
.A2(n_656),
.B(n_665),
.C(n_30),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_720),
.A2(n_28),
.A3(n_29),
.B(n_31),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_694),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_712),
.B(n_29),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_689),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_692),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_697),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_720),
.A2(n_31),
.A3(n_32),
.B(n_33),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_691),
.B(n_67),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_722),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_705),
.A2(n_148),
.B(n_220),
.Y(n_753)
);

AO31x2_ASAP7_75t_L g754 ( 
.A1(n_675),
.A2(n_35),
.A3(n_36),
.B(n_37),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_676),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_710),
.B(n_38),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_682),
.A2(n_694),
.B1(n_681),
.B2(n_708),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_709),
.A2(n_69),
.B(n_72),
.Y(n_758)
);

AO31x2_ASAP7_75t_L g759 ( 
.A1(n_726),
.A2(n_74),
.A3(n_76),
.B(n_77),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_701),
.B(n_79),
.Y(n_760)
);

OAI222xp33_ASAP7_75t_L g761 ( 
.A1(n_722),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.C1(n_86),
.C2(n_89),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_684),
.A2(n_91),
.B(n_92),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_714),
.A2(n_93),
.B(n_94),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_711),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_729),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_718),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_724),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_767)
);

AO31x2_ASAP7_75t_L g768 ( 
.A1(n_680),
.A2(n_98),
.A3(n_100),
.B(n_102),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_707),
.Y(n_769)
);

NAND3x1_ASAP7_75t_L g770 ( 
.A(n_721),
.B(n_104),
.C(n_105),
.Y(n_770)
);

AO21x1_ASAP7_75t_L g771 ( 
.A1(n_690),
.A2(n_107),
.B(n_113),
.Y(n_771)
);

AOI221xp5_ASAP7_75t_SL g772 ( 
.A1(n_713),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.C(n_119),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_695),
.A2(n_120),
.B(n_122),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_715),
.A2(n_123),
.B(n_124),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_696),
.B(n_136),
.Y(n_775)
);

AOI221xp5_ASAP7_75t_SL g776 ( 
.A1(n_731),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.C(n_141),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_688),
.A2(n_142),
.B(n_144),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_698),
.A2(n_702),
.B(n_704),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_730),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_693),
.B(n_147),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_700),
.A2(n_706),
.B(n_725),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_725),
.A2(n_149),
.B(n_150),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_749),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_764),
.Y(n_785)
);

INVx6_ASAP7_75t_L g786 ( 
.A(n_769),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_779),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_747),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_766),
.A2(n_717),
.B1(n_723),
.B2(n_719),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_778),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_754),
.Y(n_791)
);

BUFx4f_ASAP7_75t_L g792 ( 
.A(n_733),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_774),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_732),
.A2(n_723),
.B1(n_719),
.B2(n_707),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_751),
.A2(n_756),
.B1(n_765),
.B2(n_771),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_765),
.B(n_723),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_754),
.B(n_727),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_754),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_758),
.Y(n_799)
);

BUFx8_ASAP7_75t_SL g800 ( 
.A(n_734),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_744),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_739),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_751),
.A2(n_719),
.B1(n_152),
.B2(n_153),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_744),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_741),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_746),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_741),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_744),
.B(n_151),
.Y(n_808)
);

INVx6_ASAP7_75t_L g809 ( 
.A(n_760),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_750),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_775),
.B(n_229),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_750),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_733),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_SL g815 ( 
.A1(n_755),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_750),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_SL g817 ( 
.A1(n_736),
.A2(n_763),
.B1(n_757),
.B2(n_761),
.Y(n_817)
);

INVx6_ASAP7_75t_L g818 ( 
.A(n_745),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_777),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_735),
.Y(n_820)
);

INVx6_ASAP7_75t_L g821 ( 
.A(n_748),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_780),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_768),
.Y(n_823)
);

CKINVDCx6p67_ASAP7_75t_R g824 ( 
.A(n_770),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_753),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_759),
.B(n_219),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_768),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_759),
.B(n_167),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_743),
.Y(n_830)
);

INVx6_ASAP7_75t_L g831 ( 
.A(n_781),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_762),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_782),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_773),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_740),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_759),
.Y(n_836)
);

INVx4_ASAP7_75t_SL g837 ( 
.A(n_768),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_752),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_783),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_819),
.A2(n_737),
.B(n_772),
.Y(n_840)
);

AO21x2_ASAP7_75t_L g841 ( 
.A1(n_819),
.A2(n_767),
.B(n_776),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_785),
.B(n_776),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_784),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_787),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_801),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_792),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_791),
.Y(n_847)
);

NOR2x1_ASAP7_75t_R g848 ( 
.A(n_788),
.B(n_772),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_804),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_798),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_810),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_818),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_838),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_789),
.B(n_179),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_812),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_816),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_808),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_788),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_808),
.B(n_180),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_836),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_796),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_817),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_806),
.B(n_186),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_827),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_790),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_790),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_835),
.B(n_187),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_831),
.B(n_188),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_795),
.A2(n_193),
.B(n_197),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_835),
.A2(n_198),
.B(n_199),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_823),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_809),
.B(n_200),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_830),
.B(n_201),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_807),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_809),
.B(n_202),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_786),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_823),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_807),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_831),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_828),
.Y(n_882)
);

AO21x2_ASAP7_75t_L g883 ( 
.A1(n_799),
.A2(n_203),
.B(n_205),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_814),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_786),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_826),
.B(n_214),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_R g888 ( 
.A(n_876),
.B(n_805),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_870),
.A2(n_834),
.B(n_833),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_848),
.B(n_809),
.Y(n_890)
);

AO21x2_ASAP7_75t_L g891 ( 
.A1(n_840),
.A2(n_797),
.B(n_820),
.Y(n_891)
);

AO21x2_ASAP7_75t_L g892 ( 
.A1(n_840),
.A2(n_797),
.B(n_799),
.Y(n_892)
);

OA21x2_ASAP7_75t_L g893 ( 
.A1(n_845),
.A2(n_814),
.B(n_829),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_866),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_857),
.B(n_829),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_862),
.A2(n_826),
.B(n_811),
.C(n_803),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_872),
.A2(n_834),
.B(n_833),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_858),
.B(n_824),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_860),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_839),
.B(n_837),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_847),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_843),
.B(n_837),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_850),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_849),
.B(n_837),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_867),
.B(n_851),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_855),
.B(n_837),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_856),
.B(n_793),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_885),
.B(n_793),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_871),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_885),
.B(n_793),
.Y(n_911)
);

OAI221xp5_ASAP7_75t_L g912 ( 
.A1(n_854),
.A2(n_815),
.B1(n_825),
.B2(n_832),
.C(n_822),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_854),
.A2(n_792),
.B(n_824),
.C(n_794),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_844),
.B(n_831),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_869),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_873),
.B(n_818),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_879),
.B(n_215),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_882),
.B(n_818),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_861),
.B(n_818),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_868),
.A2(n_802),
.B1(n_786),
.B2(n_792),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_900),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_894),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_894),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_894),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_914),
.B(n_863),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_900),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_906),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_911),
.B(n_850),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_911),
.B(n_884),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_893),
.B(n_865),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_898),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_893),
.B(n_852),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_914),
.B(n_881),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_906),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_889),
.A2(n_868),
.B1(n_887),
.B2(n_859),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_898),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_904),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_893),
.B(n_852),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_888),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_910),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_909),
.B(n_881),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_904),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_909),
.B(n_903),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_943),
.B(n_905),
.Y(n_944)
);

OAI221xp5_ASAP7_75t_L g945 ( 
.A1(n_935),
.A2(n_889),
.B1(n_897),
.B2(n_912),
.C(n_896),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_930),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_SL g947 ( 
.A(n_939),
.B(n_915),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_943),
.B(n_905),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_930),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_943),
.B(n_907),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_943),
.B(n_907),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_927),
.B(n_893),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_941),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_932),
.B(n_909),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_922),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_932),
.B(n_909),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_922),
.Y(n_957)
);

NOR3xp33_ASAP7_75t_L g958 ( 
.A(n_935),
.B(n_897),
.C(n_912),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_922),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_925),
.Y(n_960)
);

NAND2x1_ASAP7_75t_L g961 ( 
.A(n_953),
.B(n_938),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_946),
.B(n_921),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_946),
.B(n_926),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_959),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_949),
.B(n_942),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_944),
.B(n_941),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_952),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_947),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_954),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_958),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_966),
.B(n_945),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_962),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_964),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_965),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_960),
.B(n_949),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_963),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_967),
.B(n_949),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_961),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_972),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_970),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_973),
.A2(n_945),
.B(n_958),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_974),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_973),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_984),
.B(n_974),
.Y(n_986)
);

AOI21xp33_ASAP7_75t_SL g987 ( 
.A1(n_983),
.A2(n_985),
.B(n_980),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_983),
.A2(n_978),
.B1(n_976),
.B2(n_971),
.C(n_975),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_982),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_SL g990 ( 
.A1(n_981),
.A2(n_890),
.B(n_896),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_987),
.A2(n_990),
.B(n_988),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_986),
.B(n_947),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_989),
.B(n_979),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_986),
.A2(n_890),
.B1(n_899),
.B2(n_915),
.Y(n_994)
);

AOI31xp33_ASAP7_75t_L g995 ( 
.A1(n_987),
.A2(n_899),
.A3(n_868),
.B(n_920),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_991),
.A2(n_913),
.B(n_979),
.C(n_920),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_993),
.B(n_977),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_992),
.A2(n_915),
.B1(n_953),
.B2(n_887),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_995),
.B(n_956),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_994),
.B(n_953),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_993),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_993),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_991),
.B(n_956),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_992),
.B(n_953),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_1004),
.B(n_880),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_1001),
.B(n_956),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_1002),
.B(n_874),
.C(n_877),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_956),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_996),
.A2(n_998),
.B1(n_999),
.B2(n_1000),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_997),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_1001),
.B(n_800),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_997),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_1005),
.A2(n_853),
.B(n_869),
.C(n_859),
.Y(n_1013)
);

OAI222xp33_ASAP7_75t_L g1014 ( 
.A1(n_1009),
.A2(n_915),
.B1(n_869),
.B2(n_887),
.C1(n_864),
.C2(n_936),
.Y(n_1014)
);

OAI21xp33_ASAP7_75t_SL g1015 ( 
.A1(n_1008),
.A2(n_1006),
.B(n_1010),
.Y(n_1015)
);

NOR4xp25_ASAP7_75t_L g1016 ( 
.A(n_1012),
.B(n_877),
.C(n_874),
.D(n_875),
.Y(n_1016)
);

AOI211xp5_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_917),
.B(n_846),
.C(n_800),
.Y(n_1017)
);

AOI222xp33_ASAP7_75t_L g1018 ( 
.A1(n_1007),
.A2(n_917),
.B1(n_952),
.B2(n_937),
.C1(n_931),
.C2(n_936),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1011),
.A2(n_954),
.B1(n_950),
.B2(n_951),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1010),
.B(n_954),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1011),
.A2(n_917),
.B(n_919),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_1011),
.Y(n_1022)
);

AOI221xp5_ASAP7_75t_L g1023 ( 
.A1(n_1022),
.A2(n_917),
.B1(n_942),
.B2(n_937),
.C(n_931),
.Y(n_1023)
);

AOI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_1015),
.A2(n_954),
.B1(n_919),
.B2(n_881),
.C(n_959),
.Y(n_1024)
);

AOI221xp5_ASAP7_75t_L g1025 ( 
.A1(n_1016),
.A2(n_959),
.B1(n_948),
.B2(n_951),
.C(n_944),
.Y(n_1025)
);

AOI221xp5_ASAP7_75t_L g1026 ( 
.A1(n_1020),
.A2(n_950),
.B1(n_948),
.B2(n_878),
.C(n_886),
.Y(n_1026)
);

AOI211xp5_ASAP7_75t_SL g1027 ( 
.A1(n_1014),
.A2(n_938),
.B(n_933),
.C(n_842),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_1019),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_1018),
.A2(n_878),
.B1(n_886),
.B2(n_846),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1013),
.A2(n_1017),
.B1(n_1021),
.B2(n_957),
.C(n_955),
.Y(n_1030)
);

AOI222xp33_ASAP7_75t_L g1031 ( 
.A1(n_1015),
.A2(n_895),
.B1(n_846),
.B2(n_957),
.C1(n_955),
.C2(n_903),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_SL g1032 ( 
.A(n_1016),
.B(n_895),
.C(n_901),
.Y(n_1032)
);

NOR2x1_ASAP7_75t_L g1033 ( 
.A(n_1028),
.B(n_883),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1030),
.A2(n_786),
.B1(n_846),
.B2(n_941),
.Y(n_1034)
);

NOR2x1_ASAP7_75t_L g1035 ( 
.A(n_1032),
.B(n_883),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1031),
.B(n_957),
.Y(n_1036)
);

NAND4xp75_ASAP7_75t_L g1037 ( 
.A(n_1024),
.B(n_901),
.C(n_927),
.D(n_934),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_L g1038 ( 
.A(n_1027),
.B(n_957),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1026),
.Y(n_1039)
);

OAI322xp33_ASAP7_75t_L g1040 ( 
.A1(n_1039),
.A2(n_1029),
.A3(n_1023),
.B1(n_1025),
.B2(n_955),
.C1(n_902),
.C2(n_934),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_955),
.Y(n_1041)
);

NAND4xp75_ASAP7_75t_L g1042 ( 
.A(n_1035),
.B(n_893),
.C(n_928),
.D(n_902),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1038),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1034),
.A2(n_941),
.B1(n_821),
.B2(n_928),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_SL g1045 ( 
.A1(n_1043),
.A2(n_1036),
.B1(n_1037),
.B2(n_821),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1041),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1040),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1044),
.A2(n_821),
.B1(n_902),
.B2(n_923),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_1047),
.A2(n_1046),
.B1(n_1048),
.B2(n_1045),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1046),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_SL g1051 ( 
.A1(n_1049),
.A2(n_1042),
.B1(n_821),
.B2(n_923),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_1050),
.B(n_940),
.C(n_924),
.Y(n_1052)
);

NAND4xp25_ASAP7_75t_L g1053 ( 
.A(n_1052),
.B(n_216),
.C(n_217),
.D(n_918),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1051),
.A2(n_940),
.B1(n_924),
.B2(n_929),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1053),
.B(n_1054),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1053),
.A2(n_841),
.B(n_940),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1055),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1056),
.A2(n_929),
.B1(n_916),
.B2(n_918),
.Y(n_1058)
);

AOI21xp33_ASAP7_75t_SL g1059 ( 
.A1(n_1057),
.A2(n_1058),
.B(n_841),
.Y(n_1059)
);

INVxp33_ASAP7_75t_SL g1060 ( 
.A(n_1057),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1060),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_R g1062 ( 
.A1(n_1061),
.A2(n_1059),
.B1(n_892),
.B2(n_924),
.C(n_891),
.Y(n_1062)
);

AOI211xp5_ASAP7_75t_L g1063 ( 
.A1(n_1062),
.A2(n_916),
.B(n_908),
.C(n_906),
.Y(n_1063)
);


endmodule