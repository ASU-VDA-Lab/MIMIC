module fake_netlist_1_7733_n_719 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_719);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_719;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g81 ( .A(n_34), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_36), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_23), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_59), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_0), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_43), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_7), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_11), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_56), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_60), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_76), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_24), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_66), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_53), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_16), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_2), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_71), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_33), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_27), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_75), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_11), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_51), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_1), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_54), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_63), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_29), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_28), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_61), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_30), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_49), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_5), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_8), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
INVxp33_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
BUFx5_ASAP7_75t_L g125 ( .A(n_25), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_69), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_18), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_38), .Y(n_128) );
INVxp33_ASAP7_75t_SL g129 ( .A(n_64), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_17), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
CKINVDCx8_ASAP7_75t_R g133 ( .A(n_100), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_125), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_89), .B(n_32), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_113), .B(n_0), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_113), .B(n_1), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_125), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_88), .B(n_91), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_124), .B(n_100), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_88), .B(n_3), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_85), .A2(n_35), .B(n_79), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_106), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_91), .B(n_3), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_106), .Y(n_156) );
NAND3xp33_ASAP7_75t_L g157 ( .A(n_109), .B(n_39), .C(n_78), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_99), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_109), .B(n_4), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_122), .B(n_4), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_108), .B(n_5), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_108), .B(n_6), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_122), .B(n_7), .Y(n_165) );
BUFx8_ASAP7_75t_L g166 ( .A(n_125), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_123), .B(n_8), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_83), .B(n_9), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_105), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_93), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_93), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_123), .B(n_9), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_165), .B(n_110), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_148), .B(n_130), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_166), .B(n_92), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_165), .B(n_128), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_166), .B(n_82), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
INVx4_ASAP7_75t_SL g186 ( .A(n_139), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVx5_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_131), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_135), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_137), .B(n_121), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_151), .B(n_95), .Y(n_194) );
AOI22xp33_ASAP7_75t_SL g195 ( .A1(n_169), .A2(n_120), .B1(n_126), .B2(n_81), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_169), .B(n_129), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_156), .B(n_83), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_158), .B(n_119), .Y(n_203) );
AO22x2_ASAP7_75t_L g204 ( .A1(n_142), .A2(n_128), .B1(n_104), .B2(n_103), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_166), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_135), .Y(n_206) );
NOR2x1_ASAP7_75t_L g207 ( .A(n_142), .B(n_114), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_138), .B(n_119), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_133), .B(n_96), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_138), .B(n_89), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_173), .A2(n_127), .B1(n_107), .B2(n_117), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_156), .B(n_107), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g215 ( .A(n_139), .B(n_84), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_173), .Y(n_216) );
INVx5_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_133), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_135), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_134), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_134), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_139), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_144), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_141), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_144), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_154), .B(n_84), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_147), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_135), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_154), .B(n_110), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_155), .B(n_90), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_147), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_155), .B(n_114), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_136), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_153), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_153), .Y(n_238) );
INVx6_ASAP7_75t_L g239 ( .A(n_139), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_170), .B(n_90), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_204), .A2(n_172), .B1(n_170), .B2(n_162), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_199), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_216), .A2(n_161), .B1(n_167), .B2(n_149), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_199), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_205), .B(n_153), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_204), .A2(n_172), .B1(n_162), .B2(n_164), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_203), .Y(n_247) );
BUFx8_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_176), .A2(n_164), .B1(n_161), .B2(n_167), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g252 ( .A(n_218), .B(n_145), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_211), .Y(n_253) );
AO22x1_ASAP7_75t_L g254 ( .A1(n_180), .A2(n_139), .B1(n_118), .B2(n_145), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g256 ( .A1(n_204), .A2(n_149), .B1(n_160), .B2(n_152), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_193), .B(n_160), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_175), .B(n_152), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_203), .B(n_168), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_204), .A2(n_127), .B1(n_94), .B2(n_112), .C(n_111), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_195), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_214), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_209), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_214), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_214), .B(n_171), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_175), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_199), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_201), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_178), .B(n_116), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_193), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_175), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
NOR2x1p5_ASAP7_75t_L g274 ( .A(n_194), .B(n_112), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_231), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_221), .B(n_111), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_205), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_180), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_196), .B(n_117), .Y(n_280) );
NOR2x1p5_ASAP7_75t_SL g281 ( .A(n_220), .B(n_171), .Y(n_281) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_207), .B(n_157), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_201), .B(n_157), .Y(n_284) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_231), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_179), .B(n_127), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_226), .B(n_171), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_231), .Y(n_289) );
BUFx4f_ASAP7_75t_L g290 ( .A(n_180), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_180), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_180), .A2(n_115), .B1(n_97), .B2(n_101), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_181), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_207), .B(n_163), .Y(n_294) );
BUFx4f_ASAP7_75t_L g295 ( .A(n_180), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_198), .B(n_163), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_228), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_232), .A2(n_163), .B1(n_159), .B2(n_127), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_212), .B(n_159), .Y(n_299) );
OR2x2_ASAP7_75t_SL g300 ( .A(n_240), .B(n_150), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_222), .A2(n_150), .B(n_159), .Y(n_301) );
NAND3xp33_ASAP7_75t_SL g302 ( .A(n_212), .B(n_116), .C(n_97), .Y(n_302) );
CKINVDCx6p67_ASAP7_75t_R g303 ( .A(n_182), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_235), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_233), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_186), .B(n_94), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_233), .B(n_115), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_188), .Y(n_308) );
INVx3_ASAP7_75t_SL g309 ( .A(n_186), .Y(n_309) );
NOR2xp33_ASAP7_75t_R g310 ( .A(n_215), .B(n_10), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_224), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_186), .B(n_101), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_258), .B(n_186), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_244), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_285), .A2(n_215), .B1(n_181), .B2(n_239), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_243), .B(n_181), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
BUFx8_ASAP7_75t_SL g319 ( .A(n_261), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_271), .B(n_189), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_248), .Y(n_322) );
NOR2xp67_ASAP7_75t_L g323 ( .A(n_257), .B(n_10), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_263), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_268), .Y(n_325) );
OR2x6_ASAP7_75t_L g326 ( .A(n_258), .B(n_239), .Y(n_326) );
NOR2x1_ASAP7_75t_R g327 ( .A(n_264), .B(n_239), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_265), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_258), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_260), .A2(n_102), .B(n_103), .C(n_104), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_269), .Y(n_332) );
BUFx4f_ASAP7_75t_SL g333 ( .A(n_248), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_276), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_252), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_243), .B(n_233), .Y(n_336) );
CKINVDCx11_ASAP7_75t_R g337 ( .A(n_303), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_276), .Y(n_338) );
BUFx12f_ASAP7_75t_L g339 ( .A(n_247), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_256), .A2(n_127), .B1(n_238), .B2(n_189), .Y(n_340) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_260), .B(n_200), .C(n_238), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_297), .B(n_197), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_249), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_245), .A2(n_224), .B(n_217), .Y(n_344) );
BUFx10_ASAP7_75t_L g345 ( .A(n_267), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_250), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_253), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_259), .B(n_197), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_259), .B(n_200), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_246), .A2(n_239), .B1(n_227), .B2(n_234), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_256), .A2(n_127), .B1(n_234), .B2(n_229), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_272), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_241), .A2(n_223), .B1(n_229), .B2(n_227), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_246), .A2(n_223), .B1(n_202), .B2(n_237), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_288), .B(n_202), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_262), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_275), .A2(n_217), .B1(n_188), .B2(n_220), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_301), .A2(n_150), .B(n_237), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_302), .A2(n_225), .B(n_102), .C(n_95), .Y(n_360) );
NOR2xp67_ASAP7_75t_L g361 ( .A(n_251), .B(n_12), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_273), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_242), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_242), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_279), .B(n_150), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_310), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_279), .Y(n_367) );
AOI22xp5_ASAP7_75t_SL g368 ( .A1(n_322), .A2(n_304), .B1(n_280), .B2(n_270), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_345), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_315), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_313), .A2(n_241), .B1(n_295), .B2(n_290), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_333), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_342), .A2(n_295), .B1(n_290), .B2(n_292), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_296), .B1(n_291), .B2(n_266), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_318), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_333), .Y(n_376) );
CKINVDCx6p67_ASAP7_75t_R g377 ( .A(n_337), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_353), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_337), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_361), .A2(n_302), .B1(n_274), .B2(n_280), .Y(n_381) );
INVx4_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_345), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_329), .A2(n_291), .B1(n_286), .B2(n_278), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_329), .B(n_277), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_341), .A2(n_282), .B(n_299), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_324), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_343), .A2(n_270), .B1(n_307), .B2(n_298), .C(n_294), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_328), .Y(n_392) );
AOI21xp5_ASAP7_75t_R g393 ( .A1(n_314), .A2(n_312), .B(n_306), .Y(n_393) );
BUFx2_ASAP7_75t_SL g394 ( .A(n_331), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_326), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_366), .A2(n_310), .B1(n_286), .B2(n_277), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_353), .B(n_349), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_356), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_331), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_350), .B(n_284), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_391), .B(n_340), .Y(n_401) );
AO21x2_ASAP7_75t_L g402 ( .A1(n_387), .A2(n_359), .B(n_330), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_398), .B(n_320), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_368), .B(n_334), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_393), .A2(n_352), .B1(n_336), .B2(n_323), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_398), .A2(n_338), .B1(n_339), .B2(n_336), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_396), .A2(n_352), .B1(n_317), .B2(n_354), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_389), .Y(n_408) );
INVx4_ASAP7_75t_L g409 ( .A(n_391), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_381), .A2(n_317), .B1(n_354), .B2(n_330), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_395), .A2(n_339), .B1(n_345), .B2(n_286), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_390), .B(n_360), .C(n_284), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_379), .B(n_357), .C(n_348), .D(n_346), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_372), .B(n_335), .C(n_298), .D(n_355), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_400), .A2(n_284), .B1(n_332), .B2(n_362), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_395), .A2(n_326), .B1(n_365), .B2(n_351), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g417 ( .A1(n_389), .A2(n_364), .B(n_319), .C(n_363), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_397), .B(n_326), .Y(n_418) );
BUFx12f_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_397), .A2(n_365), .B1(n_325), .B2(n_362), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_392), .Y(n_421) );
BUFx12f_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_378), .A2(n_363), .B(n_316), .C(n_325), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_400), .A2(n_332), .B1(n_319), .B2(n_365), .Y(n_425) );
CKINVDCx6p67_ASAP7_75t_R g426 ( .A(n_377), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_370), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_375), .B(n_327), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_374), .A2(n_314), .B1(n_367), .B2(n_300), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_408), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_413), .B(n_392), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_412), .B(n_399), .C(n_382), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_427), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_416), .A2(n_388), .B1(n_371), .B2(n_384), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_427), .Y(n_435) );
AOI322xp5_ASAP7_75t_L g436 ( .A1(n_404), .A2(n_375), .A3(n_385), .B1(n_388), .B2(n_383), .C1(n_369), .C2(n_377), .Y(n_436) );
AO21x2_ASAP7_75t_L g437 ( .A1(n_401), .A2(n_359), .B(n_385), .Y(n_437) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_401), .A2(n_370), .B(n_380), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_421), .B(n_380), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_403), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_407), .A2(n_369), .B1(n_383), .B2(n_373), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_410), .A2(n_254), .B1(n_314), .B2(n_146), .C(n_136), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_415), .B(n_382), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_405), .A2(n_394), .B1(n_399), .B2(n_382), .Y(n_449) );
NOR2x1_ASAP7_75t_SL g450 ( .A(n_420), .B(n_394), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_423), .A2(n_399), .B1(n_391), .B2(n_386), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_415), .B(n_391), .C(n_136), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_425), .B(n_406), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_416), .A2(n_386), .B1(n_391), .B2(n_367), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_411), .A2(n_136), .B(n_143), .C(n_146), .Y(n_456) );
OAI33xp33_ASAP7_75t_L g457 ( .A1(n_417), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_425), .B(n_386), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_418), .B(n_281), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_419), .B(n_15), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
OAI21x1_ASAP7_75t_L g463 ( .A1(n_414), .A2(n_344), .B(n_245), .Y(n_463) );
AOI31xp33_ASAP7_75t_L g464 ( .A1(n_426), .A2(n_312), .A3(n_306), .B(n_19), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_419), .B(n_305), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_422), .A2(n_367), .B1(n_347), .B2(n_255), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_442), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_434), .A2(n_358), .A3(n_255), .B(n_305), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_440), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
OAI31xp33_ASAP7_75t_L g474 ( .A1(n_434), .A2(n_283), .A3(n_19), .B(n_18), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_448), .B(n_20), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_448), .B(n_22), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_430), .B(n_146), .Y(n_477) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_452), .A2(n_283), .B(n_225), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_440), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_433), .Y(n_480) );
INVxp33_ASAP7_75t_SL g481 ( .A(n_466), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_455), .B(n_146), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_146), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_448), .B(n_26), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_433), .B(n_146), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_435), .B(n_143), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_436), .B(n_177), .C(n_174), .D(n_185), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_431), .A2(n_347), .B1(n_367), .B2(n_188), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_435), .B(n_143), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_439), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_452), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_436), .A2(n_136), .B1(n_143), .B2(n_347), .C(n_219), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_439), .B(n_143), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_453), .B(n_143), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_453), .B(n_136), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_458), .A2(n_347), .B1(n_311), .B2(n_217), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_464), .A2(n_192), .B1(n_236), .B2(n_230), .C(n_219), .Y(n_500) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_444), .A2(n_177), .B(n_185), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_454), .A2(n_192), .B(n_206), .C(n_219), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_437), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_443), .A2(n_217), .B1(n_188), .B2(n_311), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_432), .B(n_236), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_438), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_438), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_464), .A2(n_206), .B1(n_183), .B2(n_236), .C(n_230), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_459), .B(n_31), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_41), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_462), .B(n_206), .C(n_184), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_438), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_459), .B(n_42), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_447), .B(n_44), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_446), .B(n_45), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_441), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_441), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_473), .B(n_441), .Y(n_520) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_491), .Y(n_521) );
NAND4xp25_ASAP7_75t_L g522 ( .A(n_474), .B(n_460), .C(n_449), .D(n_465), .Y(n_522) );
NOR3xp33_ASAP7_75t_SL g523 ( .A(n_500), .B(n_457), .C(n_509), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_468), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_473), .B(n_461), .Y(n_526) );
AND3x2_ASAP7_75t_L g527 ( .A(n_471), .B(n_466), .C(n_462), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_487), .B(n_454), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_487), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_481), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g533 ( .A1(n_482), .A2(n_465), .A3(n_432), .B1(n_461), .B2(n_457), .B3(n_449), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_511), .B(n_461), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_511), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_483), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_483), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_496), .B(n_459), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_496), .B(n_459), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_498), .B(n_450), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_498), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_477), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_518), .B(n_450), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g545 ( .A1(n_474), .A2(n_451), .B(n_456), .C(n_445), .Y(n_545) );
OAI31xp33_ASAP7_75t_SL g546 ( .A1(n_494), .A2(n_456), .A3(n_451), .B(n_445), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_516), .A2(n_467), .B1(n_463), .B2(n_236), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_518), .B(n_463), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_516), .B(n_463), .Y(n_549) );
OAI31xp33_ASAP7_75t_L g550 ( .A1(n_512), .A2(n_46), .A3(n_47), .B(n_52), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_517), .Y(n_551) );
OAI33xp33_ASAP7_75t_L g552 ( .A1(n_517), .A2(n_187), .A3(n_213), .B1(n_210), .B2(n_191), .B3(n_190), .Y(n_552) );
OAI21xp33_ASAP7_75t_L g553 ( .A1(n_492), .A2(n_206), .B(n_236), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_470), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_470), .B(n_55), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_519), .B(n_58), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_510), .B(n_62), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_495), .B(n_65), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_470), .Y(n_559) );
AND3x1_ASAP7_75t_L g560 ( .A(n_502), .B(n_67), .C(n_68), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_519), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_502), .B(n_206), .C(n_192), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_472), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_472), .B(n_72), .Y(n_564) );
OAI33xp33_ASAP7_75t_L g565 ( .A1(n_503), .A2(n_191), .A3(n_213), .B1(n_210), .B2(n_174), .B3(n_190), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_503), .B(n_73), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_472), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_495), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_475), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_479), .B(n_77), .Y(n_570) );
INVx3_ASAP7_75t_L g571 ( .A(n_479), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_479), .B(n_80), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_475), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_475), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_479), .B(n_187), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_475), .Y(n_577) );
AOI211x1_ASAP7_75t_SL g578 ( .A1(n_522), .A2(n_515), .B(n_489), .C(n_488), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_532), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_521), .B(n_504), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_536), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_525), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_537), .B(n_504), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_538), .B(n_514), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_533), .B(n_484), .Y(n_586) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_545), .A2(n_484), .A3(n_476), .B(n_469), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_574), .A2(n_476), .B1(n_484), .B2(n_513), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_524), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
NOR2x1_ASAP7_75t_R g591 ( .A(n_555), .B(n_476), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_552), .B(n_484), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_531), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_561), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_539), .B(n_508), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_541), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_520), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_520), .Y(n_598) );
NOR2xp33_ASAP7_75t_SL g599 ( .A(n_550), .B(n_469), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_539), .B(n_508), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_551), .B(n_486), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_526), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_526), .B(n_486), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_568), .B(n_485), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_543), .Y(n_606) );
NAND2xp33_ASAP7_75t_SL g607 ( .A(n_523), .B(n_478), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_544), .B(n_508), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_542), .B(n_485), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_528), .B(n_508), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_540), .B(n_506), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_540), .B(n_506), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_562), .A2(n_513), .B(n_478), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_534), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_544), .B(n_507), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_554), .B(n_490), .Y(n_616) );
NOR2xp33_ASAP7_75t_R g617 ( .A(n_527), .B(n_499), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_530), .B(n_501), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_559), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_563), .B(n_497), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_567), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_565), .B(n_505), .C(n_497), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_576), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_527), .B(n_501), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_546), .B(n_493), .C(n_308), .D(n_478), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_541), .B(n_493), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_582), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_595), .B(n_549), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_600), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_606), .B(n_548), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_590), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_587), .B(n_560), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_617), .A2(n_523), .B(n_547), .C(n_557), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_589), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_592), .B(n_564), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_614), .B(n_577), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_588), .B(n_553), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_583), .B(n_569), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_597), .B(n_573), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_601), .B(n_535), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_589), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_599), .A2(n_557), .B1(n_566), .B2(n_558), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_627), .B(n_571), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_592), .B(n_572), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_608), .B(n_598), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_579), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_619), .B(n_571), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_593), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_581), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_588), .B(n_571), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_596), .A2(n_570), .B1(n_535), .B2(n_556), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_618), .B(n_535), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_621), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_608), .B(n_556), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_624), .Y(n_657) );
XOR2x2_ASAP7_75t_L g658 ( .A(n_580), .B(n_575), .Y(n_658) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_623), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_615), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_615), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_625), .B(n_183), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_586), .B(n_183), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_584), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_585), .Y(n_665) );
AOI221xp5_ASAP7_75t_SL g666 ( .A1(n_586), .A2(n_183), .B1(n_184), .B2(n_192), .C(n_230), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_611), .A2(n_183), .B1(n_184), .B2(n_230), .Y(n_667) );
INVx1_ASAP7_75t_SL g668 ( .A(n_604), .Y(n_668) );
AOI21xp5_ASAP7_75t_SL g669 ( .A1(n_591), .A2(n_184), .B(n_230), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_607), .A2(n_184), .B1(n_192), .B2(n_219), .C1(n_217), .C2(n_188), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_602), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_623), .A2(n_293), .B(n_308), .C(n_625), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_616), .Y(n_673) );
OAI22xp5_ASAP7_75t_SL g674 ( .A1(n_617), .A2(n_293), .B1(n_610), .B2(n_578), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_612), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_610), .B(n_293), .Y(n_676) );
NOR4xp25_ASAP7_75t_L g677 ( .A(n_626), .B(n_605), .C(n_609), .D(n_607), .Y(n_677) );
OAI31xp33_ASAP7_75t_L g678 ( .A1(n_613), .A2(n_620), .A3(n_622), .B(n_594), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_622), .A2(n_586), .B1(n_525), .B2(n_583), .C(n_607), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_587), .A2(n_617), .B(n_532), .C(n_607), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_606), .B(n_603), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_587), .A2(n_453), .B1(n_522), .B2(n_586), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_634), .A2(n_669), .B(n_680), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_660), .A2(n_637), .B1(n_661), .B2(n_675), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_677), .A2(n_679), .B(n_646), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_643), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_658), .B(n_682), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_678), .A2(n_682), .B(n_635), .C(n_644), .Y(n_688) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_672), .A2(n_660), .B(n_661), .C(n_639), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_668), .A2(n_651), .A3(n_659), .B1(n_671), .B2(n_647), .C1(n_652), .C2(n_629), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_665), .B(n_664), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_674), .A2(n_673), .B1(n_637), .B2(n_660), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_681), .A2(n_636), .B1(n_628), .B2(n_650), .C(n_633), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_636), .Y(n_694) );
AO22x2_ASAP7_75t_L g695 ( .A1(n_662), .A2(n_655), .B1(n_631), .B2(n_630), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_657), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_SL g697 ( .A1(n_689), .A2(n_662), .B(n_658), .C(n_653), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_686), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_688), .A2(n_637), .B1(n_640), .B2(n_647), .Y(n_699) );
OAI211xp5_ASAP7_75t_SL g700 ( .A1(n_683), .A2(n_663), .B(n_670), .C(n_667), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_687), .A2(n_630), .B(n_631), .Y(n_701) );
NAND3x1_ASAP7_75t_SL g702 ( .A(n_685), .B(n_666), .C(n_656), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_695), .A2(n_657), .B(n_649), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_695), .A2(n_632), .B1(n_648), .B2(n_641), .C(n_638), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_698), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_701), .A2(n_691), .B1(n_690), .B2(n_694), .Y(n_706) );
NOR2x1p5_ASAP7_75t_L g707 ( .A(n_697), .B(n_696), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_699), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_700), .B(n_692), .C(n_693), .D(n_676), .Y(n_709) );
OAI222xp33_ASAP7_75t_L g710 ( .A1(n_706), .A2(n_703), .B1(n_684), .B2(n_702), .C1(n_704), .C2(n_654), .Y(n_710) );
OAI221xp5_ASAP7_75t_R g711 ( .A1(n_707), .A2(n_642), .B1(n_629), .B2(n_656), .C(n_645), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_705), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_712), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_712), .A2(n_709), .B1(n_708), .B2(n_676), .C(n_654), .Y(n_714) );
INVx3_ASAP7_75t_L g715 ( .A(n_713), .Y(n_715) );
INVx4_ASAP7_75t_L g716 ( .A(n_714), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_711), .B1(n_710), .B2(n_642), .Y(n_717) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_717), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_716), .B1(n_715), .B2(n_645), .Y(n_719) );
endmodule