module real_aes_16809_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1595;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g921 ( .A(n_0), .B(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g650 ( .A(n_1), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g1368 ( .A1(n_2), .A2(n_297), .B1(n_599), .B2(n_626), .Y(n_1368) );
OAI22xp33_ASAP7_75t_SL g1378 ( .A1(n_2), .A2(n_297), .B1(n_476), .B2(n_1267), .Y(n_1378) );
INVx1_ASAP7_75t_L g542 ( .A(n_3), .Y(n_542) );
INVx1_ASAP7_75t_L g345 ( .A(n_4), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_4), .B(n_355), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_5), .A2(n_239), .B1(n_430), .B2(n_434), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_5), .A2(n_179), .B1(n_501), .B2(n_504), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g1618 ( .A(n_6), .Y(n_1618) );
OAI22xp33_ASAP7_75t_SL g1630 ( .A1(n_7), .A2(n_320), .B1(n_599), .B2(n_1631), .Y(n_1630) );
OAI22xp33_ASAP7_75t_L g1639 ( .A1(n_7), .A2(n_162), .B1(n_476), .B2(n_571), .Y(n_1639) );
INVx1_ASAP7_75t_L g1285 ( .A(n_8), .Y(n_1285) );
INVx1_ASAP7_75t_L g413 ( .A(n_9), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_9), .A2(n_239), .B1(n_504), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g666 ( .A(n_10), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_11), .A2(n_190), .B1(n_1400), .B2(n_1414), .Y(n_1426) );
CKINVDCx5p33_ASAP7_75t_R g1202 ( .A(n_12), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_13), .A2(n_85), .B1(n_1400), .B2(n_1402), .Y(n_1418) );
CKINVDCx5p33_ASAP7_75t_R g1221 ( .A(n_14), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_15), .A2(n_313), .B1(n_1392), .B2(n_1397), .Y(n_1515) );
OAI22xp33_ASAP7_75t_L g1375 ( .A1(n_16), .A2(n_275), .B1(n_850), .B2(n_1376), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_16), .A2(n_275), .B1(n_462), .B2(n_468), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_17), .A2(n_292), .B1(n_756), .B2(n_1160), .Y(n_1177) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_17), .A2(n_292), .B1(n_745), .B2(n_1121), .Y(n_1180) );
INVx2_ASAP7_75t_L g456 ( .A(n_18), .Y(n_456) );
INVx1_ASAP7_75t_L g999 ( .A(n_19), .Y(n_999) );
INVx1_ASAP7_75t_L g995 ( .A(n_20), .Y(n_995) );
INVx1_ASAP7_75t_L g1087 ( .A(n_21), .Y(n_1087) );
INVx1_ASAP7_75t_L g1058 ( .A(n_22), .Y(n_1058) );
INVx1_ASAP7_75t_L g1331 ( .A(n_23), .Y(n_1331) );
INVx1_ASAP7_75t_L g1280 ( .A(n_24), .Y(n_1280) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_25), .A2(n_79), .B1(n_687), .B2(n_978), .C(n_980), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_25), .A2(n_41), .B1(n_1028), .B2(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g720 ( .A(n_26), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g1423 ( .A1(n_27), .A2(n_200), .B1(n_1392), .B2(n_1397), .Y(n_1423) );
INVx1_ASAP7_75t_L g875 ( .A(n_28), .Y(n_875) );
INVx1_ASAP7_75t_L g1082 ( .A(n_29), .Y(n_1082) );
OAI211xp5_ASAP7_75t_L g1108 ( .A1(n_30), .A2(n_610), .B(n_1109), .C(n_1112), .Y(n_1108) );
INVx1_ASAP7_75t_L g1119 ( .A(n_30), .Y(n_1119) );
INVx1_ASAP7_75t_L g766 ( .A(n_31), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_32), .A2(n_78), .B1(n_462), .B2(n_571), .C(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g595 ( .A(n_32), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_33), .A2(n_296), .B1(n_597), .B2(n_850), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_33), .A2(n_296), .B1(n_462), .B2(n_468), .Y(n_1273) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_34), .Y(n_340) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_34), .B(n_338), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_35), .A2(n_174), .B1(n_1400), .B2(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g934 ( .A(n_36), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_37), .A2(n_187), .B1(n_1400), .B2(n_1402), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_38), .Y(n_832) );
INVx1_ASAP7_75t_L g1141 ( .A(n_39), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_40), .A2(n_167), .B1(n_734), .B2(n_735), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_40), .A2(n_167), .B1(n_347), .B2(n_367), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_41), .A2(n_66), .B1(n_687), .B2(n_978), .C(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1320 ( .A(n_42), .Y(n_1320) );
OAI22xp33_ASAP7_75t_L g1264 ( .A1(n_43), .A2(n_251), .B1(n_599), .B2(n_600), .Y(n_1264) );
OAI22xp33_ASAP7_75t_SL g1266 ( .A1(n_43), .A2(n_251), .B1(n_476), .B2(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g899 ( .A(n_44), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_44), .A2(n_324), .B1(n_621), .B2(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g743 ( .A(n_45), .Y(n_743) );
OAI211xp5_ASAP7_75t_L g751 ( .A1(n_45), .A2(n_610), .B(n_752), .C(n_753), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g1408 ( .A1(n_46), .A2(n_151), .B1(n_1400), .B2(n_1402), .Y(n_1408) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_47), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_48), .Y(n_404) );
INVx1_ASAP7_75t_L g937 ( .A(n_49), .Y(n_937) );
INVx1_ASAP7_75t_L g1356 ( .A(n_50), .Y(n_1356) );
INVx1_ASAP7_75t_L g989 ( .A(n_51), .Y(n_989) );
AOI22xp33_ASAP7_75t_SL g1022 ( .A1(n_51), .A2(n_244), .B1(n_434), .B2(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g546 ( .A(n_52), .Y(n_546) );
INVx1_ASAP7_75t_L g867 ( .A(n_53), .Y(n_867) );
XNOR2xp5_ASAP7_75t_L g606 ( .A(n_54), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g1065 ( .A(n_55), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_56), .B(n_455), .Y(n_574) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_56), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g1304 ( .A1(n_57), .A2(n_816), .B(n_1182), .C(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1313 ( .A(n_57), .Y(n_1313) );
OAI211xp5_ASAP7_75t_L g1626 ( .A1(n_58), .A2(n_558), .B(n_583), .C(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1638 ( .A(n_58), .Y(n_1638) );
INVx1_ASAP7_75t_L g718 ( .A(n_59), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g1610 ( .A(n_60), .Y(n_1610) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_61), .A2(n_164), .B1(n_380), .B2(n_384), .C1(n_388), .C2(n_389), .Y(n_379) );
OAI222xp33_ASAP7_75t_L g443 ( .A1(n_61), .A2(n_164), .B1(n_207), .B2(n_444), .C1(n_452), .C2(n_458), .Y(n_443) );
INVx1_ASAP7_75t_L g1284 ( .A(n_62), .Y(n_1284) );
OAI22xp33_ASAP7_75t_L g1161 ( .A1(n_63), .A2(n_276), .B1(n_347), .B2(n_626), .Y(n_1161) );
OAI22xp33_ASAP7_75t_L g1163 ( .A1(n_63), .A2(n_276), .B1(n_644), .B2(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1111 ( .A(n_64), .Y(n_1111) );
OAI211xp5_ASAP7_75t_L g1117 ( .A1(n_64), .A2(n_633), .B(n_634), .C(n_1118), .Y(n_1117) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_65), .A2(n_169), .B1(n_476), .B2(n_578), .Y(n_577) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_65), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_66), .A2(n_79), .B1(n_425), .B2(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1355 ( .A(n_67), .Y(n_1355) );
INVx1_ASAP7_75t_L g1330 ( .A(n_68), .Y(n_1330) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_69), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_70), .A2(n_156), .B1(n_745), .B2(n_746), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_70), .A2(n_156), .B1(n_621), .B2(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g1326 ( .A(n_71), .Y(n_1326) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_72), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g1258 ( .A1(n_73), .A2(n_583), .B(n_1259), .C(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1270 ( .A(n_73), .Y(n_1270) );
INVx1_ASAP7_75t_L g619 ( .A(n_74), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_74), .A2(n_633), .B(n_634), .C(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g544 ( .A(n_75), .Y(n_544) );
INVx1_ASAP7_75t_L g932 ( .A(n_76), .Y(n_932) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_77), .B(n_821), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_78), .A2(n_169), .B1(n_599), .B2(n_600), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_80), .A2(n_176), .B1(n_462), .B2(n_476), .Y(n_992) );
INVx1_ASAP7_75t_L g1005 ( .A(n_80), .Y(n_1005) );
INVx1_ASAP7_75t_L g1089 ( .A(n_81), .Y(n_1089) );
INVx1_ASAP7_75t_L g808 ( .A(n_82), .Y(n_808) );
OAI211xp5_ASAP7_75t_L g813 ( .A1(n_82), .A2(n_814), .B(n_816), .C(n_817), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_83), .A2(n_250), .B1(n_597), .B2(n_599), .Y(n_1238) );
OAI22xp5_ASAP7_75t_SL g1246 ( .A1(n_83), .A2(n_117), .B1(n_468), .B2(n_476), .Y(n_1246) );
INVx1_ASAP7_75t_L g576 ( .A(n_84), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_86), .Y(n_1241) );
INVx1_ASAP7_75t_L g1307 ( .A(n_87), .Y(n_1307) );
OAI211xp5_ASAP7_75t_L g1311 ( .A1(n_87), .A2(n_409), .B(n_613), .C(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1288 ( .A(n_88), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g1220 ( .A(n_89), .Y(n_1220) );
OAI22xp33_ASAP7_75t_L g1107 ( .A1(n_90), .A2(n_147), .B1(n_347), .B2(n_600), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_90), .A2(n_147), .B1(n_642), .B2(n_735), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g1609 ( .A(n_91), .Y(n_1609) );
INVx1_ASAP7_75t_L g1000 ( .A(n_92), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g1391 ( .A1(n_93), .A2(n_199), .B1(n_1392), .B2(n_1397), .Y(n_1391) );
XOR2xp5_ASAP7_75t_L g1604 ( .A(n_93), .B(n_1605), .Y(n_1604) );
AOI22xp33_ASAP7_75t_L g1643 ( .A1(n_93), .A2(n_1644), .B1(n_1647), .B2(n_1651), .Y(n_1643) );
INVx1_ASAP7_75t_L g1348 ( .A(n_94), .Y(n_1348) );
INVx1_ASAP7_75t_L g935 ( .A(n_95), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_96), .Y(n_835) );
INVx1_ASAP7_75t_L g1325 ( .A(n_97), .Y(n_1325) );
CKINVDCx5p33_ASAP7_75t_R g1227 ( .A(n_98), .Y(n_1227) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_99), .A2(n_131), .B1(n_599), .B2(n_626), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_99), .A2(n_115), .B1(n_476), .B2(n_745), .Y(n_963) );
INVx1_ASAP7_75t_L g928 ( .A(n_100), .Y(n_928) );
INVx1_ASAP7_75t_L g1262 ( .A(n_101), .Y(n_1262) );
INVx1_ASAP7_75t_L g939 ( .A(n_102), .Y(n_939) );
INVx1_ASAP7_75t_L g1147 ( .A(n_103), .Y(n_1147) );
OAI211xp5_ASAP7_75t_L g803 ( .A1(n_104), .A2(n_583), .B(n_804), .C(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g818 ( .A(n_104), .Y(n_818) );
INVx1_ASAP7_75t_L g338 ( .A(n_105), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_106), .A2(n_272), .B1(n_622), .B2(n_626), .Y(n_810) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_106), .A2(n_143), .B1(n_462), .B2(n_468), .Y(n_819) );
XOR2xp5_ASAP7_75t_L g363 ( .A(n_107), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g655 ( .A(n_108), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_109), .Y(n_957) );
INVx1_ASAP7_75t_L g1135 ( .A(n_110), .Y(n_1135) );
AOI22xp5_ASAP7_75t_L g1412 ( .A1(n_111), .A2(n_291), .B1(n_1392), .B2(n_1397), .Y(n_1412) );
INVx1_ASAP7_75t_L g1359 ( .A(n_112), .Y(n_1359) );
INVx1_ASAP7_75t_L g1306 ( .A(n_113), .Y(n_1306) );
INVx1_ASAP7_75t_L g1061 ( .A(n_114), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_115), .A2(n_202), .B1(n_621), .B2(n_960), .Y(n_959) );
OAI22xp33_ASAP7_75t_SL g1243 ( .A1(n_116), .A2(n_117), .B1(n_600), .B2(n_850), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_116), .A2(n_123), .B1(n_1251), .B2(n_1252), .Y(n_1250) );
INVx1_ASAP7_75t_L g1064 ( .A(n_118), .Y(n_1064) );
INVx1_ASAP7_75t_L g1371 ( .A(n_119), .Y(n_1371) );
AOI22xp5_ASAP7_75t_L g1422 ( .A1(n_120), .A2(n_203), .B1(n_1400), .B2(n_1402), .Y(n_1422) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_121), .Y(n_1198) );
INVx1_ASAP7_75t_L g716 ( .A(n_122), .Y(n_716) );
INVx1_ASAP7_75t_L g1242 ( .A(n_123), .Y(n_1242) );
INVx1_ASAP7_75t_L g1323 ( .A(n_124), .Y(n_1323) );
INVx1_ASAP7_75t_L g1062 ( .A(n_125), .Y(n_1062) );
AOI31xp33_ASAP7_75t_L g974 ( .A1(n_126), .A2(n_975), .A3(n_991), .B(n_1003), .Y(n_974) );
NAND2xp33_ASAP7_75t_SL g1020 ( .A(n_126), .B(n_1021), .Y(n_1020) );
INVxp67_ASAP7_75t_SL g1033 ( .A(n_126), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_127), .A2(n_213), .B1(n_1392), .B2(n_1397), .Y(n_1427) );
INVx1_ASAP7_75t_L g1084 ( .A(n_128), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_129), .A2(n_170), .B1(n_626), .B2(n_850), .Y(n_849) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_129), .A2(n_161), .B1(n_462), .B2(n_468), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_130), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_131), .A2(n_202), .B1(n_644), .B2(n_970), .Y(n_969) );
CKINVDCx5p33_ASAP7_75t_R g1201 ( .A(n_132), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_133), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_134), .Y(n_1224) );
OAI22xp33_ASAP7_75t_L g1308 ( .A1(n_135), .A2(n_146), .B1(n_1187), .B2(n_1309), .Y(n_1308) );
OAI22xp33_ASAP7_75t_L g1315 ( .A1(n_135), .A2(n_146), .B1(n_599), .B2(n_626), .Y(n_1315) );
INVx1_ASAP7_75t_L g1350 ( .A(n_136), .Y(n_1350) );
INVx1_ASAP7_75t_L g1091 ( .A(n_137), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g1612 ( .A(n_138), .Y(n_1612) );
OAI211xp5_ASAP7_75t_L g1154 ( .A1(n_139), .A2(n_752), .B(n_1155), .C(n_1156), .Y(n_1154) );
INVx1_ASAP7_75t_L g1167 ( .A(n_139), .Y(n_1167) );
INVx1_ASAP7_75t_L g930 ( .A(n_140), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_141), .Y(n_678) );
INVx1_ASAP7_75t_L g1157 ( .A(n_142), .Y(n_1157) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_143), .A2(n_254), .B1(n_599), .B2(n_624), .Y(n_809) );
INVx1_ASAP7_75t_L g847 ( .A(n_144), .Y(n_847) );
OAI211xp5_ASAP7_75t_L g853 ( .A1(n_144), .A2(n_814), .B(n_816), .C(n_854), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_145), .Y(n_772) );
INVx1_ASAP7_75t_L g540 ( .A(n_148), .Y(n_540) );
INVx1_ASAP7_75t_L g1059 ( .A(n_149), .Y(n_1059) );
INVx1_ASAP7_75t_L g618 ( .A(n_150), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_152), .A2(n_268), .B1(n_756), .B2(n_1160), .Y(n_1159) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_152), .A2(n_268), .B1(n_745), .B2(n_746), .Y(n_1168) );
OAI211xp5_ASAP7_75t_L g844 ( .A1(n_153), .A2(n_583), .B(n_804), .C(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g855 ( .A(n_153), .Y(n_855) );
INVx1_ASAP7_75t_L g1322 ( .A(n_154), .Y(n_1322) );
CKINVDCx5p33_ASAP7_75t_R g1615 ( .A(n_155), .Y(n_1615) );
INVx1_ASAP7_75t_L g1146 ( .A(n_157), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_158), .A2(n_237), .B1(n_621), .B2(n_623), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_158), .A2(n_237), .B1(n_630), .B2(n_631), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_159), .A2(n_161), .B1(n_599), .B2(n_624), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_159), .A2(n_170), .B1(n_476), .B2(n_571), .Y(n_852) );
INVx1_ASAP7_75t_L g675 ( .A(n_160), .Y(n_675) );
OAI22xp33_ASAP7_75t_SL g1632 ( .A1(n_162), .A2(n_279), .B1(n_622), .B2(n_626), .Y(n_1632) );
INVx1_ASAP7_75t_L g1130 ( .A(n_163), .Y(n_1130) );
INVx1_ASAP7_75t_L g1055 ( .A(n_165), .Y(n_1055) );
INVx2_ASAP7_75t_L g1395 ( .A(n_166), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_166), .B(n_1396), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_166), .B(n_274), .Y(n_1403) );
AO22x2_ASAP7_75t_L g1342 ( .A1(n_168), .A2(n_1343), .B1(n_1383), .B2(n_1384), .Y(n_1342) );
INVx1_ASAP7_75t_L g1383 ( .A(n_168), .Y(n_1383) );
AOI22xp5_ASAP7_75t_L g1407 ( .A1(n_168), .A2(n_253), .B1(n_1392), .B2(n_1397), .Y(n_1407) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_171), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_172), .Y(n_1226) );
INVx1_ASAP7_75t_L g665 ( .A(n_173), .Y(n_665) );
INVx1_ASAP7_75t_L g705 ( .A(n_175), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_176), .A2(n_259), .B1(n_597), .B2(n_850), .Y(n_1009) );
INVx1_ASAP7_75t_L g958 ( .A(n_177), .Y(n_958) );
OAI211xp5_ASAP7_75t_L g964 ( .A1(n_177), .A2(n_816), .B(n_965), .C(n_966), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_178), .A2(n_282), .B1(n_1400), .B2(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g419 ( .A(n_179), .Y(n_419) );
XOR2xp5_ASAP7_75t_L g524 ( .A(n_180), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g902 ( .A(n_181), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g917 ( .A1(n_181), .A2(n_215), .B1(n_599), .B2(n_626), .Y(n_917) );
XNOR2x2_ASAP7_75t_L g1076 ( .A(n_182), .B(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g531 ( .A(n_183), .Y(n_531) );
INVx1_ASAP7_75t_L g1042 ( .A(n_184), .Y(n_1042) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_185), .Y(n_781) );
INVx1_ASAP7_75t_L g1261 ( .A(n_186), .Y(n_1261) );
XOR2x2_ASAP7_75t_L g1255 ( .A(n_188), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g702 ( .A(n_189), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_191), .A2(n_367), .B(n_373), .C(n_393), .Y(n_366) );
INVx1_ASAP7_75t_L g477 ( .A(n_191), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_192), .Y(n_1174) );
INVx1_ASAP7_75t_L g1136 ( .A(n_193), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g1303 ( .A1(n_194), .A2(n_216), .B1(n_745), .B2(n_970), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1314 ( .A1(n_194), .A2(n_216), .B1(n_621), .B2(n_911), .Y(n_1314) );
INVx1_ASAP7_75t_L g534 ( .A(n_195), .Y(n_534) );
INVx2_ASAP7_75t_L g486 ( .A(n_196), .Y(n_486) );
INVx1_ASAP7_75t_L g514 ( .A(n_196), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_197), .Y(n_773) );
XOR2xp5_ASAP7_75t_L g696 ( .A(n_198), .B(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g1038 ( .A1(n_201), .A2(n_258), .B1(n_597), .B2(n_850), .Y(n_1038) );
OAI22xp5_ASAP7_75t_SL g1045 ( .A1(n_201), .A2(n_229), .B1(n_462), .B2(n_476), .Y(n_1045) );
INVx1_ASAP7_75t_L g877 ( .A(n_204), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_205), .A2(n_285), .B1(n_1392), .B2(n_1397), .Y(n_1417) );
INVx1_ASAP7_75t_L g387 ( .A(n_206), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_206), .A2(n_234), .B1(n_462), .B2(n_468), .Y(n_461) );
INVx1_ASAP7_75t_L g375 ( .A(n_207), .Y(n_375) );
INVx1_ASAP7_75t_L g894 ( .A(n_208), .Y(n_894) );
OA211x2_ASAP7_75t_L g912 ( .A1(n_208), .A2(n_613), .B(n_658), .C(n_913), .Y(n_912) );
BUFx3_ASAP7_75t_L g451 ( .A(n_209), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_210), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_211), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_212), .Y(n_1199) );
OAI22xp5_ASAP7_75t_SL g860 ( .A1(n_213), .A2(n_861), .B1(n_908), .B2(n_919), .Y(n_860) );
NAND4xp25_ASAP7_75t_L g861 ( .A(n_213), .B(n_862), .C(n_879), .D(n_888), .Y(n_861) );
XOR2xp5_ASAP7_75t_L g1125 ( .A(n_214), .B(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g898 ( .A(n_215), .Y(n_898) );
OA22x2_ASAP7_75t_L g1300 ( .A1(n_217), .A2(n_1301), .B1(n_1339), .B2(n_1340), .Y(n_1300) );
INVxp67_ASAP7_75t_L g1340 ( .A(n_217), .Y(n_1340) );
INVx1_ASAP7_75t_L g1176 ( .A(n_218), .Y(n_1176) );
OAI211xp5_ASAP7_75t_L g1181 ( .A1(n_218), .A2(n_816), .B(n_1182), .C(n_1184), .Y(n_1181) );
INVx1_ASAP7_75t_L g402 ( .A(n_219), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_219), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g1372 ( .A(n_220), .Y(n_1372) );
INVx1_ASAP7_75t_L g1132 ( .A(n_221), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_222), .Y(n_829) );
INVx1_ASAP7_75t_L g870 ( .A(n_223), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_224), .Y(n_777) );
INVx1_ASAP7_75t_L g714 ( .A(n_225), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_226), .A2(n_294), .B1(n_347), .B2(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_226), .A2(n_294), .B1(n_642), .B2(n_644), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g1399 ( .A1(n_227), .A2(n_247), .B1(n_1400), .B2(n_1402), .Y(n_1399) );
INVx1_ASAP7_75t_L g1041 ( .A(n_228), .Y(n_1041) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_229), .A2(n_261), .B1(n_599), .B2(n_600), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g1196 ( .A(n_230), .Y(n_1196) );
INVx1_ASAP7_75t_L g1347 ( .A(n_231), .Y(n_1347) );
INVx1_ASAP7_75t_L g657 ( .A(n_232), .Y(n_657) );
XOR2xp5_ASAP7_75t_L g1215 ( .A(n_233), .B(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g399 ( .A(n_234), .Y(n_399) );
INVx1_ASAP7_75t_L g1281 ( .A(n_235), .Y(n_1281) );
BUFx3_ASAP7_75t_L g355 ( .A(n_236), .Y(n_355) );
INVx1_ASAP7_75t_L g370 ( .A(n_236), .Y(n_370) );
INVx1_ASAP7_75t_L g1110 ( .A(n_238), .Y(n_1110) );
INVx1_ASAP7_75t_L g530 ( .A(n_240), .Y(n_530) );
INVx1_ASAP7_75t_L g893 ( .A(n_241), .Y(n_893) );
INVx1_ASAP7_75t_L g878 ( .A(n_242), .Y(n_878) );
INVx1_ASAP7_75t_L g1277 ( .A(n_243), .Y(n_1277) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_244), .A2(n_264), .B1(n_522), .B2(n_896), .Y(n_976) );
INVx1_ASAP7_75t_L g1094 ( .A(n_245), .Y(n_1094) );
INVx1_ASAP7_75t_L g701 ( .A(n_246), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_248), .A2(n_583), .B(n_658), .C(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1050 ( .A(n_248), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1613 ( .A(n_249), .Y(n_1613) );
NOR2xp33_ASAP7_75t_L g1245 ( .A(n_250), .B(n_462), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_252), .Y(n_1229) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_254), .A2(n_272), .B1(n_476), .B2(n_571), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g1616 ( .A(n_255), .Y(n_1616) );
INVx1_ASAP7_75t_L g874 ( .A(n_256), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_257), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_258), .A2(n_261), .B1(n_468), .B2(n_571), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_259), .A2(n_298), .B1(n_468), .B2(n_571), .Y(n_1001) );
INVx1_ASAP7_75t_L g449 ( .A(n_260), .Y(n_449) );
INVx1_ASAP7_75t_L g467 ( .A(n_260), .Y(n_467) );
INVx1_ASAP7_75t_L g1093 ( .A(n_262), .Y(n_1093) );
INVx1_ASAP7_75t_L g1086 ( .A(n_263), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_264), .A2(n_300), .B1(n_425), .B2(n_1025), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_265), .A2(n_314), .B1(n_621), .B2(n_911), .Y(n_1113) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_265), .A2(n_314), .B1(n_745), .B2(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g871 ( .A(n_266), .Y(n_871) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_267), .A2(n_634), .B(n_737), .C(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g754 ( .A(n_267), .Y(n_754) );
INVx1_ASAP7_75t_L g1628 ( .A(n_269), .Y(n_1628) );
OAI211xp5_ASAP7_75t_SL g1635 ( .A1(n_269), .A2(n_634), .B(n_1636), .C(n_1637), .Y(n_1635) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_270), .A2(n_271), .B1(n_347), .B2(n_626), .Y(n_1178) );
OAI22xp33_ASAP7_75t_L g1186 ( .A1(n_270), .A2(n_271), .B1(n_644), .B2(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g533 ( .A(n_273), .Y(n_533) );
INVx1_ASAP7_75t_L g1396 ( .A(n_274), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_274), .B(n_1395), .Y(n_1401) );
INVx1_ASAP7_75t_L g1278 ( .A(n_277), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_278), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g1634 ( .A1(n_279), .A2(n_320), .B1(n_462), .B2(n_468), .Y(n_1634) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_280), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_281), .A2(n_319), .B1(n_1392), .B2(n_1397), .Y(n_1433) );
INVx1_ASAP7_75t_L g1287 ( .A(n_283), .Y(n_1287) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_284), .Y(n_846) );
INVx1_ASAP7_75t_L g1358 ( .A(n_286), .Y(n_1358) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_287), .Y(n_422) );
OAI211xp5_ASAP7_75t_SL g1239 ( .A1(n_288), .A2(n_558), .B(n_583), .C(n_1240), .Y(n_1239) );
OAI211xp5_ASAP7_75t_SL g1247 ( .A1(n_288), .A2(n_634), .B(n_1248), .C(n_1249), .Y(n_1247) );
INVx1_ASAP7_75t_L g1056 ( .A(n_289), .Y(n_1056) );
INVx1_ASAP7_75t_L g575 ( .A(n_290), .Y(n_575) );
XOR2x2_ASAP7_75t_L g1035 ( .A(n_291), .B(n_1036), .Y(n_1035) );
OAI211xp5_ASAP7_75t_L g1172 ( .A1(n_293), .A2(n_613), .B(n_1155), .C(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1185 ( .A(n_293), .Y(n_1185) );
OAI211xp5_ASAP7_75t_L g954 ( .A1(n_295), .A2(n_613), .B(n_955), .C(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g968 ( .A(n_295), .Y(n_968) );
INVxp67_ASAP7_75t_SL g1007 ( .A(n_298), .Y(n_1007) );
INVx1_ASAP7_75t_L g1158 ( .A(n_299), .Y(n_1158) );
OAI211xp5_ASAP7_75t_L g1165 ( .A1(n_299), .A2(n_816), .B(n_945), .C(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g987 ( .A(n_300), .Y(n_987) );
OAI211xp5_ASAP7_75t_SL g609 ( .A1(n_301), .A2(n_610), .B(n_613), .C(n_615), .Y(n_609) );
INVx1_ASAP7_75t_L g638 ( .A(n_301), .Y(n_638) );
INVx1_ASAP7_75t_L g652 ( .A(n_302), .Y(n_652) );
INVx1_ASAP7_75t_L g1319 ( .A(n_303), .Y(n_1319) );
CKINVDCx5p33_ASAP7_75t_R g1619 ( .A(n_304), .Y(n_1619) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_305), .Y(n_1192) );
INVx1_ASAP7_75t_L g866 ( .A(n_306), .Y(n_866) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
INVx1_ASAP7_75t_L g1351 ( .A(n_308), .Y(n_1351) );
INVx1_ASAP7_75t_L g1140 ( .A(n_309), .Y(n_1140) );
CKINVDCx5p33_ASAP7_75t_R g1195 ( .A(n_310), .Y(n_1195) );
INVx1_ASAP7_75t_L g709 ( .A(n_311), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_312), .Y(n_806) );
XNOR2xp5_ASAP7_75t_L g1648 ( .A(n_315), .B(n_1649), .Y(n_1648) );
CKINVDCx5p33_ASAP7_75t_R g1629 ( .A(n_316), .Y(n_1629) );
CKINVDCx5p33_ASAP7_75t_R g1223 ( .A(n_317), .Y(n_1223) );
INVx1_ASAP7_75t_L g1374 ( .A(n_318), .Y(n_1374) );
XOR2x2_ASAP7_75t_L g1169 ( .A(n_319), .B(n_1170), .Y(n_1169) );
INVx2_ASAP7_75t_L g439 ( .A(n_321), .Y(n_439) );
INVx1_ASAP7_75t_L g491 ( .A(n_321), .Y(n_491) );
INVx1_ASAP7_75t_L g513 ( .A(n_321), .Y(n_513) );
INVx1_ASAP7_75t_L g742 ( .A(n_322), .Y(n_742) );
INVx1_ASAP7_75t_L g926 ( .A(n_323), .Y(n_926) );
INVx1_ASAP7_75t_L g904 ( .A(n_324), .Y(n_904) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_325), .A2(n_425), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g497 ( .A(n_325), .Y(n_497) );
INVx1_ASAP7_75t_L g895 ( .A(n_326), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_327), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_328), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_356), .B(n_1385), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx4f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_341), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g1642 ( .A(n_335), .B(n_344), .Y(n_1642) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g1646 ( .A(n_337), .B(n_340), .Y(n_1646) );
INVx1_ASAP7_75t_L g1653 ( .A(n_337), .Y(n_1653) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g1656 ( .A(n_340), .B(n_1653), .Y(n_1656) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI21xp5_ASAP7_75t_SL g365 ( .A1(n_344), .A2(n_366), .B(n_400), .Y(n_365) );
AND2x4_ASAP7_75t_L g601 ( .A(n_344), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g420 ( .A(n_345), .B(n_355), .Y(n_420) );
AND2x4_ASAP7_75t_L g428 ( .A(n_345), .B(n_354), .Y(n_428) );
AND2x4_ASAP7_75t_SL g1641 ( .A(n_346), .B(n_1642), .Y(n_1641) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
BUFx4f_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
OR2x6_ASAP7_75t_L g622 ( .A(n_348), .B(n_369), .Y(n_622) );
OR2x2_ASAP7_75t_L g850 ( .A(n_348), .B(n_369), .Y(n_850) );
INVx1_ASAP7_75t_L g1295 ( .A(n_348), .Y(n_1295) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx3_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
BUFx4f_ASAP7_75t_L g674 ( .A(n_349), .Y(n_674) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g371 ( .A(n_351), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_352), .Y(n_378) );
INVx1_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
INVx2_ASAP7_75t_L g398 ( .A(n_351), .Y(n_398) );
NAND2x1_ASAP7_75t_L g412 ( .A(n_351), .B(n_352), .Y(n_412) );
INVx2_ASAP7_75t_L g418 ( .A(n_351), .Y(n_418) );
INVx2_ASAP7_75t_L g372 ( .A(n_352), .Y(n_372) );
BUFx2_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_352), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g417 ( .A(n_352), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g433 ( .A(n_352), .Y(n_433) );
AND2x2_ASAP7_75t_L g435 ( .A(n_352), .B(n_398), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_353), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_384) );
OR2x6_ASAP7_75t_L g599 ( .A(n_353), .B(n_388), .Y(n_599) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
AND2x4_ASAP7_75t_L g390 ( .A(n_355), .B(n_391), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_1211), .B2(n_1212), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
XNOR2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_760), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_604), .B2(n_759), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
XOR2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_524), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_436), .B(n_440), .Y(n_364) );
INVx3_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g600 ( .A(n_368), .Y(n_600) );
CKINVDCx16_ASAP7_75t_R g626 ( .A(n_368), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_368), .A2(n_1005), .B1(n_1006), .B2(n_1007), .Y(n_1004) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_371), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_376), .C(n_379), .Y(n_373) );
INVx1_ASAP7_75t_L g386 ( .A(n_374), .Y(n_386) );
OR2x2_ASAP7_75t_L g395 ( .A(n_374), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g588 ( .A(n_374), .B(n_383), .Y(n_588) );
AND2x2_ASAP7_75t_L g593 ( .A(n_374), .B(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g617 ( .A(n_374), .B(n_383), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_376), .A2(n_575), .B1(n_576), .B2(n_588), .C1(n_589), .C2(n_590), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_376), .B(n_1374), .Y(n_1373) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g614 ( .A(n_377), .B(n_382), .Y(n_614) );
BUFx3_ASAP7_75t_L g1025 ( .A(n_377), .Y(n_1025) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g586 ( .A(n_378), .Y(n_586) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_381), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_381), .A2(n_590), .B1(n_846), .B2(n_847), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_381), .A2(n_390), .B1(n_995), .B2(n_999), .Y(n_1011) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g584 ( .A(n_382), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g597 ( .A(n_382), .B(n_396), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_385), .A2(n_475), .B1(n_477), .B2(n_478), .Y(n_474) );
BUFx3_ASAP7_75t_L g554 ( .A(n_388), .Y(n_554) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_388), .Y(n_564) );
BUFx3_ASAP7_75t_L g651 ( .A(n_388), .Y(n_651) );
INVx2_ASAP7_75t_SL g1329 ( .A(n_388), .Y(n_1329) );
INVx2_ASAP7_75t_L g807 ( .A(n_389), .Y(n_807) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g590 ( .A(n_390), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_390), .A2(n_617), .B1(n_742), .B2(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g915 ( .A(n_390), .Y(n_915) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_399), .Y(n_393) );
INVx2_ASAP7_75t_L g1631 ( .A(n_394), .Y(n_1631) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g624 ( .A(n_395), .Y(n_624) );
INVx2_ASAP7_75t_L g757 ( .A(n_395), .Y(n_757) );
INVx8_ASAP7_75t_L g407 ( .A(n_396), .Y(n_407) );
BUFx2_ASAP7_75t_L g884 ( .A(n_396), .Y(n_884) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_408), .B(n_421), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g883 ( .A1(n_403), .A2(n_866), .B1(n_877), .B2(n_884), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_403), .A2(n_826), .B1(n_871), .B2(n_875), .Y(n_887) );
OAI22xp33_ASAP7_75t_L g1149 ( .A1(n_403), .A2(n_405), .B1(n_1130), .B2(n_1146), .Y(n_1149) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_404), .A2(n_422), .B1(n_516), .B2(n_518), .C(n_521), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_405), .A2(n_725), .B1(n_1136), .B2(n_1141), .Y(n_1152) );
OAI22xp33_ASAP7_75t_L g1318 ( .A1(n_405), .A2(n_927), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_405), .A2(n_1328), .B1(n_1330), .B2(n_1331), .Y(n_1327) );
INVx5_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx6_ASAP7_75t_L g653 ( .A(n_406), .Y(n_653) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx4_ASAP7_75t_L g555 ( .A(n_407), .Y(n_555) );
INVx2_ASAP7_75t_L g566 ( .A(n_407), .Y(n_566) );
INVx1_ASAP7_75t_L g677 ( .A(n_407), .Y(n_677) );
INVx1_ASAP7_75t_L g726 ( .A(n_407), .Y(n_726) );
INVx2_ASAP7_75t_SL g826 ( .A(n_407), .Y(n_826) );
INVx2_ASAP7_75t_L g938 ( .A(n_407), .Y(n_938) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B1(n_414), .B2(n_419), .C(n_420), .Y(n_408) );
OAI22xp5_ASAP7_75t_SL g885 ( .A1(n_409), .A2(n_799), .B1(n_870), .B2(n_874), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_409), .A2(n_414), .B1(n_867), .B2(n_878), .Y(n_886) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g797 ( .A(n_410), .Y(n_797) );
INVx1_ASAP7_75t_L g804 ( .A(n_410), .Y(n_804) );
INVx2_ASAP7_75t_L g955 ( .A(n_410), .Y(n_955) );
INVx4_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx4f_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_411), .Y(n_558) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_411), .Y(n_562) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_411), .Y(n_612) );
BUFx4f_ASAP7_75t_L g729 ( .A(n_411), .Y(n_729) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g660 ( .A(n_412), .Y(n_660) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g656 ( .A(n_416), .Y(n_656) );
INVx2_ASAP7_75t_L g796 ( .A(n_416), .Y(n_796) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g557 ( .A(n_417), .Y(n_557) );
INVx1_ASAP7_75t_L g561 ( .A(n_417), .Y(n_561) );
BUFx2_ASAP7_75t_L g664 ( .A(n_417), .Y(n_664) );
BUFx2_ASAP7_75t_L g799 ( .A(n_417), .Y(n_799) );
AND2x2_ASAP7_75t_L g432 ( .A(n_418), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_420), .B(n_489), .Y(n_568) );
AND2x4_ASAP7_75t_L g668 ( .A(n_420), .B(n_669), .Y(n_668) );
OAI211xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_423), .B(n_424), .C(n_429), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_423), .A2(n_728), .B1(n_1132), .B2(n_1147), .Y(n_1151) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g1023 ( .A(n_431), .Y(n_1023) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_432), .Y(n_594) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g1031 ( .A(n_435), .Y(n_1031) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x6_ASAP7_75t_L g547 ( .A(n_438), .B(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g551 ( .A(n_438), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g791 ( .A(n_438), .B(n_548), .Y(n_791) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g982 ( .A(n_439), .Y(n_982) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_483), .B(n_492), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_474), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_461), .C(n_471), .Y(n_442) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_444), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_528) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g633 ( .A(n_445), .Y(n_633) );
INVx1_ASAP7_75t_L g719 ( .A(n_445), .Y(n_719) );
INVx1_ASAP7_75t_L g945 ( .A(n_445), .Y(n_945) );
INVx1_ASAP7_75t_L g965 ( .A(n_445), .Y(n_965) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_446), .Y(n_545) );
INVx3_ASAP7_75t_L g775 ( .A(n_446), .Y(n_775) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g684 ( .A(n_447), .Y(n_684) );
BUFx2_ASAP7_75t_L g739 ( .A(n_447), .Y(n_739) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
BUFx2_ASAP7_75t_L g460 ( .A(n_448), .Y(n_460) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_449), .B(n_451), .Y(n_470) );
INVx2_ASAP7_75t_L g473 ( .A(n_449), .Y(n_473) );
BUFx2_ASAP7_75t_L g457 ( .A(n_450), .Y(n_457) );
AND2x4_ASAP7_75t_L g507 ( .A(n_450), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g1252 ( .A(n_450), .Y(n_1252) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g465 ( .A(n_451), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g472 ( .A(n_451), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g482 ( .A(n_451), .Y(n_482) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g572 ( .A1(n_453), .A2(n_459), .B1(n_573), .B2(n_574), .C1(n_575), .C2(n_576), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_453), .A2(n_459), .B1(n_806), .B2(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_453), .A2(n_459), .B1(n_846), .B2(n_855), .Y(n_854) );
AOI222xp33_ASAP7_75t_L g892 ( .A1(n_453), .A2(n_640), .B1(n_893), .B2(n_894), .C1(n_895), .C2(n_896), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_453), .A2(n_459), .B1(n_999), .B2(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_453), .A2(n_459), .B1(n_1041), .B2(n_1050), .Y(n_1049) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_453), .A2(n_1241), .B1(n_1250), .B2(n_1253), .Y(n_1249) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_457), .Y(n_453) );
AND2x2_ASAP7_75t_L g459 ( .A(n_454), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g637 ( .A(n_454), .B(n_457), .Y(n_637) );
AND2x4_ASAP7_75t_L g640 ( .A(n_454), .B(n_460), .Y(n_640) );
AND2x4_ASAP7_75t_L g967 ( .A(n_454), .B(n_457), .Y(n_967) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND3x4_ASAP7_75t_L g981 ( .A(n_455), .B(n_486), .C(n_982), .Y(n_981) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_455), .B(n_1254), .Y(n_1253) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g464 ( .A(n_456), .Y(n_464) );
NAND2xp33_ASAP7_75t_SL g495 ( .A(n_456), .B(n_486), .Y(n_495) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_459), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_459), .A2(n_967), .B1(n_1261), .B2(n_1270), .Y(n_1269) );
AOI32xp33_ASAP7_75t_L g1637 ( .A1(n_459), .A2(n_1251), .A3(n_1253), .B1(n_1629), .B2(n_1638), .Y(n_1637) );
BUFx2_ASAP7_75t_L g630 ( .A(n_462), .Y(n_630) );
BUFx3_ASAP7_75t_L g745 ( .A(n_462), .Y(n_745) );
INVx2_ASAP7_75t_SL g905 ( .A(n_462), .Y(n_905) );
OR2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
AND2x2_ASAP7_75t_L g478 ( .A(n_463), .B(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g645 ( .A(n_463), .B(n_479), .Y(n_645) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x6_ASAP7_75t_L g468 ( .A(n_464), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g471 ( .A(n_464), .B(n_472), .Y(n_471) );
OR2x4_ASAP7_75t_L g476 ( .A(n_464), .B(n_465), .Y(n_476) );
NAND3x1_ASAP7_75t_L g511 ( .A(n_464), .B(n_512), .C(n_514), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_464), .B(n_514), .Y(n_548) );
BUFx4f_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
BUFx3_ASAP7_75t_L g682 ( .A(n_465), .Y(n_682) );
BUFx3_ASAP7_75t_L g694 ( .A(n_465), .Y(n_694) );
INVx2_ASAP7_75t_L g788 ( .A(n_465), .Y(n_788) );
INVx1_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g481 ( .A(n_467), .Y(n_481) );
INVx2_ASAP7_75t_L g579 ( .A(n_468), .Y(n_579) );
INVx1_ASAP7_75t_L g747 ( .A(n_468), .Y(n_747) );
INVx1_ASAP7_75t_L g900 ( .A(n_468), .Y(n_900) );
BUFx3_ASAP7_75t_L g970 ( .A(n_468), .Y(n_970) );
BUFx3_ASAP7_75t_L g688 ( .A(n_469), .Y(n_688) );
INVx1_ASAP7_75t_L g712 ( .A(n_469), .Y(n_712) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g520 ( .A(n_470), .Y(n_520) );
CKINVDCx8_ASAP7_75t_R g634 ( .A(n_471), .Y(n_634) );
CKINVDCx8_ASAP7_75t_R g816 ( .A(n_471), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_471), .B(n_891), .Y(n_890) );
BUFx2_ASAP7_75t_L g504 ( .A(n_472), .Y(n_504) );
BUFx2_ASAP7_75t_L g573 ( .A(n_472), .Y(n_573) );
BUFx2_ASAP7_75t_L g896 ( .A(n_472), .Y(n_896) );
BUFx3_ASAP7_75t_L g986 ( .A(n_472), .Y(n_986) );
INVx2_ASAP7_75t_L g997 ( .A(n_472), .Y(n_997) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_472), .Y(n_1048) );
INVx1_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
INVx1_ASAP7_75t_L g1187 ( .A(n_475), .Y(n_1187) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g643 ( .A(n_476), .Y(n_643) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_476), .Y(n_734) );
INVx1_ASAP7_75t_L g903 ( .A(n_476), .Y(n_903) );
INVx2_ASAP7_75t_L g571 ( .A(n_478), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_478), .A2(n_898), .B1(n_899), .B2(n_900), .Y(n_897) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_479), .Y(n_499) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_479), .Y(n_687) );
INVx2_ASAP7_75t_L g690 ( .A(n_479), .Y(n_690) );
INVx1_ASAP7_75t_L g715 ( .A(n_479), .Y(n_715) );
INVx2_ASAP7_75t_L g949 ( .A(n_479), .Y(n_949) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
BUFx8_ASAP7_75t_L g539 ( .A(n_480), .Y(n_539) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_480), .Y(n_708) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x4_ASAP7_75t_L g502 ( .A(n_482), .B(n_503), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g628 ( .A1(n_483), .A2(n_629), .A3(n_632), .B(n_641), .Y(n_628) );
BUFx2_ASAP7_75t_L g1122 ( .A(n_483), .Y(n_1122) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_484), .B(n_487), .Y(n_483) );
AND2x2_ASAP7_75t_L g580 ( .A(n_484), .B(n_487), .Y(n_580) );
AND2x2_ASAP7_75t_L g748 ( .A(n_484), .B(n_487), .Y(n_748) );
AND2x4_ASAP7_75t_L g907 ( .A(n_484), .B(n_487), .Y(n_907) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_484), .B(n_487), .Y(n_1002) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g494 ( .A(n_489), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g670 ( .A(n_489), .Y(n_670) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g603 ( .A(n_490), .Y(n_603) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_496), .B1(n_509), .B2(n_515), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g527 ( .A1(n_493), .A2(n_528), .A3(n_532), .B1(n_537), .B2(n_543), .B3(n_547), .Y(n_527) );
OAI33xp33_ASAP7_75t_L g863 ( .A1(n_493), .A2(n_547), .A3(n_864), .B1(n_868), .B2(n_872), .B3(n_876), .Y(n_863) );
OAI33xp33_ASAP7_75t_L g1332 ( .A1(n_493), .A2(n_950), .A3(n_1333), .B1(n_1336), .B2(n_1337), .B3(n_1338), .Y(n_1332) );
OAI33xp33_ASAP7_75t_L g1360 ( .A1(n_493), .A2(n_547), .A3(n_1361), .B1(n_1362), .B2(n_1363), .B3(n_1366), .Y(n_1360) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx8_ASAP7_75t_L g680 ( .A(n_494), .Y(n_680) );
BUFx4f_ASAP7_75t_L g770 ( .A(n_494), .Y(n_770) );
BUFx4f_ASAP7_75t_L g1096 ( .A(n_494), .Y(n_1096) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_500), .C(n_505), .Y(n_496) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_498), .A2(n_518), .B1(n_1322), .B2(n_1330), .Y(n_1336) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g988 ( .A(n_501), .Y(n_988) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx8_ASAP7_75t_L g523 ( .A(n_502), .Y(n_523) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx5_ASAP7_75t_L g979 ( .A(n_507), .Y(n_979) );
INVx1_ASAP7_75t_L g1254 ( .A(n_508), .Y(n_1254) );
OAI33xp33_ASAP7_75t_L g679 ( .A1(n_509), .A2(n_680), .A3(n_681), .B1(n_685), .B2(n_689), .B3(n_691), .Y(n_679) );
OAI33xp33_ASAP7_75t_L g699 ( .A1(n_509), .A2(n_680), .A3(n_700), .B1(n_704), .B2(n_713), .B3(n_717), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g950 ( .A(n_510), .Y(n_950) );
INVx2_ASAP7_75t_L g1104 ( .A(n_510), .Y(n_1104) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g1144 ( .A(n_511), .Y(n_1144) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_516), .A2(n_533), .B1(n_534), .B2(n_535), .Y(n_532) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g783 ( .A(n_517), .Y(n_783) );
BUFx2_ASAP7_75t_L g869 ( .A(n_517), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_518), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
OAI22xp33_ASAP7_75t_SL g948 ( .A1(n_518), .A2(n_932), .B1(n_939), .B2(n_949), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_518), .A2(n_707), .B1(n_1086), .B2(n_1093), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_518), .A2(n_1138), .B1(n_1140), .B2(n_1141), .Y(n_1137) );
CKINVDCx8_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g541 ( .A(n_519), .Y(n_541) );
INVx3_ASAP7_75t_L g779 ( .A(n_519), .Y(n_779) );
INVx3_ASAP7_75t_L g1071 ( .A(n_519), .Y(n_1071) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g536 ( .A(n_520), .Y(n_536) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_569), .C(n_581), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_549), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_529), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_529), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g1072 ( .A1(n_529), .A2(n_719), .B1(n_1056), .B2(n_1062), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_529), .A2(n_774), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_529), .A2(n_684), .B1(n_1229), .B2(n_1230), .Y(n_1228) );
OAI22xp33_ASAP7_75t_L g1276 ( .A1(n_529), .A2(n_545), .B1(n_1277), .B2(n_1278), .Y(n_1276) );
OAI22xp33_ASAP7_75t_L g1286 ( .A1(n_529), .A2(n_684), .B1(n_1287), .B2(n_1288), .Y(n_1286) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_529), .A2(n_774), .B1(n_1350), .B2(n_1358), .Y(n_1361) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_529), .A2(n_684), .B1(n_1351), .B2(n_1359), .Y(n_1366) );
OAI22xp33_ASAP7_75t_L g1608 ( .A1(n_529), .A2(n_545), .B1(n_1609), .B2(n_1610), .Y(n_1608) );
OAI22xp33_ASAP7_75t_L g1617 ( .A1(n_529), .A2(n_684), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_530), .A2(n_544), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_531), .A2(n_546), .B1(n_560), .B2(n_562), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_533), .A2(n_540), .B1(n_557), .B2(n_558), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_534), .A2(n_542), .B1(n_564), .B2(n_565), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_535), .A2(n_869), .B1(n_870), .B2(n_871), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_535), .A2(n_873), .B1(n_874), .B2(n_875), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g1282 ( .A1(n_535), .A2(n_1283), .B1(n_1284), .B2(n_1285), .Y(n_1282) );
OAI22xp5_ASAP7_75t_L g1614 ( .A1(n_535), .A2(n_1069), .B1(n_1615), .B2(n_1616), .Y(n_1614) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g1365 ( .A(n_536), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_538), .A2(n_785), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_538), .A2(n_1348), .B1(n_1356), .B2(n_1364), .Y(n_1363) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g873 ( .A(n_539), .Y(n_873) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_539), .Y(n_1283) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_541), .A2(n_830), .B1(n_836), .B2(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_545), .A2(n_787), .B1(n_825), .B2(n_832), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_545), .A2(n_682), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g1183 ( .A(n_545), .Y(n_1183) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_545), .A2(n_943), .B1(n_1320), .B2(n_1326), .Y(n_1338) );
INVx1_ASAP7_75t_L g990 ( .A(n_547), .Y(n_990) );
OAI33xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_553), .A3(n_556), .B1(n_559), .B2(n_563), .B3(n_567), .Y(n_549) );
OAI33xp33_ASAP7_75t_L g792 ( .A1(n_550), .A2(n_793), .A3(n_795), .B1(n_798), .B2(n_800), .B3(n_801), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g1289 ( .A1(n_550), .A2(n_567), .A3(n_1290), .B1(n_1291), .B2(n_1292), .B3(n_1293), .Y(n_1289) );
OAI33xp33_ASAP7_75t_L g1620 ( .A1(n_550), .A2(n_567), .A3(n_1621), .B1(n_1622), .B2(n_1623), .B3(n_1624), .Y(n_1620) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g648 ( .A(n_551), .Y(n_648) );
INVx2_ASAP7_75t_L g723 ( .A(n_551), .Y(n_723) );
INVx2_ASAP7_75t_L g1080 ( .A(n_551), .Y(n_1080) );
INVx1_ASAP7_75t_L g1193 ( .A(n_551), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_554), .A2(n_565), .B1(n_1220), .B2(n_1229), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_554), .A2(n_555), .B1(n_1224), .B2(n_1227), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_554), .A2(n_565), .B1(n_1355), .B2(n_1356), .Y(n_1354) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_555), .A2(n_778), .B1(n_784), .B2(n_794), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g1293 ( .A1(n_555), .A2(n_1281), .B1(n_1285), .B2(n_1294), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1621 ( .A1(n_555), .A2(n_794), .B1(n_1609), .B2(n_1618), .Y(n_1621) );
OAI22xp5_ASAP7_75t_L g1624 ( .A1(n_555), .A2(n_1294), .B1(n_1613), .B2(n_1616), .Y(n_1624) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_557), .A2(n_955), .B1(n_1221), .B2(n_1230), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_557), .A2(n_729), .B1(n_1358), .B2(n_1359), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_560), .A2(n_658), .B1(n_934), .B2(n_935), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_560), .A2(n_804), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_560), .A2(n_612), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1321 ( .A1(n_560), .A2(n_658), .B1(n_1322), .B2(n_1323), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_560), .A2(n_612), .B1(n_1325), .B2(n_1326), .Y(n_1324) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g1234 ( .A(n_561), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_562), .A2(n_796), .B1(n_832), .B2(n_833), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_562), .A2(n_796), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_562), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_562), .A2(n_1234), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_565), .A2(n_772), .B1(n_789), .B2(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_565), .A2(n_794), .B1(n_835), .B2(n_836), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_565), .A2(n_794), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI33xp33_ASAP7_75t_L g1231 ( .A1(n_567), .A2(n_723), .A3(n_1232), .B1(n_1233), .B2(n_1235), .B3(n_1236), .Y(n_1231) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g801 ( .A(n_568), .Y(n_801) );
AOI33xp33_ASAP7_75t_L g1021 ( .A1(n_568), .A2(n_882), .A3(n_1022), .B1(n_1024), .B2(n_1026), .B3(n_1027), .Y(n_1021) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_577), .B(n_580), .Y(n_569) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g631 ( .A(n_579), .Y(n_631) );
OAI31xp33_ASAP7_75t_SL g811 ( .A1(n_580), .A2(n_812), .A3(n_813), .B(n_819), .Y(n_811) );
OAI31xp33_ASAP7_75t_SL g851 ( .A1(n_580), .A2(n_852), .A3(n_853), .B(n_856), .Y(n_851) );
OAI31xp33_ASAP7_75t_SL g1244 ( .A1(n_580), .A2(n_1245), .A3(n_1246), .B(n_1247), .Y(n_1244) );
OAI31xp33_ASAP7_75t_L g1265 ( .A1(n_580), .A2(n_1266), .A3(n_1268), .B(n_1273), .Y(n_1265) );
OAI31xp33_ASAP7_75t_SL g1633 ( .A1(n_580), .A2(n_1634), .A3(n_1635), .B(n_1639), .Y(n_1633) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_598), .B(n_601), .Y(n_581) );
NAND3xp33_ASAP7_75t_SL g582 ( .A(n_583), .B(n_587), .C(n_591), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g1015 ( .A(n_584), .Y(n_1015) );
INVx1_ASAP7_75t_L g1014 ( .A(n_585), .Y(n_1014) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_588), .A2(n_1174), .B1(n_1175), .B2(n_1176), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_588), .A2(n_1175), .B1(n_1306), .B2(n_1313), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_588), .A2(n_590), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
AOI22xp5_ASAP7_75t_L g1627 ( .A1(n_588), .A2(n_807), .B1(n_1628), .B2(n_1629), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_590), .A2(n_616), .B1(n_618), .B2(n_619), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_590), .A2(n_617), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1240 ( .A1(n_590), .A2(n_617), .B1(n_1241), .B2(n_1242), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_590), .A2(n_617), .B1(n_1261), .B2(n_1262), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_591) );
INVx3_ASAP7_75t_L g1029 ( .A(n_594), .Y(n_1029) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g1006 ( .A(n_599), .Y(n_1006) );
BUFx2_ASAP7_75t_L g627 ( .A(n_601), .Y(n_627) );
BUFx2_ASAP7_75t_SL g758 ( .A(n_601), .Y(n_758) );
INVx1_ASAP7_75t_L g1016 ( .A(n_601), .Y(n_1016) );
OAI31xp33_ASAP7_75t_L g1037 ( .A1(n_601), .A2(n_1038), .A3(n_1039), .B(n_1043), .Y(n_1037) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_601), .Y(n_1114) );
OAI31xp33_ASAP7_75t_L g1237 ( .A1(n_601), .A2(n_1238), .A3(n_1239), .B(n_1243), .Y(n_1237) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g759 ( .A(n_604), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_695), .B2(n_696), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_628), .C(n_646), .Y(n_607) );
OAI31xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_620), .A3(n_625), .B(n_627), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_612), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_613), .B(n_1370), .C(n_1373), .Y(n_1369) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g752 ( .A(n_614), .Y(n_752) );
INVx1_ASAP7_75t_L g1112 ( .A(n_614), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_616), .A2(n_914), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
BUFx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_617), .A2(n_893), .B1(n_895), .B2(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_617), .A2(n_807), .B1(n_957), .B2(n_958), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_617), .A2(n_807), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_618), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_635) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_622), .Y(n_1160) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI31xp33_ASAP7_75t_L g802 ( .A1(n_627), .A2(n_803), .A3(n_809), .B(n_810), .Y(n_802) );
OAI31xp33_ASAP7_75t_L g843 ( .A1(n_627), .A2(n_844), .A3(n_848), .B(n_849), .Y(n_843) );
INVx1_ASAP7_75t_L g918 ( .A(n_627), .Y(n_918) );
OAI31xp33_ASAP7_75t_L g953 ( .A1(n_627), .A2(n_954), .A3(n_959), .B(n_961), .Y(n_953) );
OAI31xp33_ASAP7_75t_L g1367 ( .A1(n_627), .A2(n_1368), .A3(n_1369), .B(n_1375), .Y(n_1367) );
OAI31xp33_ASAP7_75t_L g1625 ( .A1(n_627), .A2(n_1626), .A3(n_1630), .B(n_1632), .Y(n_1625) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_633), .A2(n_652), .B1(n_666), .B2(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g1145 ( .A1(n_633), .A2(n_1131), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1208 ( .A1(n_633), .A2(n_692), .B1(n_1192), .B2(n_1199), .Y(n_1208) );
NAND3xp33_ASAP7_75t_L g1379 ( .A(n_634), .B(n_1380), .C(n_1381), .Y(n_1379) );
BUFx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx3_ASAP7_75t_L g741 ( .A(n_637), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_639), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_639), .A2(n_741), .B1(n_1110), .B2(n_1119), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_640), .A2(n_957), .B1(n_967), .B2(n_968), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g1166 ( .A1(n_640), .A2(n_967), .B1(n_1157), .B2(n_1167), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_640), .A2(n_967), .B1(n_1174), .B2(n_1185), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_640), .A2(n_967), .B1(n_1306), .B2(n_1307), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_640), .A2(n_967), .B1(n_1371), .B2(n_1374), .Y(n_1380) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g735 ( .A(n_645), .Y(n_735) );
INVx1_ASAP7_75t_L g1267 ( .A(n_645), .Y(n_1267) );
INVx1_ASAP7_75t_L g1309 ( .A(n_645), .Y(n_1309) );
NOR2xp33_ASAP7_75t_SL g646 ( .A(n_647), .B(n_679), .Y(n_646) );
OAI33xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .A3(n_654), .B1(n_661), .B2(n_667), .B3(n_671), .Y(n_647) );
INVx2_ASAP7_75t_SL g882 ( .A(n_648), .Y(n_882) );
OAI33xp33_ASAP7_75t_L g924 ( .A1(n_648), .A2(n_925), .A3(n_929), .B1(n_933), .B2(n_936), .B3(n_940), .Y(n_924) );
INVx2_ASAP7_75t_SL g1353 ( .A(n_648), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_652), .B2(n_653), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_650), .A2(n_665), .B1(n_682), .B2(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_651), .A2(n_653), .B1(n_709), .B2(n_716), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_651), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_651), .A2(n_653), .B1(n_1093), .B2(n_1094), .Y(n_1092) );
OAI22xp5_ASAP7_75t_SL g1081 ( .A1(n_653), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_653), .A2(n_927), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1200 ( .A1(n_653), .A2(n_927), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_655), .A2(n_675), .B1(n_686), .B2(n_688), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_656), .A2(n_660), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_657), .A2(n_678), .B1(n_688), .B2(n_690), .Y(n_689) );
INVx5_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_662), .B1(n_665), .B2(n_666), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_660), .A2(n_662), .B1(n_702), .B2(n_720), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_660), .A2(n_773), .B1(n_790), .B2(n_799), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_660), .A2(n_796), .B1(n_829), .B2(n_830), .Y(n_828) );
BUFx2_ASAP7_75t_SL g1090 ( .A(n_660), .Y(n_1090) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_660), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1292 ( .A1(n_660), .A2(n_1234), .B1(n_1278), .B2(n_1288), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_662), .A2(n_1089), .B1(n_1090), .B2(n_1091), .Y(n_1088) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx4_ASAP7_75t_L g728 ( .A(n_663), .Y(n_728) );
INVx2_ASAP7_75t_L g931 ( .A(n_663), .Y(n_931) );
INVx4_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI33xp33_ASAP7_75t_L g721 ( .A1(n_667), .A2(n_722), .A3(n_724), .B1(n_727), .B2(n_730), .B3(n_731), .Y(n_721) );
OAI33xp33_ASAP7_75t_L g1079 ( .A1(n_667), .A2(n_1080), .A3(n_1081), .B1(n_1085), .B2(n_1088), .B3(n_1092), .Y(n_1079) );
OAI33xp33_ASAP7_75t_L g1148 ( .A1(n_667), .A2(n_722), .A3(n_1149), .B1(n_1150), .B2(n_1151), .B3(n_1152), .Y(n_1148) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_668), .Y(n_940) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .B1(n_676), .B2(n_678), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g725 ( .A(n_673), .Y(n_725) );
INVx3_ASAP7_75t_L g927 ( .A(n_673), .Y(n_927) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx4_ASAP7_75t_L g794 ( .A(n_674), .Y(n_794) );
INVx3_ASAP7_75t_L g1083 ( .A(n_674), .Y(n_1083) );
BUFx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g1349 ( .A1(n_677), .A2(n_794), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
OAI33xp33_ASAP7_75t_L g941 ( .A1(n_680), .A2(n_942), .A3(n_946), .B1(n_948), .B2(n_950), .B3(n_951), .Y(n_941) );
OAI33xp33_ASAP7_75t_L g1203 ( .A1(n_680), .A2(n_950), .A3(n_1204), .B1(n_1205), .B2(n_1207), .B3(n_1208), .Y(n_1203) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_682), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_682), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_684), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_684), .A2(n_787), .B1(n_789), .B2(n_790), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_684), .A2(n_787), .B1(n_827), .B2(n_833), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g1067 ( .A1(n_684), .A2(n_787), .B1(n_1055), .B2(n_1061), .Y(n_1067) );
INVx2_ASAP7_75t_L g1101 ( .A(n_684), .Y(n_1101) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g1206 ( .A(n_687), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_688), .A2(n_930), .B1(n_937), .B2(n_947), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_688), .A2(n_841), .B1(n_1087), .B2(n_1094), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1337 ( .A1(n_688), .A2(n_947), .B1(n_1323), .B2(n_1331), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_690), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_690), .A2(n_779), .B1(n_829), .B2(n_835), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_690), .A2(n_1059), .B1(n_1065), .B2(n_1071), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_690), .A2(n_779), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g944 ( .A(n_694), .Y(n_944) );
INVxp67_ASAP7_75t_SL g1099 ( .A(n_694), .Y(n_1099) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_732), .C(n_749), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_721), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_701), .A2(n_718), .B1(n_725), .B2(n_726), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_709), .B2(n_710), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_705), .A2(n_714), .B1(n_728), .B2(n_729), .Y(n_727) );
BUFx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx8_ASAP7_75t_L g1139 ( .A(n_707), .Y(n_1139) );
OAI22xp33_ASAP7_75t_SL g1362 ( .A1(n_707), .A2(n_785), .B1(n_1347), .B2(n_1355), .Y(n_1362) );
INVx5_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g841 ( .A(n_708), .Y(n_841) );
INVx3_ASAP7_75t_L g1069 ( .A(n_708), .Y(n_1069) );
OAI22xp33_ASAP7_75t_SL g1134 ( .A1(n_710), .A2(n_1069), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_710), .A2(n_1195), .B1(n_1201), .B2(n_1206), .Y(n_1205) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_710), .A2(n_949), .B1(n_1196), .B2(n_1202), .Y(n_1207) );
INVx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g785 ( .A(n_712), .Y(n_785) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI33xp33_ASAP7_75t_L g823 ( .A1(n_723), .A2(n_801), .A3(n_824), .B1(n_828), .B2(n_831), .B3(n_834), .Y(n_823) );
OAI33xp33_ASAP7_75t_L g1053 ( .A1(n_723), .A2(n_801), .A3(n_1054), .B1(n_1057), .B2(n_1060), .B3(n_1063), .Y(n_1053) );
OAI22xp33_ASAP7_75t_L g1290 ( .A1(n_726), .A2(n_794), .B1(n_1277), .B2(n_1287), .Y(n_1290) );
OAI22xp33_ASAP7_75t_L g1150 ( .A1(n_728), .A2(n_804), .B1(n_1135), .B2(n_1140), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_729), .A2(n_796), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_729), .A2(n_1223), .B1(n_1226), .B2(n_1234), .Y(n_1233) );
OAI31xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .A3(n_744), .B(n_748), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_SL g1133 ( .A(n_738), .Y(n_1133) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g815 ( .A(n_739), .Y(n_815) );
INVx1_ASAP7_75t_L g1335 ( .A(n_739), .Y(n_1335) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI31xp33_ASAP7_75t_L g962 ( .A1(n_748), .A2(n_963), .A3(n_964), .B(n_969), .Y(n_962) );
OAI31xp33_ASAP7_75t_L g1162 ( .A1(n_748), .A2(n_1163), .A3(n_1165), .B(n_1168), .Y(n_1162) );
OAI31xp33_ASAP7_75t_L g1179 ( .A1(n_748), .A2(n_1180), .A3(n_1181), .B(n_1186), .Y(n_1179) );
OAI31xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .A3(n_755), .B(n_758), .Y(n_749) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g911 ( .A(n_757), .Y(n_911) );
INVxp67_ASAP7_75t_SL g960 ( .A(n_757), .Y(n_960) );
INVx1_ASAP7_75t_L g1376 ( .A(n_757), .Y(n_1376) );
OAI31xp33_ASAP7_75t_L g1171 ( .A1(n_758), .A2(n_1172), .A3(n_1177), .B(n_1178), .Y(n_1171) );
OAI31xp33_ASAP7_75t_SL g1257 ( .A1(n_758), .A2(n_1258), .A3(n_1263), .B(n_1264), .Y(n_1257) );
OAI31xp33_ASAP7_75t_L g1310 ( .A1(n_758), .A2(n_1311), .A3(n_1314), .B(n_1315), .Y(n_1310) );
XNOR2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_1074), .Y(n_760) );
XOR2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_857), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
XNOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_820), .Y(n_764) );
XNOR2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
AND3x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_802), .C(n_811), .Y(n_767) );
NOR2xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_792), .Y(n_768) );
OAI33xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .A3(n_776), .B1(n_780), .B2(n_786), .B3(n_791), .Y(n_769) );
OAI33xp33_ASAP7_75t_L g837 ( .A1(n_770), .A2(n_791), .A3(n_838), .B1(n_839), .B2(n_840), .B3(n_842), .Y(n_837) );
OAI33xp33_ASAP7_75t_L g1066 ( .A1(n_770), .A2(n_791), .A3(n_1067), .B1(n_1068), .B2(n_1070), .B3(n_1072), .Y(n_1066) );
OAI33xp33_ASAP7_75t_L g1218 ( .A1(n_770), .A2(n_791), .A3(n_1219), .B1(n_1222), .B2(n_1225), .B3(n_1228), .Y(n_1218) );
OAI33xp33_ASAP7_75t_L g1275 ( .A1(n_770), .A2(n_791), .A3(n_1276), .B1(n_1279), .B2(n_1282), .B3(n_1286), .Y(n_1275) );
OAI33xp33_ASAP7_75t_L g1607 ( .A1(n_770), .A2(n_791), .A3(n_1608), .B1(n_1611), .B2(n_1614), .B3(n_1617), .Y(n_1607) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_774), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
INVx3_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g952 ( .A(n_775), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_777), .A2(n_781), .B1(n_796), .B2(n_797), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_779), .A2(n_1058), .B1(n_1064), .B2(n_1069), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_784), .B2(n_785), .Y(n_780) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g947 ( .A(n_783), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g1611 ( .A1(n_785), .A2(n_1283), .B1(n_1612), .B2(n_1613), .Y(n_1611) );
INVx2_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g865 ( .A(n_788), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_794), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_794), .A2(n_826), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1291 ( .A1(n_797), .A2(n_1234), .B1(n_1280), .B2(n_1284), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g1622 ( .A1(n_797), .A2(n_1234), .B1(n_1612), .B2(n_1615), .Y(n_1622) );
OAI22xp5_ASAP7_75t_L g1623 ( .A1(n_797), .A2(n_1234), .B1(n_1610), .B2(n_1619), .Y(n_1623) );
OAI33xp33_ASAP7_75t_L g880 ( .A1(n_801), .A2(n_881), .A3(n_883), .B1(n_885), .B2(n_886), .B3(n_887), .Y(n_880) );
OAI33xp33_ASAP7_75t_L g1345 ( .A1(n_801), .A2(n_1346), .A3(n_1349), .B1(n_1352), .B2(n_1354), .B3(n_1357), .Y(n_1345) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_814), .A2(n_1084), .B1(n_1091), .B2(n_1098), .Y(n_1105) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND3xp33_ASAP7_75t_SL g993 ( .A(n_816), .B(n_994), .C(n_998), .Y(n_993) );
NAND3xp33_ASAP7_75t_SL g1046 ( .A(n_816), .B(n_1047), .C(n_1049), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_816), .B(n_1269), .C(n_1271), .Y(n_1268) );
AND3x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_843), .C(n_851), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_837), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_826), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_841), .A2(n_1071), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B1(n_972), .B2(n_1073), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_920), .B1(n_921), .B2(n_971), .Y(n_859) );
INVx1_ASAP7_75t_L g971 ( .A(n_860), .Y(n_971) );
INVxp67_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NOR4xp25_ASAP7_75t_L g919 ( .A(n_863), .B(n_880), .C(n_889), .D(n_908), .Y(n_919) );
BUFx4f_ASAP7_75t_SL g1131 ( .A(n_865), .Y(n_1131) );
INVxp67_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVxp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AOI31xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_897), .A3(n_901), .B(n_906), .Y(n_889) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g1121 ( .A(n_900), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_901) );
INVx1_ASAP7_75t_L g1164 ( .A(n_903), .Y(n_1164) );
CKINVDCx14_ASAP7_75t_R g906 ( .A(n_907), .Y(n_906) );
OAI31xp33_ASAP7_75t_L g1302 ( .A1(n_907), .A2(n_1303), .A3(n_1304), .B(n_1308), .Y(n_1302) );
AOI31xp67_ASAP7_75t_SL g908 ( .A1(n_909), .A2(n_912), .A3(n_916), .B(n_918), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g1175 ( .A(n_915), .Y(n_1175) );
INVxp67_ASAP7_75t_SL g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_953), .C(n_962), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_941), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_926), .A2(n_934), .B1(n_943), .B2(n_945), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g951 ( .A1(n_928), .A2(n_935), .B1(n_943), .B2(n_952), .Y(n_951) );
OAI33xp33_ASAP7_75t_L g1189 ( .A1(n_940), .A2(n_1190), .A3(n_1193), .B1(n_1194), .B2(n_1197), .B3(n_1200), .Y(n_1189) );
OAI33xp33_ASAP7_75t_L g1317 ( .A1(n_940), .A2(n_1080), .A3(n_1318), .B1(n_1321), .B2(n_1324), .B3(n_1327), .Y(n_1317) );
OAI22xp33_ASAP7_75t_L g1204 ( .A1(n_943), .A2(n_952), .B1(n_1191), .B2(n_1198), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_943), .A2(n_1319), .B1(n_1325), .B2(n_1334), .Y(n_1333) );
INVx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g1636 ( .A(n_967), .Y(n_1636) );
INVx2_ASAP7_75t_L g1073 ( .A(n_972), .Y(n_1073) );
XNOR2x1_ASAP7_75t_L g972 ( .A(n_973), .B(n_1035), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_974), .B(n_1017), .Y(n_973) );
INVx1_ASAP7_75t_L g1019 ( .A(n_975), .Y(n_1019) );
AOI21xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .B(n_983), .Y(n_975) );
INVx2_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
OAI221xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_987), .B1(n_988), .B2(n_989), .C(n_990), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_986), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_991), .B(n_1003), .Y(n_1018) );
OAI31xp33_ASAP7_75t_SL g991 ( .A1(n_992), .A2(n_993), .A3(n_1001), .B(n_1002), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1000), .B(n_1013), .Y(n_1012) );
OAI31xp33_ASAP7_75t_SL g1044 ( .A1(n_1002), .A2(n_1045), .A3(n_1046), .B(n_1051), .Y(n_1044) );
OAI31xp33_ASAP7_75t_L g1377 ( .A1(n_1002), .A2(n_1378), .A3(n_1379), .B(n_1382), .Y(n_1377) );
AO21x1_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1008), .B(n_1016), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
NAND3xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .C(n_1015), .Y(n_1010) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
OAI31xp33_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1019), .A3(n_1020), .B(n_1032), .Y(n_1017) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1021), .Y(n_1034) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1034), .Y(n_1032) );
NAND3xp33_ASAP7_75t_SL g1036 ( .A(n_1037), .B(n_1044), .C(n_1052), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1042), .B(n_1048), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1048), .B(n_1372), .Y(n_1381) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1066), .Y(n_1052) );
XNOR2xp5_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1123), .Y(n_1074) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1076), .Y(n_1075) );
NAND3xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1106), .C(n_1115), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1095), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_1082), .A2(n_1089), .B1(n_1098), .B2(n_1100), .Y(n_1097) );
OAI33xp33_ASAP7_75t_L g1095 ( .A1(n_1096), .A2(n_1097), .A3(n_1102), .B1(n_1103), .B2(n_1104), .B3(n_1105), .Y(n_1095) );
OAI33xp33_ASAP7_75t_L g1128 ( .A1(n_1096), .A2(n_1129), .A3(n_1134), .B1(n_1137), .B2(n_1142), .B3(n_1145), .Y(n_1128) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
OAI31xp33_ASAP7_75t_L g1106 ( .A1(n_1107), .A2(n_1108), .A3(n_1113), .B(n_1114), .Y(n_1106) );
OAI31xp33_ASAP7_75t_SL g1153 ( .A1(n_1114), .A2(n_1154), .A3(n_1159), .B(n_1161), .Y(n_1153) );
OAI31xp33_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1117), .A3(n_1120), .B(n_1122), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1169), .B1(n_1209), .B2(n_1210), .Y(n_1123) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1124), .Y(n_1209) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1153), .C(n_1162), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1148), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_1130), .A2(n_1131), .B1(n_1132), .B2(n_1133), .Y(n_1129) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1169), .Y(n_1210) );
NAND3xp33_ASAP7_75t_SL g1170 ( .A(n_1171), .B(n_1179), .C(n_1188), .Y(n_1170) );
INVx2_ASAP7_75t_SL g1182 ( .A(n_1183), .Y(n_1182) );
NOR2xp33_ASAP7_75t_SL g1188 ( .A(n_1189), .B(n_1203), .Y(n_1188) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
XNOR2xp5_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1298), .Y(n_1212) );
AOI22xp5_ASAP7_75t_L g1213 ( .A1(n_1214), .A2(n_1255), .B1(n_1296), .B2(n_1297), .Y(n_1213) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1214), .Y(n_1296) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
NAND3xp33_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1237), .C(n_1244), .Y(n_1216) );
NOR2xp33_ASAP7_75t_SL g1217 ( .A(n_1218), .B(n_1231), .Y(n_1217) );
INVx3_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx2_ASAP7_75t_SL g1297 ( .A(n_1255), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1265), .C(n_1274), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1262), .B(n_1272), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1289), .Y(n_1274) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1341), .B2(n_1342), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1301), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1310), .C(n_1316), .Y(n_1301) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1332), .Y(n_1316) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx3_ASAP7_75t_SL g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1343), .Y(n_1384) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1367), .C(n_1377), .Y(n_1343) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1360), .Y(n_1344) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
OAI221xp5_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1600), .B1(n_1602), .B2(n_1640), .C(n_1643), .Y(n_1385) );
AOI211xp5_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1512), .B(n_1516), .C(n_1575), .Y(n_1386) );
NAND5xp2_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1447), .C(n_1463), .D(n_1482), .E(n_1504), .Y(n_1387) );
AOI211xp5_ASAP7_75t_L g1388 ( .A1(n_1389), .A2(n_1419), .B(n_1428), .C(n_1440), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1404), .Y(n_1389) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1390), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1390), .B(n_1406), .Y(n_1457) );
AOI311xp33_ASAP7_75t_L g1482 ( .A1(n_1390), .A2(n_1483), .A3(n_1488), .B(n_1492), .C(n_1500), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1508 ( .A(n_1390), .B(n_1441), .Y(n_1508) );
OR2x2_ASAP7_75t_L g1534 ( .A(n_1390), .B(n_1535), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1390), .B(n_1415), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1390), .B(n_1411), .Y(n_1573) );
OR2x2_ASAP7_75t_L g1590 ( .A(n_1390), .B(n_1411), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1399), .Y(n_1390) );
AND2x4_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1394), .Y(n_1392) );
AND2x6_ASAP7_75t_L g1397 ( .A(n_1393), .B(n_1398), .Y(n_1397) );
AND2x6_ASAP7_75t_L g1400 ( .A(n_1393), .B(n_1401), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1393), .B(n_1403), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1393), .B(n_1403), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1393), .B(n_1403), .Y(n_1514) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1393), .B(n_1394), .Y(n_1601) );
HB1xp67_ASAP7_75t_L g1654 ( .A(n_1394), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1396), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1409), .Y(n_1404) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1405), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1405), .B(n_1490), .Y(n_1489) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_1405), .B(n_1445), .Y(n_1501) );
OAI21xp33_ASAP7_75t_L g1522 ( .A1(n_1405), .A2(n_1523), .B(n_1524), .Y(n_1522) );
OAI332xp33_ASAP7_75t_L g1567 ( .A1(n_1405), .A2(n_1508), .A3(n_1568), .B1(n_1570), .B2(n_1571), .B3(n_1572), .C1(n_1573), .C2(n_1574), .Y(n_1567) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1405), .B(n_1569), .Y(n_1568) );
CKINVDCx5p33_ASAP7_75t_R g1405 ( .A(n_1406), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1466 ( .A(n_1406), .B(n_1467), .Y(n_1466) );
INVx3_ASAP7_75t_L g1471 ( .A(n_1406), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1406), .B(n_1499), .Y(n_1505) );
NOR2xp33_ASAP7_75t_L g1531 ( .A(n_1406), .B(n_1474), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1535 ( .A(n_1406), .B(n_1409), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1589 ( .A(n_1406), .B(n_1590), .Y(n_1589) );
AND2x4_ASAP7_75t_SL g1406 ( .A(n_1407), .B(n_1408), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1409), .B(n_1457), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1415), .Y(n_1409) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1410), .B(n_1416), .Y(n_1441) );
AOI322xp5_ASAP7_75t_L g1504 ( .A1(n_1410), .A2(n_1490), .A3(n_1505), .B1(n_1506), .B2(n_1507), .C1(n_1509), .C2(n_1511), .Y(n_1504) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1411), .B(n_1416), .Y(n_1439) );
NOR2xp33_ASAP7_75t_L g1455 ( .A(n_1411), .B(n_1456), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1411), .B(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1411), .B(n_1438), .Y(n_1526) );
NOR3xp33_ASAP7_75t_SL g1560 ( .A(n_1411), .B(n_1436), .C(n_1512), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1413), .Y(n_1411) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1416), .Y(n_1469) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1416), .Y(n_1475) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1416), .B(n_1438), .Y(n_1569) );
NAND2x1_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1419), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1424), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1421), .Y(n_1443) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1421), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1421), .B(n_1424), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1421), .B(n_1425), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1423), .Y(n_1421) );
OR2x2_ASAP7_75t_L g1478 ( .A(n_1424), .B(n_1430), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1424), .B(n_1431), .Y(n_1491) );
HB1xp67_ASAP7_75t_SL g1540 ( .A(n_1424), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_1424), .B(n_1529), .Y(n_1572) );
CKINVDCx5p33_ASAP7_75t_R g1424 ( .A(n_1425), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1425), .B(n_1446), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1450 ( .A(n_1425), .B(n_1431), .Y(n_1450) );
HB1xp67_ASAP7_75t_SL g1476 ( .A(n_1425), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1425), .B(n_1443), .Y(n_1511) );
AND2x4_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1427), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1434), .Y(n_1428) );
OAI32xp33_ASAP7_75t_L g1564 ( .A1(n_1429), .A2(n_1430), .A3(n_1494), .B1(n_1524), .B2(n_1565), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1574 ( .A(n_1429), .B(n_1460), .Y(n_1574) );
INVx2_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1430), .B(n_1510), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1430), .B(n_1547), .Y(n_1580) );
INVx2_ASAP7_75t_SL g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1431), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1431), .B(n_1471), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1433), .Y(n_1431) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
O2A1O1Ixp33_ASAP7_75t_L g1530 ( .A1(n_1435), .A2(n_1531), .B(n_1532), .C(n_1533), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1437), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1461 ( .A(n_1436), .B(n_1462), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g1447 ( .A1(n_1437), .A2(n_1448), .B1(n_1451), .B2(n_1455), .C(n_1458), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1439), .Y(n_1437) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1438), .B(n_1441), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1438), .B(n_1469), .Y(n_1468) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1438), .B(n_1474), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_1438), .B(n_1471), .Y(n_1481) );
OR2x2_ASAP7_75t_L g1519 ( .A(n_1438), .B(n_1520), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1438), .B(n_1487), .Y(n_1524) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1438), .B(n_1480), .Y(n_1583) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1439), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1439), .B(n_1457), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1439), .B(n_1471), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1442), .Y(n_1440) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1441), .Y(n_1486) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1442), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1444), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1443), .B(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1443), .Y(n_1499) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1443), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1443), .B(n_1498), .Y(n_1596) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1445), .Y(n_1523) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1445), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1446), .B(n_1465), .Y(n_1464) );
INVx2_ASAP7_75t_L g1498 ( .A(n_1446), .Y(n_1498) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1449), .B(n_1453), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1449), .B(n_1471), .Y(n_1563) );
INVx2_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
NOR2xp33_ASAP7_75t_L g1598 ( .A(n_1450), .B(n_1471), .Y(n_1598) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
OAI332xp33_ASAP7_75t_L g1549 ( .A1(n_1454), .A2(n_1489), .A3(n_1535), .B1(n_1550), .B2(n_1551), .B3(n_1552), .C1(n_1553), .C2(n_1556), .Y(n_1549) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1457), .B(n_1487), .Y(n_1494) );
NOR2xp33_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1461), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
AOI21xp33_ASAP7_75t_L g1500 ( .A1(n_1462), .A2(n_1501), .B(n_1502), .Y(n_1500) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1462), .Y(n_1545) );
AOI221xp5_ASAP7_75t_L g1463 ( .A1(n_1464), .A2(n_1466), .B1(n_1470), .B2(n_1476), .C(n_1477), .Y(n_1463) );
OAI31xp33_ASAP7_75t_L g1576 ( .A1(n_1465), .A2(n_1518), .A3(n_1577), .B(n_1579), .Y(n_1576) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
A2O1A1Ixp33_ASAP7_75t_L g1597 ( .A1(n_1469), .A2(n_1557), .B(n_1598), .C(n_1599), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
NOR2xp33_ASAP7_75t_L g1527 ( .A(n_1471), .B(n_1478), .Y(n_1527) );
CKINVDCx14_ASAP7_75t_R g1544 ( .A(n_1471), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1472), .B(n_1498), .Y(n_1578) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1474), .Y(n_1487) );
A2O1A1Ixp33_ASAP7_75t_L g1517 ( .A1(n_1476), .A2(n_1518), .B(n_1521), .C(n_1529), .Y(n_1517) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1479), .Y(n_1477) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1478), .Y(n_1506) );
OAI22xp33_ASAP7_75t_L g1586 ( .A1(n_1478), .A2(n_1495), .B1(n_1502), .B2(n_1587), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1481), .Y(n_1479) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1481), .Y(n_1496) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1487), .Y(n_1485) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1486), .B(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1490), .Y(n_1548) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1537 ( .A(n_1491), .B(n_1538), .Y(n_1537) );
AOI21xp5_ASAP7_75t_L g1492 ( .A1(n_1493), .A2(n_1495), .B(n_1497), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
OAI22xp5_ASAP7_75t_L g1533 ( .A1(n_1497), .A2(n_1534), .B1(n_1536), .B2(n_1537), .Y(n_1533) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1497), .Y(n_1584) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1499), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1498), .B(n_1499), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1498), .B(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1498), .Y(n_1571) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1506), .B(n_1507), .Y(n_1528) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
NOR2xp33_ASAP7_75t_SL g1556 ( .A(n_1511), .B(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1511), .Y(n_1591) );
INVx3_ASAP7_75t_L g1529 ( .A(n_1512), .Y(n_1529) );
NOR2xp33_ASAP7_75t_L g1557 ( .A(n_1512), .B(n_1538), .Y(n_1557) );
NOR3xp33_ASAP7_75t_L g1588 ( .A(n_1512), .B(n_1589), .C(n_1591), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1515), .Y(n_1512) );
NAND4xp25_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1530), .C(n_1539), .D(n_1558), .Y(n_1516) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_1518), .A2(n_1547), .B1(n_1593), .B2(n_1596), .Y(n_1592) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1520), .Y(n_1565) );
NAND3xp33_ASAP7_75t_SL g1521 ( .A(n_1522), .B(n_1525), .C(n_1528), .Y(n_1521) );
INVx2_ASAP7_75t_L g1536 ( .A(n_1524), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1524), .B(n_1544), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1527), .Y(n_1525) );
CKINVDCx14_ASAP7_75t_R g1550 ( .A(n_1526), .Y(n_1550) );
CKINVDCx14_ASAP7_75t_R g1551 ( .A(n_1529), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1529), .B(n_1538), .Y(n_1566) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1537), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1593 ( .A(n_1537), .B(n_1594), .Y(n_1593) );
AOI211xp5_ASAP7_75t_L g1539 ( .A1(n_1540), .A2(n_1541), .B(n_1542), .C(n_1549), .Y(n_1539) );
AOI21xp33_ASAP7_75t_L g1542 ( .A1(n_1543), .A2(n_1546), .B(n_1548), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1545), .Y(n_1543) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
CKINVDCx14_ASAP7_75t_R g1585 ( .A(n_1551), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
OAI21xp5_ASAP7_75t_L g1561 ( .A1(n_1554), .A2(n_1562), .B(n_1564), .Y(n_1561) );
INVxp67_ASAP7_75t_SL g1570 ( .A(n_1557), .Y(n_1570) );
AOI221xp5_ASAP7_75t_L g1558 ( .A1(n_1559), .A2(n_1560), .B1(n_1561), .B2(n_1566), .C(n_1567), .Y(n_1558) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
NAND4xp25_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1581), .C(n_1592), .D(n_1597), .Y(n_1575) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
AOI311xp33_ASAP7_75t_L g1581 ( .A1(n_1582), .A2(n_1584), .A3(n_1585), .B(n_1586), .C(n_1588), .Y(n_1581) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1587), .Y(n_1599) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
BUFx2_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
HB1xp67_ASAP7_75t_L g1650 ( .A(n_1605), .Y(n_1650) );
NAND3xp33_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1625), .C(n_1633), .Y(n_1605) );
NOR2xp33_ASAP7_75t_SL g1606 ( .A(n_1607), .B(n_1620), .Y(n_1606) );
CKINVDCx5p33_ASAP7_75t_R g1640 ( .A(n_1641), .Y(n_1640) );
HB1xp67_ASAP7_75t_SL g1644 ( .A(n_1645), .Y(n_1644) );
BUFx3_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
INVxp33_ASAP7_75t_SL g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
HB1xp67_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
OAI21xp5_ASAP7_75t_L g1652 ( .A1(n_1653), .A2(n_1654), .B(n_1655), .Y(n_1652) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
endmodule