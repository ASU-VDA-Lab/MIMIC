module fake_netlist_5_1877_n_758 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_758);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_758;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_685;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_736;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_174;
wire n_745;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

BUFx5_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_47),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_85),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_86),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_40),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_36),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_27),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_60),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_79),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_51),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_41),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_99),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_50),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_33),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_92),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_100),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

BUFx2_ASAP7_75t_SL g180 ( 
.A(n_107),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_26),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_72),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_8),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_15),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_120),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_35),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_121),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_73),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_15),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_62),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_101),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_24),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_54),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_9),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_205),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_191),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_18),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_192),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_3),
.B(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_150),
.B(n_4),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_19),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

BUFx8_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_247),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_R g253 ( 
.A(n_220),
.B(n_201),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_170),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_161),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_246),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_220),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_5),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_R g266 ( 
.A(n_245),
.B(n_162),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_230),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_R g272 ( 
.A(n_245),
.B(n_165),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_166),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_211),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_245),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_221),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_171),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_221),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_224),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_206),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_240),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_240),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_240),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_240),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_219),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_219),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_219),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_232),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_219),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_226),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_226),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_234),
.C(n_215),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_243),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_243),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_243),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_282),
.B(n_215),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_293),
.B(n_173),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

AO221x1_ASAP7_75t_L g312 ( 
.A1(n_268),
.A2(n_222),
.B1(n_238),
.B2(n_241),
.C(n_226),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_265),
.B(n_174),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_222),
.B(n_216),
.C(n_235),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_216),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_238),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_238),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_238),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_222),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_241),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_241),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_241),
.Y(n_327)
);

BUFx8_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_175),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_176),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_210),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_233),
.B(n_235),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_273),
.B(n_229),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_208),
.C(n_181),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_271),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_279),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_273),
.B(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_260),
.A2(n_229),
.B(n_208),
.C(n_217),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_272),
.B(n_210),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_269),
.B(n_182),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_210),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_275),
.B(n_187),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_250),
.B(n_188),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_275),
.B(n_193),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

BUFx8_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_257),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_258),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_282),
.A2(n_233),
.B1(n_195),
.B2(n_203),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_252),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_252),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_282),
.B(n_217),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_212),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_282),
.B(n_217),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_268),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_280),
.B(n_196),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_202),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_233),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

OAI221xp5_ASAP7_75t_L g371 ( 
.A1(n_302),
.A2(n_227),
.B1(n_225),
.B2(n_213),
.C(n_212),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_213),
.B1(n_212),
.B2(n_227),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

NAND3xp33_ASAP7_75t_SL g375 ( 
.A(n_348),
.B(n_5),
.C(n_6),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_304),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_20),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

NOR2x2_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_6),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_315),
.B(n_213),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_315),
.B(n_213),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_225),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

NOR3xp33_ASAP7_75t_SL g391 ( 
.A(n_347),
.B(n_7),
.C(n_8),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_308),
.B(n_225),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_21),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_308),
.A2(n_227),
.B1(n_225),
.B2(n_11),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_322),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_356),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_322),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_334),
.A2(n_227),
.B1(n_9),
.B2(n_11),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_339),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_305),
.A2(n_307),
.B1(n_306),
.B2(n_309),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_350),
.B(n_7),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_310),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_22),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_361),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_23),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

OR2x6_ASAP7_75t_L g412 ( 
.A(n_326),
.B(n_12),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_321),
.A2(n_82),
.B1(n_147),
.B2(n_145),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_320),
.B(n_25),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_325),
.B(n_12),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_324),
.B(n_361),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_314),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_323),
.B(n_28),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_334),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_313),
.B(n_14),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_312),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_303),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_330),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_402),
.B(n_337),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_349),
.B(n_331),
.Y(n_435)
);

OR2x6_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_353),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_402),
.B(n_328),
.Y(n_438)
);

OA22x2_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_328),
.B1(n_352),
.B2(n_16),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_396),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_352),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_405),
.B(n_29),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_397),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_409),
.B(n_34),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_392),
.A2(n_37),
.B(n_38),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_400),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_409),
.B(n_44),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_380),
.A2(n_381),
.B(n_413),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_417),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_45),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_46),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_378),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_379),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_413),
.A2(n_48),
.B(n_49),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_53),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_R g460 ( 
.A(n_399),
.B(n_55),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_422),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_425),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_419),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_422),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_412),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_386),
.A2(n_65),
.B(n_66),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_388),
.A2(n_67),
.B(n_68),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_369),
.A2(n_70),
.B(n_71),
.C(n_75),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_420),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_424),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_390),
.A2(n_80),
.B(n_81),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_376),
.Y(n_474)
);

AOI22x1_ASAP7_75t_L g475 ( 
.A1(n_428),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_383),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_427),
.A2(n_90),
.B(n_91),
.C(n_93),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_377),
.B(n_94),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_410),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_367),
.B(n_407),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_385),
.B(n_103),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_434),
.A2(n_423),
.B(n_416),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_448),
.Y(n_487)
);

INVx6_ASAP7_75t_SL g488 ( 
.A(n_436),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_449),
.A2(n_435),
.B(n_459),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_408),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_433),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_455),
.A2(n_408),
.B(n_372),
.Y(n_492)
);

INVx3_ASAP7_75t_SL g493 ( 
.A(n_440),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_431),
.B(n_394),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_390),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_453),
.A2(n_411),
.B(n_387),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_464),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_393),
.B(n_371),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_480),
.A2(n_414),
.B(n_395),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_458),
.A2(n_395),
.B(n_372),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_438),
.A2(n_375),
.B(n_394),
.Y(n_502)
);

NAND2x1p5_ASAP7_75t_L g503 ( 
.A(n_464),
.B(n_479),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_457),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_436),
.B(n_415),
.Y(n_505)
);

AO21x2_ASAP7_75t_L g506 ( 
.A1(n_469),
.A2(n_391),
.B(n_393),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_479),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_430),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

AO21x2_ASAP7_75t_L g511 ( 
.A1(n_444),
.A2(n_447),
.B(n_462),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_467),
.A2(n_393),
.B(n_429),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

AO21x2_ASAP7_75t_L g514 ( 
.A1(n_478),
.A2(n_385),
.B(n_429),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_452),
.B(n_412),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_452),
.B(n_412),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_466),
.A2(n_104),
.B(n_105),
.Y(n_517)
);

INVx3_ASAP7_75t_SL g518 ( 
.A(n_439),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_468),
.A2(n_445),
.B(n_463),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_475),
.A2(n_106),
.B(n_110),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_471),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_470),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_473),
.A2(n_115),
.B(n_116),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_474),
.B(n_118),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_476),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_450),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_502),
.A2(n_442),
.B1(n_446),
.B2(n_472),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_487),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_494),
.B(n_483),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_497),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_524),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_507),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_465),
.B1(n_443),
.B2(n_441),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_513),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_489),
.A2(n_481),
.B(n_460),
.Y(n_541)
);

INVx8_ASAP7_75t_L g542 ( 
.A(n_513),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_484),
.A2(n_149),
.B(n_119),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_526),
.Y(n_544)
);

AOI21x1_ASAP7_75t_L g545 ( 
.A1(n_499),
.A2(n_122),
.B(n_123),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_498),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_492),
.B(n_124),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_521),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_509),
.B(n_125),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_490),
.Y(n_553)
);

AOI21x1_ASAP7_75t_L g554 ( 
.A1(n_499),
.A2(n_484),
.B(n_496),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_493),
.Y(n_555)
);

NAND2x1p5_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_126),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_513),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_493),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_503),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_504),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_520),
.Y(n_562)
);

BUFx2_ASAP7_75t_SL g563 ( 
.A(n_522),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_498),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_492),
.A2(n_128),
.B(n_129),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_508),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_501),
.B(n_131),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_518),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_559),
.B(n_518),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_555),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_535),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_511),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_531),
.B(n_508),
.Y(n_574)
);

AND2x4_ASAP7_75t_SL g575 ( 
.A(n_564),
.B(n_505),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_533),
.B(n_511),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_536),
.B(n_490),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_538),
.A2(n_516),
.B1(n_515),
.B2(n_505),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_546),
.B(n_510),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_546),
.B(n_516),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_536),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_515),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_561),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_529),
.A2(n_506),
.B1(n_505),
.B2(n_500),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_561),
.A2(n_504),
.B1(n_506),
.B2(n_527),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_544),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_565),
.A2(n_525),
.B1(n_514),
.B2(n_527),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_548),
.A2(n_488),
.B1(n_525),
.B2(n_514),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_548),
.A2(n_512),
.B(n_503),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_555),
.B(n_495),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_559),
.Y(n_593)
);

NOR2x1p5_ASAP7_75t_L g594 ( 
.A(n_551),
.B(n_522),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_542),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_530),
.B(n_485),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_495),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_560),
.B(n_488),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_560),
.B(n_138),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_563),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_539),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_547),
.B(n_139),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_547),
.B(n_140),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_568),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_549),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_542),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_540),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_537),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_540),
.B(n_558),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_540),
.B(n_558),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_543),
.A2(n_563),
.B1(n_567),
.B2(n_556),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

INVx8_ASAP7_75t_L g615 ( 
.A(n_542),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_608),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_584),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_597),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_602),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_573),
.B(n_567),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_576),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_574),
.B(n_573),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_606),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_582),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_583),
.B(n_553),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_543),
.Y(n_626)
);

AND2x4_ASAP7_75t_SL g627 ( 
.A(n_608),
.B(n_580),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_609),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_588),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_577),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_553),
.Y(n_632)
);

OAI33xp33_ASAP7_75t_L g633 ( 
.A1(n_572),
.A2(n_550),
.A3(n_557),
.B1(n_552),
.B2(n_562),
.B3(n_545),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_596),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_575),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_587),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_570),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_579),
.B(n_537),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_587),
.B(n_554),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_578),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_599),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_578),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_579),
.B(n_558),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_610),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_614),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_603),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_612),
.B(n_562),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_586),
.B(n_591),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_604),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_585),
.B(n_542),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_557),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_594),
.B(n_556),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_600),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_571),
.B(n_534),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_622),
.B(n_640),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_618),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_599),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_619),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_SL g660 ( 
.A1(n_637),
.A2(n_605),
.B1(n_590),
.B2(n_589),
.C(n_613),
.Y(n_660)
);

OR2x6_ASAP7_75t_SL g661 ( 
.A(n_655),
.B(n_593),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_641),
.B(n_592),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_652),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_625),
.B(n_601),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_640),
.B(n_600),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_617),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_655),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_620),
.B(n_592),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_592),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_623),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_623),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_628),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_647),
.B(n_569),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_627),
.B(n_632),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_628),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_621),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_627),
.B(n_607),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_624),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_637),
.B(n_615),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_643),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_630),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_656),
.B(n_663),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_656),
.B(n_638),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_671),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_673),
.B(n_653),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_663),
.B(n_652),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_658),
.B(n_626),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_657),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_659),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_667),
.B(n_626),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_671),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_676),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_667),
.B(n_620),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_678),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_668),
.B(n_649),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_682),
.B(n_680),
.Y(n_697)
);

OA222x2_ASAP7_75t_L g698 ( 
.A1(n_696),
.A2(n_679),
.B1(n_649),
.B2(n_662),
.C1(n_631),
.C2(n_681),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_694),
.B(n_674),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_689),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_R g701 ( 
.A1(n_697),
.A2(n_664),
.B(n_644),
.C(n_639),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_683),
.B(n_669),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_690),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_687),
.B(n_679),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_693),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_683),
.B(n_675),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_700),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_703),
.Y(n_708)
);

OAI221xp5_ASAP7_75t_L g709 ( 
.A1(n_701),
.A2(n_686),
.B1(n_660),
.B2(n_704),
.C(n_705),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_706),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_701),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_702),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_712),
.B(n_635),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_710),
.B(n_704),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_711),
.B(n_684),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_SL g717 ( 
.A1(n_709),
.A2(n_686),
.B(n_665),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_SL g719 ( 
.A(n_717),
.B(n_660),
.C(n_651),
.Y(n_719)
);

OAI221xp5_ASAP7_75t_L g720 ( 
.A1(n_714),
.A2(n_708),
.B1(n_695),
.B2(n_697),
.C(n_635),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_716),
.B(n_661),
.Y(n_721)
);

AOI211xp5_ASAP7_75t_L g722 ( 
.A1(n_713),
.A2(n_698),
.B(n_650),
.C(n_661),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_722),
.A2(n_665),
.B1(n_679),
.B2(n_669),
.Y(n_723)
);

NAND4xp25_ASAP7_75t_L g724 ( 
.A(n_718),
.B(n_642),
.C(n_632),
.D(n_669),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_724),
.A2(n_721),
.B(n_719),
.C(n_720),
.Y(n_725)
);

OAI221xp5_ASAP7_75t_L g726 ( 
.A1(n_723),
.A2(n_642),
.B1(n_647),
.B2(n_654),
.C(n_692),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_723),
.A2(n_692),
.B1(n_685),
.B2(n_666),
.C(n_670),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_725),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_726),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_SL g730 ( 
.A1(n_727),
.A2(n_636),
.B(n_634),
.C(n_654),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_726),
.B(n_699),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_725),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_725),
.B(n_616),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_733),
.B(n_685),
.Y(n_734)
);

NOR3xp33_ASAP7_75t_L g735 ( 
.A(n_728),
.B(n_598),
.C(n_541),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_732),
.B(n_541),
.C(n_645),
.Y(n_736)
);

NOR4xp25_ASAP7_75t_L g737 ( 
.A(n_729),
.B(n_629),
.C(n_672),
.D(n_646),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_SL g738 ( 
.A(n_731),
.B(n_677),
.C(n_691),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_737),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_738),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_734),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_735),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_740),
.A2(n_736),
.B1(n_730),
.B2(n_632),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_741),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_739),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_742),
.B1(n_595),
.B2(n_616),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_616),
.B1(n_595),
.B2(n_646),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_743),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_748),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_746),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_747),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_748),
.A2(n_616),
.B1(n_595),
.B2(n_615),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_L g753 ( 
.A1(n_746),
.A2(n_615),
.B1(n_616),
.B2(n_646),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_749),
.Y(n_754)
);

OAI21xp33_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_752),
.B(n_750),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_751),
.B1(n_753),
.B2(n_688),
.Y(n_756)
);

OR2x6_ASAP7_75t_L g757 ( 
.A(n_756),
.B(n_648),
.Y(n_757)
);

AOI211xp5_ASAP7_75t_L g758 ( 
.A1(n_757),
.A2(n_675),
.B(n_681),
.C(n_633),
.Y(n_758)
);


endmodule