module real_jpeg_5751_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_1),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_1),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_2),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_2),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_2),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_3),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_3),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_3),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_3),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_3),
.B(n_152),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_3),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_3),
.B(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_4),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_4),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_5),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_5),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_5),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_5),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_5),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_5),
.B(n_454),
.Y(n_453)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_7),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_8),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_8),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_8),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_8),
.B(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_9),
.Y(n_228)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_11),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_11),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_11),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_152),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_12),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_12),
.Y(n_211)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_12),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_12),
.Y(n_300)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_13),
.Y(n_285)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_13),
.Y(n_439)
);

BUFx5_ASAP7_75t_L g454 ( 
.A(n_13),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_14),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_14),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_14),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_14),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_15),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_15),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_15),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_15),
.B(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_163),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_162),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_20),
.B(n_102),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_47),
.B2(n_48),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_44),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_30),
.B(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.C(n_40),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_31),
.A2(n_37),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_31),
.Y(n_140)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_35),
.Y(n_270)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_36),
.Y(n_249)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_37),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_37),
.A2(n_139),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_37),
.B(n_144),
.C(n_188),
.Y(n_337)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_39),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_40),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_40),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_44),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_44),
.A2(n_86),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_44),
.B(n_355),
.C(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_44),
.A2(n_86),
.B1(n_151),
.B2(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_46),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_46),
.Y(n_258)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_70),
.B2(n_71),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_62),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_88),
.C(n_93),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_62),
.B1(n_63),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_55),
.A2(n_93),
.B1(n_94),
.B2(n_101),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_55),
.A2(n_101),
.B1(n_231),
.B2(n_239),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_55),
.B(n_117),
.C(n_232),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_57),
.Y(n_395)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_57),
.Y(n_412)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_58),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_63),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_62),
.A2(n_63),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_63),
.B(n_205),
.C(n_210),
.Y(n_297)
);

OR2x2_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_66),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_66),
.Y(n_323)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_76),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_95),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_67),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_81),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_74),
.A2(n_75),
.B1(n_279),
.B2(n_286),
.Y(n_278)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_75),
.B(n_357),
.C(n_358),
.Y(n_356)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_81),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_78),
.B(n_128),
.C(n_135),
.Y(n_157)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_99),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_83),
.A2(n_84),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_143),
.C(n_151),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_87),
.B(n_99),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_94),
.B1(n_111),
.B2(n_115),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_93),
.A2(n_94),
.B1(n_188),
.B2(n_290),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_107),
.C(n_111),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_94),
.B(n_183),
.C(n_188),
.Y(n_182)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_97),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_98),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_98),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_153),
.C(n_159),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_103),
.B(n_153),
.CI(n_159),
.CON(n_499),
.SN(n_499)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_136),
.C(n_142),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_104),
.A2(n_105),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.C(n_125),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_106),
.B(n_366),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_144),
.C(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_111),
.B(n_316),
.C(n_321),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_111),
.A2(n_115),
.B1(n_144),
.B2(n_291),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_111),
.A2(n_115),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_112),
.Y(n_429)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_113),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_116),
.B(n_125),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_121),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_117),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_117),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_117),
.A2(n_237),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_120),
.B(n_121),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_124),
.Y(n_422)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_132),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_132),
.B(n_264),
.C(n_267),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_136),
.B(n_142),
.Y(n_502)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_143),
.B(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_144),
.A2(n_188),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_144),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_144),
.A2(n_291),
.B1(n_405),
.B2(n_406),
.Y(n_423)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_147),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_147),
.Y(n_344)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_150),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_151),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_158),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_154),
.A2(n_155),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_157),
.B(n_158),
.Y(n_506)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_497),
.B(n_511),
.Y(n_163)
);

AO21x2_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_361),
.B(n_377),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_331),
.B(n_360),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_306),
.B(n_330),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_167),
.B(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_272),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_168),
.B(n_272),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_229),
.C(n_259),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_169),
.B(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_201),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_170),
.B(n_202),
.C(n_213),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_182),
.C(n_191),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_171),
.B(n_326),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_171),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_176),
.CI(n_180),
.CON(n_171),
.SN(n_171)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_172),
.B(n_176),
.C(n_180),
.Y(n_271)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_182),
.A2(n_191),
.B1(n_192),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_182),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_183),
.B(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_188),
.Y(n_290)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_324)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_196),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_196),
.Y(n_448)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_213),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_205),
.A2(n_212),
.B1(n_245),
.B2(n_246),
.Y(n_413)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_215),
.B(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_214),
.B(n_222),
.C(n_224),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_220),
.B(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_225),
.B(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_225),
.B(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_225),
.B(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_229),
.B(n_259),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_240),
.C(n_242),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_230),
.A2(n_240),
.B1(n_241),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_242),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.C(n_255),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_243),
.A2(n_244),
.B1(n_484),
.B2(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_250),
.A2(n_251),
.B1(n_255),
.B2(n_256),
.Y(n_485)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_262),
.C(n_271),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_275),
.C(n_305),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_292),
.B1(n_304),
.B2(n_305),
.Y(n_274)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_287),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_277),
.B(n_278),
.C(n_287),
.Y(n_348)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_284),
.Y(n_358)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_291),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_301),
.C(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_328),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_307),
.B(n_328),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.C(n_325),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_308),
.A2(n_309),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_312),
.B(n_325),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_324),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_313),
.B(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_315),
.B(n_324),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_316),
.A2(n_317),
.B1(n_321),
.B2(n_322),
.Y(n_402)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_332),
.B(n_361),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_334),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_362),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_334),
.B(n_362),
.Y(n_496)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_347),
.CI(n_359),
.CON(n_334),
.SN(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_343),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_336)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_337),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_342),
.C(n_343),
.Y(n_369)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_350),
.C(n_352),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_363),
.B(n_365),
.C(n_367),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_370),
.B2(n_376),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_368),
.B(n_371),
.C(n_373),
.Y(n_507)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

OAI31xp33_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_493),
.A3(n_494),
.B(n_496),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_487),
.B(n_492),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_472),
.B(n_486),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_424),
.B(n_471),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_414),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_382),
.B(n_414),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_403),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_400),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_384),
.B(n_400),
.C(n_403),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_391),
.C(n_396),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_385),
.A2(n_386),
.B1(n_391),
.B2(n_392),
.Y(n_416)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_396),
.B(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_409),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_404),
.B(n_481),
.C(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_413),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_417),
.C(n_423),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_415),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_417),
.A2(n_423),
.B1(n_463),
.B2(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_465),
.B(n_470),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_450),
.B(n_464),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_434),
.B(n_449),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_445),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_445),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_440),
.B(n_444),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_440),
.Y(n_444)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_444),
.A2(n_452),
.B1(n_458),
.B2(n_459),
.Y(n_451)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx8_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_460),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_460),
.Y(n_464)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_452),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_453),
.A2(n_455),
.B(n_458),
.Y(n_466)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_462),
.B(n_463),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_466),
.B(n_467),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_474),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_476),
.B1(n_478),
.B2(n_479),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_480),
.C(n_483),
.Y(n_488)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.Y(n_479)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_489),
.Y(n_492)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_508),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_498),
.A2(n_512),
.B(n_513),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_500),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_499),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.C(n_507),
.Y(n_500)
);

FAx1_ASAP7_75t_SL g510 ( 
.A(n_501),
.B(n_504),
.CI(n_507),
.CON(n_510),
.SN(n_510)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_502),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_510),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_510),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_510),
.Y(n_517)
);


endmodule