module fake_jpeg_17662_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_19),
.B1(n_24),
.B2(n_27),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_54),
.B1(n_58),
.B2(n_65),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_24),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_56),
.B1(n_62),
.B2(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_19),
.B1(n_27),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_33),
.B1(n_23),
.B2(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_38),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_30),
.B1(n_21),
.B2(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_77),
.B1(n_82),
.B2(n_35),
.Y(n_128)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_74),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.C(n_43),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_75),
.C(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_23),
.B1(n_20),
.B2(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_81),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_1),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_35),
.B1(n_20),
.B2(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_38),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_23),
.B1(n_28),
.B2(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_40),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_89),
.Y(n_105)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_52),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_43),
.B1(n_63),
.B2(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_47),
.B1(n_64),
.B2(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_33),
.B1(n_28),
.B2(n_34),
.Y(n_125)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_102),
.Y(n_106)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_43),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_43),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_54),
.B1(n_46),
.B2(n_63),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_111),
.A2(n_130),
.B1(n_101),
.B2(n_35),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_18),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_107),
.B(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_128),
.B1(n_71),
.B2(n_103),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_34),
.B1(n_33),
.B2(n_18),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_73),
.B1(n_91),
.B2(n_67),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_12),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_94),
.B1(n_80),
.B2(n_69),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_138),
.A2(n_145),
.B1(n_156),
.B2(n_162),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_72),
.C(n_75),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_141),
.C(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_78),
.C(n_100),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_81),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_131),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_66),
.B(n_86),
.C(n_73),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_147),
.B(n_159),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_78),
.B1(n_93),
.B2(n_66),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_86),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_105),
.A2(n_99),
.B1(n_98),
.B2(n_83),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_149),
.A2(n_113),
.B1(n_39),
.B2(n_35),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_157),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_111),
.C(n_108),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_160),
.B1(n_147),
.B2(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_70),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_155),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_43),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_161),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_85),
.B(n_90),
.C(n_84),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_39),
.C(n_44),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_106),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_39),
.C(n_44),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_121),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_18),
.B(n_35),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_129),
.C(n_132),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g221 ( 
.A1(n_165),
.A2(n_195),
.B(n_17),
.Y(n_221)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_176),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_185),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_177),
.B1(n_162),
.B2(n_159),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_120),
.B1(n_133),
.B2(n_124),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_167),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_191),
.C(n_192),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_115),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_109),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_109),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_135),
.A2(n_113),
.B(n_31),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_150),
.B(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_136),
.B1(n_160),
.B2(n_135),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_208),
.B1(n_216),
.B2(n_221),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_137),
.B1(n_138),
.B2(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_161),
.C(n_156),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_191),
.C(n_166),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_169),
.B(n_182),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_219),
.Y(n_240)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_223),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_185),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_170),
.B(n_149),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_9),
.B(n_15),
.C(n_11),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_184),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_229),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_194),
.B1(n_183),
.B2(n_189),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_239),
.B1(n_217),
.B2(n_214),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_188),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_166),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_180),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_192),
.C(n_174),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_209),
.C(n_208),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_193),
.C(n_177),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_171),
.B1(n_187),
.B2(n_178),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_173),
.C(n_195),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_222),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_219),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_201),
.B1(n_198),
.B2(n_199),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_255),
.B1(n_261),
.B2(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_218),
.C(n_201),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_252),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_240),
.B1(n_238),
.B2(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_260),
.B1(n_262),
.B2(n_225),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_217),
.C(n_223),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_271),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_254),
.A2(n_215),
.B1(n_173),
.B2(n_220),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_266),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_246),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_259),
.B1(n_257),
.B2(n_249),
.Y(n_283)
);

AOI222xp33_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_197),
.B1(n_17),
.B2(n_39),
.C1(n_9),
.C2(n_10),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_9),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_17),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_3),
.C(n_4),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_275),
.C(n_257),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_3),
.C(n_4),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_245),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_282),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_286),
.C(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_269),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_264),
.B1(n_270),
.B2(n_267),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_4),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_253),
.C(n_6),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.C(n_295),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_274),
.B1(n_6),
.B2(n_7),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_7),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_5),
.C(n_6),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_277),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_284),
.B(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_287),
.B(n_277),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_5),
.B(n_7),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_295),
.C(n_296),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_292),
.B(n_301),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_308),
.A2(n_290),
.B(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_307),
.Y(n_312)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_305),
.A3(n_301),
.B(n_291),
.Y(n_313)
);


endmodule