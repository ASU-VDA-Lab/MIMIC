module fake_jpeg_15772_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_73),
.Y(n_75)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_82),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_55),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_59),
.B1(n_65),
.B2(n_51),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_66),
.B1(n_56),
.B2(n_64),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_50),
.B1(n_54),
.B2(n_60),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_58),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_107),
.B(n_91),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_52),
.Y(n_117)
);

AO21x2_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_94),
.B(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_116),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_98),
.B1(n_96),
.B2(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_119),
.CI(n_104),
.CON(n_122),
.SN(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_27),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_26),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_28),
.B(n_40),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_21),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_47),
.B(n_20),
.C(n_1),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_29),
.B(n_41),
.C(n_2),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_19),
.C(n_39),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_18),
.B1(n_35),
.B2(n_4),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_31),
.B(n_37),
.C(n_5),
.Y(n_134)
);


endmodule