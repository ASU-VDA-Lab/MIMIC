module fake_jpeg_21983_n_307 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NAND2x1_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_30),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g107 ( 
.A(n_50),
.B(n_10),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_23),
.B1(n_21),
.B2(n_37),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_65),
.B1(n_67),
.B2(n_33),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_19),
.B(n_30),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_23),
.B1(n_37),
.B2(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_23),
.B1(n_37),
.B2(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_22),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_27),
.B1(n_18),
.B2(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_66),
.B1(n_0),
.B2(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_22),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_18),
.B1(n_30),
.B2(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_31),
.B1(n_34),
.B2(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_79),
.B1(n_8),
.B2(n_14),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_27),
.B1(n_25),
.B2(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_10),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_28),
.B1(n_33),
.B2(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_1),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_87),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_33),
.B1(n_48),
.B2(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_80),
.B1(n_74),
.B2(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_94),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_101),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_91),
.B(n_6),
.Y(n_142)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_109),
.B1(n_112),
.B2(n_82),
.Y(n_144)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_61),
.B1(n_69),
.B2(n_68),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_102),
.B(n_110),
.C(n_9),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_106),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_7),
.C(n_9),
.Y(n_137)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_114),
.Y(n_143)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_69),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_118),
.B1(n_60),
.B2(n_63),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_17),
.B1(n_7),
.B2(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_128),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_77),
.B1(n_76),
.B2(n_66),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_125),
.B1(n_136),
.B2(n_145),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_3),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_127),
.A2(n_129),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_74),
.C(n_5),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_138),
.C(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_74),
.B1(n_6),
.B2(n_4),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_4),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_4),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_91),
.B(n_87),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_12),
.B1(n_13),
.B2(n_84),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_114),
.B1(n_102),
.B2(n_113),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_92),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_89),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_6),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_112),
.B1(n_95),
.B2(n_110),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_171),
.B1(n_176),
.B2(n_180),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_130),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_159),
.B(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_169),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_100),
.B(n_109),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_100),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_168),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_116),
.B1(n_83),
.B2(n_96),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_167),
.B1(n_133),
.B2(n_141),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_108),
.B1(n_89),
.B2(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_119),
.A2(n_106),
.B1(n_99),
.B2(n_94),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_134),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_7),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_91),
.B(n_115),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_127),
.B(n_149),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_86),
.B(n_84),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_179),
.B(n_137),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_134),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_154),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_12),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_119),
.A2(n_129),
.B1(n_124),
.B2(n_135),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_182),
.B(n_126),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_192),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_196),
.B1(n_168),
.B2(n_152),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_125),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_194),
.C(n_199),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_127),
.B(n_129),
.Y(n_195)
);

XOR2x2_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_173),
.Y(n_231)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_133),
.B1(n_136),
.B2(n_148),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_200),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_139),
.C(n_122),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_208),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_156),
.A2(n_141),
.B(n_147),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_205),
.B1(n_159),
.B2(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_122),
.B1(n_147),
.B2(n_126),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_142),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_165),
.Y(n_221)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_227),
.B1(n_232),
.B2(n_188),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_223),
.B1(n_230),
.B2(n_203),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_163),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_233),
.B(n_179),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_180),
.B1(n_176),
.B2(n_161),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_155),
.C(n_174),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_208),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_161),
.B1(n_166),
.B2(n_155),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_155),
.B1(n_160),
.B2(n_162),
.Y(n_230)
);

OA21x2_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_195),
.B(n_186),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_205),
.B1(n_187),
.B2(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_238),
.B1(n_244),
.B2(n_247),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_193),
.C(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_239),
.C(n_240),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_197),
.B1(n_188),
.B2(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_201),
.C(n_194),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_160),
.C(n_162),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_249),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_196),
.B(n_157),
.C(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_196),
.B1(n_184),
.B2(n_211),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_250),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_196),
.B1(n_211),
.B2(n_189),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_196),
.B1(n_207),
.B2(n_163),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_173),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

AO221x1_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_224),
.B1(n_212),
.B2(n_213),
.C(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_225),
.B(n_234),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_263),
.B(n_264),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_217),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_256),
.Y(n_269)
);

AO21x1_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_226),
.B(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

AO221x1_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_213),
.B1(n_123),
.B2(n_233),
.C(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_154),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_228),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_245),
.B1(n_243),
.B2(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_237),
.C(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_240),
.C(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_279),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_243),
.B1(n_236),
.B2(n_235),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_244),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_250),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_249),
.C(n_236),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_229),
.A3(n_214),
.B1(n_222),
.B2(n_218),
.C1(n_173),
.C2(n_230),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_285),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_259),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_286),
.B(n_288),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_218),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_259),
.C(n_255),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_284),
.B(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_278),
.B1(n_258),
.B2(n_275),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_279),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_269),
.C(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_258),
.C(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_229),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_260),
.A3(n_277),
.B1(n_257),
.B2(n_214),
.C1(n_179),
.C2(n_158),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_169),
.C(n_179),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_123),
.Y(n_307)
);


endmodule