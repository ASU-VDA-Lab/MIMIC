module fake_netlist_5_1340_n_1976 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1976);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1976;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_1014;
wire n_279;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_61),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_97),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_19),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_126),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_24),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_62),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_79),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_53),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_10),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_76),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_134),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_109),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_164),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_45),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_38),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_77),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_130),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_186),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_81),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_116),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_66),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_148),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_106),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_18),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_46),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_175),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_72),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_180),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_18),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_137),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_8),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_104),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_75),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_91),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_21),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_27),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_11),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_102),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_11),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_19),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_74),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_115),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_8),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_17),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_183),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_110),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_71),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_100),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_154),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_150),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_146),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_84),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_55),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_57),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_168),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_30),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_108),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_50),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_187),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_49),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_27),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_50),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_192),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_167),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_83),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_101),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_151),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_35),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_96),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_125),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_159),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_82),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_136),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_4),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_158),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_127),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_48),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_153),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_131),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_178),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_57),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_49),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_51),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_13),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_14),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_54),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_7),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_63),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_140),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_89),
.Y(n_328)
);

BUFx8_ASAP7_75t_SL g329 ( 
.A(n_44),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_6),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_53),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_32),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_87),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_70),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_44),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_118),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_36),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_138),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_95),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_43),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_59),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_161),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_68),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_193),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_40),
.Y(n_345)
);

BUFx10_ASAP7_75t_L g346 ( 
.A(n_30),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_93),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_33),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_3),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_17),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_47),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_62),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_42),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_56),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_10),
.Y(n_355)
);

BUFx5_ASAP7_75t_L g356 ( 
.A(n_86),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_43),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_65),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_52),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_157),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_144),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_16),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_34),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_9),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_56),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_60),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_32),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_133),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_73),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_64),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_0),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_4),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_149),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_112),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_121),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_60),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_155),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_98),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_185),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_14),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_21),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_22),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_55),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_36),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_141),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_78),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_135),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_94),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_99),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_59),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_182),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_33),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_173),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_80),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_207),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_207),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_207),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_207),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_206),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_207),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_207),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_207),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_214),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_207),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_206),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_329),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_354),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_238),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_245),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_249),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_354),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_267),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_255),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_222),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_202),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_222),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_212),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_229),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_234),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_356),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_241),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_250),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_258),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_270),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_259),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_278),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_289),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_297),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_197),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_247),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_298),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_231),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_374),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_305),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_307),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_320),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_325),
.Y(n_450)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_197),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_332),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_282),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_337),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_265),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_356),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_341),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_348),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_271),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_273),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_351),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_359),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_274),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_365),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_309),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_346),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_277),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_198),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_201),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_310),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_324),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_272),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_324),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_317),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_272),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_209),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_370),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_209),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_237),
.Y(n_481)
);

BUFx6f_ASAP7_75t_SL g482 ( 
.A(n_368),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_237),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_284),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_272),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_211),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_211),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_385),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_284),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_291),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_291),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_252),
.Y(n_492)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_346),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_269),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_316),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_204),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_356),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_301),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_230),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_407),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_407),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_399),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_230),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_423),
.B(n_316),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_395),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_445),
.B(n_304),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_395),
.B(n_347),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_399),
.B(n_199),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_413),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_402),
.B(n_253),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_399),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_399),
.B(n_199),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_492),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_396),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_431),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_397),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_414),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_412),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_487),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_406),
.B(n_368),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_406),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_402),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_415),
.A2(n_296),
.B1(n_380),
.B2(n_384),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_405),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_405),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_437),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_400),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_478),
.Y(n_547)
);

OA21x2_ASAP7_75t_L g548 ( 
.A1(n_478),
.A2(n_393),
.B(n_347),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_406),
.B(n_200),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_437),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_480),
.A2(n_393),
.B(n_213),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_481),
.A2(n_215),
.B(n_208),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_427),
.B(n_216),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

NOR2x1_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_224),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_403),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_483),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_404),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_497),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

INVx6_ASAP7_75t_L g566 ( 
.A(n_406),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_443),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_484),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_470),
.B(n_233),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_L g571 ( 
.A(n_406),
.B(n_218),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_489),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_410),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_489),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_490),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_498),
.A2(n_420),
.B1(n_460),
.B2(n_455),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_542),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_501),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_508),
.B(n_434),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_498),
.B(n_451),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_542),
.Y(n_582)
);

AO21x2_ASAP7_75t_L g583 ( 
.A1(n_515),
.A2(n_242),
.B(n_240),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_524),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_500),
.B(n_507),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_500),
.B(n_446),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_521),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_500),
.B(n_471),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_512),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_559),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_558),
.B(n_455),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_514),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_558),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_507),
.B(n_496),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_511),
.B(n_356),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_534),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_527),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_527),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_513),
.B(n_460),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_530),
.B(n_461),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_536),
.B(n_421),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_499),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_535),
.A2(n_227),
.B1(n_323),
.B2(n_319),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_512),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

AND3x1_ASAP7_75t_L g614 ( 
.A(n_541),
.B(n_425),
.C(n_421),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_559),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_537),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_537),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_520),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_559),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_546),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_546),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_517),
.B(n_243),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_521),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_535),
.A2(n_464),
.B1(n_468),
.B2(n_486),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_520),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_509),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_507),
.B(n_464),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_574),
.B(n_494),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g633 ( 
.A(n_562),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_543),
.B(n_410),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_543),
.B(n_268),
.C(n_468),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_509),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_517),
.B(n_368),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_551),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_551),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_559),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_559),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_517),
.B(n_200),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_508),
.B(n_425),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_551),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_509),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_555),
.Y(n_647)
);

NAND2x1p5_ASAP7_75t_L g648 ( 
.A(n_554),
.B(n_244),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_559),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_511),
.B(n_356),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

INVxp33_ASAP7_75t_L g652 ( 
.A(n_534),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_508),
.B(n_490),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_556),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_510),
.B(n_467),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_556),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_563),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_519),
.B(n_203),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_550),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_555),
.B(n_491),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_510),
.B(n_493),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_563),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_505),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_506),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_541),
.A2(n_312),
.B1(n_287),
.B2(n_290),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_536),
.A2(n_217),
.B1(n_321),
.B2(n_315),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_572),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_506),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_555),
.B(n_246),
.Y(n_671)
);

XOR2x2_ASAP7_75t_L g672 ( 
.A(n_550),
.B(n_519),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_505),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_509),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_499),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_518),
.B(n_436),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_571),
.B(n_440),
.C(n_439),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_506),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_506),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_518),
.B(n_441),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_522),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_523),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_523),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_572),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_570),
.A2(n_495),
.B1(n_491),
.B2(n_444),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_532),
.Y(n_687)
);

AND3x2_ASAP7_75t_L g688 ( 
.A(n_519),
.B(n_387),
.C(n_264),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_571),
.B(n_448),
.C(n_447),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_525),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_572),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_572),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_549),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_570),
.A2(n_495),
.B1(n_457),
.B2(n_454),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_549),
.B(n_482),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_525),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_562),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_528),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_528),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_565),
.B(n_449),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_572),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_529),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_531),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_531),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_565),
.B(n_482),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_539),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_509),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_570),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_526),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_515),
.B(n_221),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_499),
.B(n_299),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_572),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_565),
.B(n_482),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_572),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_526),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_540),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_568),
.B(n_473),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_540),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_526),
.Y(n_721)
);

NOR2x1p5_ASAP7_75t_L g722 ( 
.A(n_503),
.B(n_218),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_540),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_526),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_526),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_568),
.B(n_203),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_533),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_630),
.B(n_568),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_595),
.B(n_540),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_595),
.B(n_540),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_624),
.A2(n_294),
.B1(n_236),
.B2(n_355),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_581),
.B(n_453),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_599),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_608),
.Y(n_734)
);

NOR3xp33_ASAP7_75t_L g735 ( 
.A(n_597),
.B(n_452),
.C(n_450),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_610),
.B(n_570),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_610),
.B(n_540),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_SL g738 ( 
.A(n_586),
.B(n_554),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_693),
.B(n_540),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_664),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_710),
.B(n_552),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_580),
.B(n_466),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_577),
.B(n_557),
.C(n_570),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_693),
.B(n_544),
.Y(n_744)
);

AND2x6_ASAP7_75t_L g745 ( 
.A(n_695),
.B(n_248),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_602),
.B(n_472),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_624),
.B(n_205),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_664),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_580),
.B(n_647),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_673),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_719),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_647),
.B(n_712),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_652),
.B(n_476),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_673),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_647),
.B(n_205),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_647),
.B(n_544),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_587),
.B(n_544),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_676),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_632),
.B(n_458),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_592),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_632),
.B(n_459),
.Y(n_761)
);

INVx8_ASAP7_75t_L g762 ( 
.A(n_719),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_578),
.B(n_582),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_592),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_676),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_655),
.B(n_210),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_682),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_590),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_593),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_635),
.B(n_463),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_710),
.B(n_544),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_675),
.A2(n_538),
.B(n_504),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_671),
.B(n_544),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_682),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_593),
.Y(n_775)
);

BUFx6f_ASAP7_75t_SL g776 ( 
.A(n_579),
.Y(n_776)
);

BUFx8_ASAP7_75t_L g777 ( 
.A(n_589),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_643),
.B(n_479),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_658),
.B(n_488),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_589),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_677),
.B(n_544),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_645),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_662),
.B(n_210),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_671),
.B(n_544),
.Y(n_785)
);

AOI22x1_ASAP7_75t_L g786 ( 
.A1(n_648),
.A2(n_386),
.B1(n_342),
.B2(n_334),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_671),
.B(n_504),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_660),
.A2(n_591),
.B(n_600),
.C(n_653),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_726),
.B(n_532),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_671),
.B(n_504),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_671),
.A2(n_557),
.B1(n_261),
.B2(n_308),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_644),
.B(n_465),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_608),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_690),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_656),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_677),
.B(n_681),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_700),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_681),
.A2(n_251),
.B(n_257),
.C(n_391),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_700),
.B(n_219),
.Y(n_800)
);

NOR2x1p5_ASAP7_75t_L g801 ( 
.A(n_697),
.B(n_236),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_627),
.B(n_567),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_644),
.B(n_473),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_696),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_696),
.A2(n_302),
.B(n_377),
.C(n_375),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_706),
.B(n_219),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_614),
.A2(n_363),
.B1(n_330),
.B2(n_331),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_659),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_671),
.B(n_533),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_715),
.B(n_220),
.Y(n_810)
);

AO22x2_ASAP7_75t_L g811 ( 
.A1(n_638),
.A2(n_475),
.B1(n_318),
.B2(n_333),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_615),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_699),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_703),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_588),
.B(n_533),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_666),
.B(n_220),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_703),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_633),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_707),
.B(n_538),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_713),
.B(n_533),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_605),
.B(n_567),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_636),
.B(n_667),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_687),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_590),
.A2(n_330),
.B1(n_331),
.B2(n_382),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_607),
.A2(n_382),
.B1(n_350),
.B2(n_352),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_588),
.B(n_533),
.Y(n_826)
);

AO22x2_ASAP7_75t_L g827 ( 
.A1(n_606),
.A2(n_475),
.B1(n_262),
.B2(n_260),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_719),
.B(n_469),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_694),
.A2(n_686),
.B1(n_678),
.B2(n_689),
.C(n_607),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_656),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_683),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_607),
.A2(n_366),
.B1(n_367),
.B2(n_364),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_683),
.B(n_545),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_719),
.B(n_223),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_684),
.B(n_545),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_607),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_545),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_672),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_672),
.B(n_426),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_609),
.B(n_225),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_697),
.B(n_225),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_698),
.B(n_545),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_698),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_702),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_702),
.B(n_545),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_709),
.A2(n_548),
.B(n_552),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_704),
.B(n_511),
.Y(n_847)
);

BUFx6f_ASAP7_75t_SL g848 ( 
.A(n_579),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_704),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_R g850 ( 
.A(n_626),
.B(n_254),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_661),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_722),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_661),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_579),
.B(n_226),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_705),
.B(n_511),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_594),
.B(n_548),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_626),
.A2(n_362),
.B1(n_350),
.B2(n_352),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_708),
.B(n_226),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_688),
.B(n_709),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_708),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_583),
.B(n_346),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_598),
.Y(n_863)
);

BUFx6f_ASAP7_75t_SL g864 ( 
.A(n_584),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_596),
.B(n_511),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_629),
.B(n_228),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_648),
.B(n_228),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_594),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_583),
.A2(n_288),
.B1(n_286),
.B2(n_285),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_603),
.B(n_548),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_603),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_604),
.B(n_548),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_648),
.B(n_426),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_598),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_615),
.B(n_232),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_631),
.B(n_232),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_604),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_612),
.A2(n_313),
.B(n_336),
.C(n_358),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_583),
.A2(n_554),
.B1(n_552),
.B2(n_511),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_612),
.B(n_548),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_646),
.B(n_235),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_615),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_616),
.B(n_617),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_616),
.B(n_554),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_611),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_611),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_718),
.B(n_235),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_617),
.Y(n_888)
);

INVx5_ASAP7_75t_L g889 ( 
.A(n_615),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_720),
.A2(n_275),
.B1(n_266),
.B2(n_263),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_723),
.A2(n_293),
.B1(n_256),
.B2(n_276),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_615),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_613),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_843),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_838),
.A2(n_364),
.B1(n_392),
.B2(n_376),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_782),
.B(n_596),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_797),
.B(n_596),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_797),
.B(n_239),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_843),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_749),
.A2(n_736),
.B1(n_822),
.B2(n_743),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_884),
.B(n_619),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_782),
.B(n_736),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_831),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_844),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_788),
.B(n_619),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_849),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_733),
.B(n_729),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_742),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_798),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_734),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_853),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_740),
.B(n_621),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_840),
.A2(n_357),
.B(n_353),
.Y(n_913)
);

AO21x1_ASAP7_75t_L g914 ( 
.A1(n_867),
.A2(n_360),
.B(n_601),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_748),
.B(n_621),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_759),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_761),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_882),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_861),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_762),
.B(n_751),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_750),
.B(n_621),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_781),
.B(n_371),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_754),
.B(n_641),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_734),
.B(n_239),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_762),
.B(n_428),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_SL g926 ( 
.A(n_776),
.B(n_328),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_734),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_758),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_729),
.B(n_641),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_765),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_730),
.B(n_737),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_873),
.A2(n_554),
.B1(n_601),
.B2(n_650),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_767),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_818),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_SL g935 ( 
.A1(n_731),
.A2(n_371),
.B1(n_363),
.B2(n_366),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_873),
.A2(n_650),
.B1(n_552),
.B2(n_623),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_808),
.B(n_585),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_794),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_873),
.A2(n_552),
.B1(n_622),
.B2(n_620),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_770),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_774),
.Y(n_941)
);

AO22x1_ASAP7_75t_L g942 ( 
.A1(n_731),
.A2(n_357),
.B1(n_362),
.B2(n_367),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_828),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_823),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_728),
.B(n_641),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_760),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_793),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_795),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_762),
.B(n_836),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_804),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_813),
.B(n_685),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_814),
.B(n_685),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_823),
.B(n_428),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_794),
.B(n_328),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_764),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_794),
.B(n_338),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_882),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_817),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_L g959 ( 
.A(n_745),
.B(n_356),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_730),
.B(n_685),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_752),
.A2(n_691),
.B1(n_692),
.B2(n_701),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_882),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_803),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_SL g964 ( 
.A(n_732),
.B(n_392),
.C(n_376),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_737),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_892),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_769),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_747),
.B(n_691),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_786),
.A2(n_620),
.B1(n_622),
.B2(n_623),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_739),
.B(n_691),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_800),
.B(n_692),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_SL g972 ( 
.A(n_824),
.B(n_322),
.C(n_292),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_868),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_792),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_892),
.B(n_634),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_777),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_SL g977 ( 
.A1(n_779),
.A2(n_371),
.B1(n_378),
.B2(n_373),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_739),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_792),
.B(n_429),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_852),
.B(n_429),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_777),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_763),
.B(n_430),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_801),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_871),
.Y(n_984)
);

NOR2x2_ASAP7_75t_L g985 ( 
.A(n_816),
.B(n_575),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_775),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_SL g987 ( 
.A(n_858),
.B(n_338),
.C(n_339),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_778),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_744),
.B(n_692),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_780),
.B(n_701),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_744),
.B(n_701),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_834),
.B(n_339),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_757),
.B(n_714),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_768),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_745),
.A2(n_714),
.B1(n_637),
.B2(n_674),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_839),
.B(n_714),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_827),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_746),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_877),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_827),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_892),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_756),
.A2(n_634),
.B(n_637),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_862),
.B(n_639),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_888),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_738),
.B(n_639),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_883),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_812),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_811),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_883),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_741),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_850),
.B(n_343),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_SL g1012 ( 
.A(n_807),
.B(n_343),
.C(n_344),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_SL g1013 ( 
.A(n_807),
.B(n_344),
.C(n_361),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_841),
.B(n_634),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_820),
.B(n_640),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_812),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_819),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_869),
.B(n_361),
.Y(n_1018)
);

NAND2x1p5_ASAP7_75t_L g1019 ( 
.A(n_812),
.B(n_637),
.Y(n_1019)
);

AND2x2_ASAP7_75t_SL g1020 ( 
.A(n_789),
.B(n_674),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_753),
.B(n_430),
.Y(n_1021)
);

OR2x4_ASAP7_75t_L g1022 ( 
.A(n_860),
.B(n_432),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_766),
.B(n_674),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_745),
.B(n_640),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_784),
.B(n_829),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_864),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_783),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_809),
.B(n_642),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_821),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_745),
.B(n_651),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_864),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_812),
.B(n_642),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_791),
.A2(n_727),
.B1(n_725),
.B2(n_724),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_811),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_859),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_735),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_796),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_741),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_809),
.B(n_642),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_830),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_851),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_799),
.Y(n_1042)
);

NAND2xp33_ASAP7_75t_L g1043 ( 
.A(n_787),
.B(n_356),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_854),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_863),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_874),
.B(n_651),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_885),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_886),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_846),
.A2(n_727),
.B(n_725),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_893),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_815),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_773),
.B(n_642),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_802),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_866),
.B(n_654),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_815),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_826),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_826),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_855),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_847),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_SL g1060 ( 
.A(n_825),
.B(n_389),
.C(n_369),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_889),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_856),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_833),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_785),
.B(n_642),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_825),
.A2(n_832),
.B(n_810),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_835),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_837),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_876),
.B(n_654),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_806),
.B(n_832),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_875),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_842),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_845),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_890),
.B(n_369),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_865),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_857),
.A2(n_663),
.B(n_657),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_755),
.B(n_432),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_657),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_771),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_887),
.B(n_663),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_884),
.B(n_649),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_857),
.B(n_649),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1021),
.B(n_433),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1006),
.A2(n_872),
.B1(n_870),
.B2(n_880),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_918),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1041),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_928),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_944),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_930),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_998),
.B(n_776),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_933),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1007),
.A2(n_889),
.B(n_790),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_963),
.B(n_891),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_1069),
.B(n_848),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_941),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1009),
.B(n_870),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_963),
.B(n_998),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_947),
.Y(n_1097)
);

AO32x1_ASAP7_75t_L g1098 ( 
.A1(n_1008),
.A2(n_433),
.A3(n_435),
.B1(n_462),
.B2(n_419),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_965),
.B(n_872),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1029),
.B(n_848),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_918),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_948),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_SL g1103 ( 
.A1(n_932),
.A2(n_880),
.B(n_879),
.Y(n_1103)
);

OR2x6_ASAP7_75t_SL g1104 ( 
.A(n_953),
.B(n_935),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1007),
.A2(n_889),
.B(n_649),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1065),
.A2(n_805),
.B(n_878),
.C(n_772),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1007),
.A2(n_889),
.B(n_669),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_965),
.B(n_547),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_978),
.B(n_547),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_978),
.B(n_553),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1007),
.A2(n_669),
.B(n_649),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_897),
.B(n_553),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1041),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_898),
.A2(n_573),
.B(n_576),
.C(n_569),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1053),
.B(n_373),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_897),
.B(n_560),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_916),
.B(n_418),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_981),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_938),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_913),
.A2(n_935),
.B(n_977),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_950),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1020),
.B(n_378),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_944),
.B(n_379),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1061),
.A2(n_669),
.B(n_649),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1061),
.A2(n_669),
.B(n_716),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_958),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1061),
.A2(n_669),
.B(n_716),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_SL g1128 ( 
.A(n_976),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1025),
.A2(n_724),
.B(n_721),
.C(n_717),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_940),
.B(n_560),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1020),
.B(n_379),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_917),
.B(n_388),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_1014),
.A2(n_618),
.B(n_625),
.C(n_613),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1025),
.A2(n_561),
.B1(n_573),
.B2(n_569),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_903),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_974),
.B(n_388),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_934),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_974),
.B(n_389),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_943),
.B(n_418),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1061),
.A2(n_716),
.B(n_717),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_908),
.B(n_716),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_994),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_909),
.B(n_716),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_905),
.A2(n_1005),
.B(n_931),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1049),
.A2(n_721),
.B(n_711),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_918),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_902),
.B(n_1056),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_SL g1148 ( 
.A(n_964),
.B(n_279),
.C(n_280),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1057),
.B(n_665),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1060),
.A2(n_576),
.B(n_564),
.C(n_561),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_943),
.Y(n_1151)
);

OAI21xp33_ASAP7_75t_SL g1152 ( 
.A1(n_932),
.A2(n_711),
.B(n_680),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1081),
.A2(n_680),
.B(n_679),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_996),
.B(n_281),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_SL g1155 ( 
.A1(n_992),
.A2(n_419),
.B(n_566),
.C(n_516),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_936),
.A2(n_575),
.B1(n_283),
.B2(n_327),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_949),
.B(n_665),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1080),
.A2(n_939),
.B(n_936),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_996),
.B(n_668),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_973),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_946),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_939),
.A2(n_679),
.B(n_670),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_982),
.B(n_668),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_984),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_900),
.B(n_937),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_979),
.B(n_295),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1000),
.A2(n_575),
.B1(n_300),
.B2(n_326),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1035),
.A2(n_303),
.B1(n_306),
.B2(n_311),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_955),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_982),
.B(n_670),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_909),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_1026),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1000),
.A2(n_394),
.B1(n_314),
.B2(n_618),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1036),
.B(n_0),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_990),
.A2(n_968),
.B(n_971),
.C(n_1036),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_926),
.B(n_195),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1014),
.A2(n_628),
.B(n_625),
.C(n_566),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1002),
.A2(n_628),
.B(n_566),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_931),
.A2(n_516),
.B(n_566),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_914),
.A2(n_990),
.B(n_1023),
.C(n_1018),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_968),
.A2(n_971),
.B(n_1042),
.C(n_945),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_999),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_918),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_967),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_977),
.A2(n_566),
.B1(n_516),
.B2(n_3),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1026),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_896),
.A2(n_566),
.B(n_516),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1051),
.B(n_511),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_938),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1003),
.A2(n_516),
.B1(n_2),
.B2(n_5),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1019),
.A2(n_516),
.B(n_511),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_957),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_907),
.A2(n_1073),
.B(n_1011),
.C(n_924),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1019),
.A2(n_511),
.B(n_191),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_983),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_957),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1070),
.A2(n_511),
.B1(n_190),
.B2(n_184),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_997),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_945),
.A2(n_12),
.A3(n_15),
.B(n_16),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1058),
.B(n_12),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1004),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_993),
.A2(n_177),
.B(n_174),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_960),
.A2(n_169),
.B(n_166),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_949),
.B(n_105),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_979),
.B(n_15),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1034),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_957),
.Y(n_1207)
);

INVx8_ASAP7_75t_L g1208 ( 
.A(n_949),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_904),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1055),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_906),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_SL g1212 ( 
.A(n_1016),
.B(n_25),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_911),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_970),
.A2(n_991),
.B(n_989),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_910),
.B(n_162),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1022),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_919),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1078),
.B(n_26),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_1031),
.B(n_124),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1017),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_986),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_907),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_980),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_988),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1078),
.B(n_37),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1028),
.A2(n_123),
.B(n_120),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1028),
.A2(n_111),
.B(n_107),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1063),
.B(n_103),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1022),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1037),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1027),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1040),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1054),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1076),
.B(n_41),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1076),
.B(n_47),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1076),
.A2(n_88),
.B1(n_85),
.B2(n_67),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_922),
.B(n_980),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1086),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1165),
.A2(n_1075),
.B(n_1024),
.Y(n_1239)
);

NAND3x1_ASAP7_75t_L g1240 ( 
.A(n_1234),
.B(n_927),
.C(n_972),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1088),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1101),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1207),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1151),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_SL g1245 ( 
.A(n_1147),
.B(n_957),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1118),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1181),
.A2(n_1015),
.B(n_929),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1147),
.B(n_1066),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1145),
.A2(n_1178),
.B(n_1153),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1095),
.B(n_1067),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1090),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1094),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1175),
.A2(n_929),
.B(n_969),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1095),
.B(n_1072),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1158),
.A2(n_1023),
.A3(n_1030),
.B(n_1079),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1099),
.B(n_1074),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1214),
.A2(n_1077),
.B(n_1068),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1179),
.A2(n_1052),
.B(n_1064),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1187),
.A2(n_1162),
.B(n_1155),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1216),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1082),
.B(n_895),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1097),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_R g1263 ( 
.A(n_1137),
.B(n_927),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1112),
.B(n_1116),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1103),
.A2(n_1039),
.B(n_1064),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1083),
.B(n_1059),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_SL g1267 ( 
.A(n_1142),
.B(n_962),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1223),
.B(n_920),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1102),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1177),
.A2(n_969),
.B(n_952),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1195),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1171),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1180),
.A2(n_1039),
.B(n_1052),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1120),
.A2(n_956),
.B1(n_954),
.B2(n_1062),
.Y(n_1274)
);

INVx3_ASAP7_75t_SL g1275 ( 
.A(n_1172),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1129),
.A2(n_921),
.B(n_951),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1083),
.B(n_1071),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1229),
.B(n_920),
.Y(n_1279)
);

NOR4xp25_ASAP7_75t_L g1280 ( 
.A(n_1198),
.B(n_959),
.C(n_1043),
.D(n_1013),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1140),
.A2(n_923),
.B(n_915),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1144),
.A2(n_975),
.B(n_1016),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1101),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1108),
.B(n_1050),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1126),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1193),
.A2(n_1106),
.B(n_1237),
.C(n_1092),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1134),
.A2(n_912),
.A3(n_1046),
.B(n_899),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1160),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1152),
.A2(n_1033),
.B(n_901),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1101),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1104),
.A2(n_1012),
.B1(n_1013),
.B2(n_925),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1207),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1115),
.B(n_942),
.Y(n_1293)
);

AOI221x1_ASAP7_75t_L g1294 ( 
.A1(n_1185),
.A2(n_894),
.B1(n_1047),
.B2(n_1044),
.C(n_1038),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_SL g1295 ( 
.A1(n_1233),
.A2(n_1001),
.B(n_1038),
.C(n_1010),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_925),
.B1(n_972),
.B2(n_987),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1182),
.Y(n_1297)
);

O2A1O1Ixp5_ASAP7_75t_L g1298 ( 
.A1(n_1122),
.A2(n_1010),
.B(n_1001),
.C(n_1048),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1144),
.A2(n_975),
.B(n_1016),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1091),
.A2(n_961),
.B(n_1032),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1183),
.Y(n_1301)
);

OAI22x1_ASAP7_75t_L g1302 ( 
.A1(n_1235),
.A2(n_985),
.B1(n_987),
.B2(n_925),
.Y(n_1302)
);

AO22x2_ASAP7_75t_L g1303 ( 
.A1(n_1185),
.A2(n_1198),
.B1(n_1206),
.B2(n_1233),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1186),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1174),
.A2(n_920),
.B(n_1045),
.C(n_1032),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1228),
.A2(n_995),
.B(n_901),
.Y(n_1306)
);

AOI221xp5_ASAP7_75t_L g1307 ( 
.A1(n_1206),
.A2(n_1210),
.B1(n_1190),
.B2(n_1200),
.C(n_1222),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1228),
.A2(n_966),
.B(n_962),
.C(n_1016),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_SL g1309 ( 
.A1(n_1226),
.A2(n_901),
.B(n_966),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1123),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1201),
.A2(n_966),
.B1(n_901),
.B2(n_54),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1109),
.B(n_51),
.Y(n_1312)
);

AOI221x1_ASAP7_75t_L g1313 ( 
.A1(n_1190),
.A2(n_52),
.B1(n_58),
.B2(n_61),
.C(n_1093),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1183),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1133),
.A2(n_58),
.B(n_1149),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1149),
.A2(n_1159),
.B(n_1170),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1096),
.A2(n_1220),
.B(n_1131),
.C(n_1210),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1111),
.A2(n_1124),
.B(n_1125),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1110),
.B(n_1163),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1209),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1211),
.A2(n_1217),
.B1(n_1213),
.B2(n_1230),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1105),
.A2(n_1107),
.B(n_1127),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1218),
.A2(n_1225),
.B(n_1114),
.C(n_1148),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1134),
.B(n_1135),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1227),
.A2(n_1150),
.B(n_1141),
.C(n_1202),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1208),
.Y(n_1326)
);

AOI221x1_ASAP7_75t_L g1327 ( 
.A1(n_1167),
.A2(n_1173),
.B1(n_1203),
.B2(n_1156),
.C(n_1194),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_SL g1329 ( 
.A(n_1168),
.B(n_1176),
.C(n_1236),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1154),
.A2(n_1188),
.B(n_1143),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1191),
.A2(n_1188),
.B(n_1232),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1192),
.Y(n_1332)
);

OAI22x1_ASAP7_75t_L g1333 ( 
.A1(n_1204),
.A2(n_1089),
.B1(n_1136),
.B2(n_1100),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1156),
.A2(n_1173),
.B(n_1167),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1130),
.B(n_1166),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1084),
.A2(n_1146),
.B(n_1215),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1161),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1208),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1197),
.A2(n_1184),
.B(n_1224),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1139),
.B(n_1117),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1084),
.A2(n_1146),
.B(n_1221),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1169),
.B(n_1231),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1085),
.B(n_1113),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1098),
.A2(n_1157),
.B(n_1219),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1205),
.A2(n_1098),
.B(n_1208),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1098),
.A2(n_1157),
.B(n_1212),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1119),
.A2(n_1189),
.B(n_1196),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1196),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1199),
.B(n_1128),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1128),
.A2(n_732),
.B(n_802),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1199),
.A2(n_932),
.B(n_1025),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1199),
.B(n_742),
.Y(n_1352)
);

INVx6_ASAP7_75t_SL g1353 ( 
.A(n_1204),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_SL g1354 ( 
.A1(n_1147),
.A2(n_1193),
.B(n_1228),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1120),
.A2(n_1025),
.B(n_1065),
.C(n_1193),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1086),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1158),
.A2(n_1103),
.B(n_1214),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1214),
.A2(n_1061),
.B(n_1007),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1237),
.A2(n_732),
.B1(n_753),
.B2(n_746),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1118),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1086),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1237),
.B(n_732),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1237),
.B(n_732),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1181),
.A2(n_1025),
.B(n_1175),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1145),
.A2(n_1178),
.B(n_1153),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1237),
.A2(n_732),
.B1(n_753),
.B2(n_746),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1181),
.A2(n_1175),
.B(n_1165),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1207),
.B(n_938),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1237),
.B(n_1053),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1082),
.B(n_599),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1375)
);

AOI221x1_ASAP7_75t_L g1376 ( 
.A1(n_1120),
.A2(n_1185),
.B1(n_1065),
.B2(n_1190),
.C(n_1175),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1087),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1207),
.B(n_938),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1177),
.A2(n_1181),
.B(n_1180),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1237),
.B(n_1053),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1147),
.B(n_1006),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1120),
.B(n_732),
.C(n_581),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1095),
.A2(n_797),
.B1(n_1009),
.B2(n_1006),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1086),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1082),
.B(n_742),
.Y(n_1386)
);

AOI221x1_ASAP7_75t_L g1387 ( 
.A1(n_1120),
.A2(n_1185),
.B1(n_1065),
.B2(n_1190),
.C(n_1175),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_SL g1388 ( 
.A1(n_1175),
.A2(n_1181),
.B(n_1165),
.C(n_1228),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1120),
.A2(n_728),
.B(n_822),
.C(n_581),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1145),
.A2(n_1178),
.B(n_1153),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1334),
.A2(n_1367),
.B(n_1357),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1318),
.A2(n_1258),
.B(n_1322),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1340),
.B(n_1386),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1257),
.A2(n_1388),
.B(n_1357),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_1326),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1334),
.A2(n_1367),
.B(n_1289),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1238),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1263),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1331),
.A2(n_1281),
.B(n_1300),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1241),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1354),
.A2(n_1245),
.B(n_1317),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1389),
.A2(n_1355),
.B(n_1383),
.C(n_1351),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1310),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1246),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1251),
.B(n_1269),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1358),
.A2(n_1364),
.B(n_1363),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1293),
.A2(n_1286),
.B(n_1323),
.C(n_1350),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1307),
.A2(n_1375),
.B(n_1358),
.C(n_1382),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1288),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1259),
.A2(n_1282),
.B(n_1299),
.Y(n_1412)
);

INVx4_ASAP7_75t_SL g1413 ( 
.A(n_1283),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1244),
.B(n_1312),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1273),
.A2(n_1359),
.B(n_1309),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1374),
.B(n_1375),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1356),
.B(n_1362),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1294),
.A2(n_1387),
.B(n_1376),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_SL g1420 ( 
.A(n_1361),
.B(n_1271),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1239),
.A2(n_1341),
.B(n_1265),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1305),
.B(n_1333),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1247),
.A2(n_1330),
.B(n_1316),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1252),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1247),
.A2(n_1346),
.B(n_1253),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1262),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1283),
.Y(n_1428)
);

AOI221x1_ASAP7_75t_L g1429 ( 
.A1(n_1303),
.A2(n_1311),
.B1(n_1291),
.B2(n_1349),
.C(n_1315),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1276),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1327),
.A2(n_1253),
.B(n_1266),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1307),
.A2(n_1291),
.B1(n_1296),
.B2(n_1302),
.C(n_1311),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1266),
.A2(n_1278),
.B(n_1325),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1285),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1278),
.A2(n_1308),
.B(n_1313),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1297),
.Y(n_1436)
);

AO32x2_ASAP7_75t_L g1437 ( 
.A1(n_1384),
.A2(n_1296),
.A3(n_1321),
.B1(n_1303),
.B2(n_1295),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1377),
.B(n_1382),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1320),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1316),
.A2(n_1380),
.B(n_1306),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1349),
.A2(n_1324),
.B(n_1298),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1380),
.A2(n_1306),
.B(n_1345),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1336),
.A2(n_1277),
.B(n_1270),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1277),
.A2(n_1270),
.B(n_1324),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1360),
.A2(n_1369),
.B(n_1264),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1385),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1370),
.A2(n_1264),
.B(n_1280),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1321),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1344),
.A2(n_1384),
.B(n_1256),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1344),
.A2(n_1256),
.B(n_1250),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1248),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1250),
.A2(n_1254),
.B(n_1248),
.Y(n_1452)
);

NAND2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1267),
.B(n_1243),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1244),
.B(n_1312),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1279),
.B(n_1337),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1254),
.A2(n_1284),
.B(n_1319),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1243),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1329),
.A2(n_1328),
.B1(n_1370),
.B2(n_1261),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1319),
.B(n_1284),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1372),
.A2(n_1381),
.B1(n_1335),
.B2(n_1240),
.Y(n_1460)
);

AOI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1274),
.A2(n_1339),
.B(n_1268),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1342),
.A2(n_1343),
.B(n_1287),
.Y(n_1462)
);

NAND2x1p5_ASAP7_75t_L g1463 ( 
.A(n_1292),
.B(n_1242),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1378),
.A2(n_1279),
.B1(n_1304),
.B2(n_1343),
.C(n_1275),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1348),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1292),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1283),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1379),
.A2(n_1371),
.B(n_1347),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1353),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1255),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1255),
.A2(n_1287),
.B(n_1242),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1301),
.B(n_1332),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1290),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1290),
.B(n_1314),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1287),
.A2(n_1332),
.B(n_1314),
.Y(n_1475)
);

INVx8_ASAP7_75t_L g1476 ( 
.A(n_1290),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1353),
.B(n_1314),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1340),
.B(n_1365),
.Y(n_1478)
);

OAI21xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1334),
.A2(n_1363),
.B(n_1358),
.Y(n_1479)
);

BUFx5_ASAP7_75t_L g1480 ( 
.A(n_1352),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1357),
.A2(n_1294),
.B(n_1367),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1249),
.A2(n_1178),
.B(n_1368),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1370),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1383),
.B(n_732),
.C(n_1389),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1272),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1383),
.A2(n_1120),
.B1(n_1303),
.B2(n_1307),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1357),
.A2(n_1294),
.B(n_1367),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1260),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1294),
.A2(n_1357),
.A3(n_1376),
.B(n_1387),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1305),
.B(n_1333),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1238),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1357),
.A2(n_1294),
.B(n_1367),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1383),
.A2(n_1120),
.B1(n_1303),
.B2(n_1307),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1338),
.B(n_1326),
.Y(n_1495)
);

AO31x2_ASAP7_75t_L g1496 ( 
.A1(n_1294),
.A2(n_1357),
.A3(n_1376),
.B(n_1387),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1389),
.A2(n_1120),
.B1(n_1383),
.B2(n_1307),
.C(n_731),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1238),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1383),
.A2(n_1310),
.B1(n_732),
.B2(n_1365),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1389),
.A2(n_1334),
.B(n_1355),
.C(n_1120),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1260),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1354),
.A2(n_1245),
.B(n_1334),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1338),
.B(n_1326),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1238),
.Y(n_1505)
);

INVx4_ASAP7_75t_SL g1506 ( 
.A(n_1283),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1507)
);

BUFx8_ASAP7_75t_L g1508 ( 
.A(n_1246),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1340),
.B(n_1386),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1357),
.A2(n_1294),
.B(n_1367),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1238),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1249),
.A2(n_1178),
.B(n_1368),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1340),
.B(n_1386),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1383),
.A2(n_1389),
.B(n_581),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1249),
.A2(n_1178),
.B(n_1368),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1383),
.B(n_1365),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1238),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1238),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1249),
.A2(n_1390),
.B(n_1368),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1272),
.Y(n_1522)
);

AO21x1_ASAP7_75t_L g1523 ( 
.A1(n_1334),
.A2(n_1389),
.B(n_1311),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1238),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1383),
.A2(n_1120),
.B1(n_1303),
.B2(n_1307),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1357),
.A2(n_1294),
.B(n_1367),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1249),
.A2(n_1178),
.B(n_1368),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1389),
.A2(n_1120),
.B1(n_1383),
.B2(n_1307),
.C(n_731),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1383),
.A2(n_1389),
.B(n_581),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1272),
.Y(n_1530)
);

O2A1O1Ixp5_ASAP7_75t_L g1531 ( 
.A1(n_1334),
.A2(n_1367),
.B(n_1357),
.C(n_1355),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1243),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1365),
.A2(n_732),
.B1(n_1366),
.B2(n_1383),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1305),
.B(n_1333),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1238),
.Y(n_1535)
);

AOI22x1_ASAP7_75t_L g1536 ( 
.A1(n_1334),
.A2(n_1333),
.B1(n_1354),
.B2(n_1303),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1389),
.A2(n_1383),
.B(n_1355),
.C(n_1334),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1533),
.A2(n_1411),
.B1(n_1460),
.B2(n_1458),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1458),
.A2(n_1518),
.B1(n_1493),
.B2(n_1525),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1518),
.A2(n_1500),
.B1(n_1528),
.B2(n_1497),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1394),
.B(n_1509),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1478),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1445),
.A2(n_1484),
.B1(n_1523),
.B2(n_1525),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1501),
.A2(n_1409),
.B(n_1514),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1486),
.A2(n_1493),
.B1(n_1501),
.B2(n_1404),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1459),
.B(n_1416),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1406),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1430),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1486),
.A2(n_1464),
.B1(n_1408),
.B2(n_1425),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1417),
.B(n_1438),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1399),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1403),
.A2(n_1409),
.B1(n_1414),
.B2(n_1454),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1529),
.A2(n_1537),
.B(n_1407),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1455),
.B(n_1418),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1430),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1556)
);

AOI211xp5_ASAP7_75t_L g1557 ( 
.A1(n_1403),
.A2(n_1432),
.B(n_1479),
.C(n_1461),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1508),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1485),
.B(n_1522),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1440),
.A2(n_1442),
.B(n_1429),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1434),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1410),
.B(n_1491),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1531),
.A2(n_1391),
.B(n_1397),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1436),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1491),
.B(n_1498),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1439),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1433),
.A2(n_1453),
.B(n_1397),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1498),
.B(n_1505),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1531),
.A2(n_1503),
.B(n_1402),
.C(n_1534),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1442),
.A2(n_1426),
.B(n_1443),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1422),
.A2(n_1490),
.B1(n_1534),
.B2(n_1536),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1422),
.B(n_1490),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1485),
.B(n_1522),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1398),
.B(n_1401),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1488),
.A2(n_1502),
.B1(n_1530),
.B2(n_1399),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1424),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1511),
.B(n_1519),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1520),
.B(n_1524),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1427),
.B(n_1446),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1441),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1396),
.A2(n_1504),
.B(n_1495),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1481),
.A2(n_1510),
.B(n_1526),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1405),
.A2(n_1469),
.B1(n_1477),
.B2(n_1396),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1535),
.B(n_1465),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1481),
.A2(n_1492),
.B(n_1487),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1423),
.A2(n_1475),
.B(n_1449),
.C(n_1450),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1457),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1473),
.B(n_1480),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1480),
.B(n_1462),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1480),
.B(n_1472),
.Y(n_1591)
);

BUFx12f_ASAP7_75t_L g1592 ( 
.A(n_1508),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1413),
.B(n_1506),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1457),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1456),
.B(n_1480),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1474),
.A2(n_1419),
.B(n_1431),
.C(n_1435),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1449),
.A2(n_1450),
.B(n_1468),
.C(n_1419),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1480),
.B(n_1532),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1467),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1466),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1469),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1467),
.B(n_1463),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1435),
.A2(n_1431),
.B1(n_1428),
.B2(n_1487),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1444),
.A2(n_1412),
.B(n_1415),
.Y(n_1604)
);

AOI211xp5_ASAP7_75t_L g1605 ( 
.A1(n_1420),
.A2(n_1415),
.B(n_1468),
.C(n_1421),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1437),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1489),
.B(n_1496),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_SL g1608 ( 
.A1(n_1489),
.A2(n_1496),
.B(n_1492),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1496),
.B(n_1510),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1470),
.A2(n_1405),
.B(n_1506),
.C(n_1413),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1428),
.B(n_1476),
.Y(n_1611)
);

O2A1O1Ixp5_ASAP7_75t_L g1612 ( 
.A1(n_1412),
.A2(n_1400),
.B(n_1393),
.C(n_1527),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1428),
.A2(n_1476),
.B1(n_1482),
.B2(n_1515),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1392),
.B(n_1494),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1494),
.Y(n_1615)
);

O2A1O1Ixp5_ASAP7_75t_L g1616 ( 
.A1(n_1512),
.A2(n_1499),
.B(n_1507),
.C(n_1516),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1499),
.B(n_1507),
.Y(n_1617)
);

O2A1O1Ixp5_ASAP7_75t_L g1618 ( 
.A1(n_1517),
.A2(n_1523),
.B(n_1334),
.C(n_1531),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1521),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1521),
.B(n_1414),
.Y(n_1620)
);

A2O1A1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1531),
.A2(n_1501),
.B(n_1334),
.C(n_1389),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1394),
.B(n_1509),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_SL g1623 ( 
.A(n_1422),
.B(n_1490),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1483),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1531),
.A2(n_1501),
.B(n_1334),
.C(n_1389),
.Y(n_1625)
);

BUFx4f_ASAP7_75t_SL g1626 ( 
.A(n_1405),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1394),
.B(n_1509),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1518),
.B(n_1459),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1394),
.B(n_1509),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1508),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1394),
.B(n_1509),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1483),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1483),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1440),
.A2(n_1395),
.B(n_1471),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1394),
.B(n_1509),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1485),
.B(n_1522),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1411),
.A2(n_935),
.B1(n_977),
.B2(n_1533),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1414),
.B(n_1454),
.Y(n_1638)
);

O2A1O1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1500),
.A2(n_1408),
.B(n_1389),
.C(n_1355),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1501),
.A2(n_1286),
.B(n_1355),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1579),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1620),
.B(n_1591),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1548),
.B(n_1564),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1559),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1576),
.B(n_1586),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1556),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1555),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1597),
.A2(n_1585),
.B(n_1582),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1595),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1561),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1566),
.Y(n_1652)
);

OAI332xp33_ASAP7_75t_L g1653 ( 
.A1(n_1637),
.A2(n_1538),
.A3(n_1539),
.B1(n_1549),
.B2(n_1545),
.B3(n_1552),
.C1(n_1628),
.C2(n_1571),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1567),
.B(n_1553),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1587),
.A2(n_1563),
.B(n_1625),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1590),
.B(n_1607),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1550),
.B(n_1546),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1638),
.B(n_1540),
.Y(n_1658)
);

AO31x2_ASAP7_75t_L g1659 ( 
.A1(n_1603),
.A2(n_1587),
.A3(n_1621),
.B(n_1625),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1542),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1632),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1559),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1633),
.B(n_1609),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1572),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1580),
.B(n_1606),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1580),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_R g1667 ( 
.A(n_1551),
.B(n_1593),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1581),
.B(n_1572),
.Y(n_1668)
);

AO31x2_ASAP7_75t_L g1669 ( 
.A1(n_1615),
.A2(n_1619),
.A3(n_1623),
.B(n_1613),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1547),
.B(n_1572),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1573),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1570),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1612),
.A2(n_1616),
.B(n_1608),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1604),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1596),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1618),
.A2(n_1543),
.B(n_1617),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1560),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1604),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1562),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1573),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1565),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1568),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1639),
.B(n_1554),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1557),
.B(n_1584),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1574),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1577),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1544),
.B(n_1578),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1569),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1653),
.A2(n_1640),
.B1(n_1630),
.B2(n_1558),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1672),
.Y(n_1690)
);

OAI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1684),
.A2(n_1575),
.B1(n_1610),
.B2(n_1630),
.C1(n_1631),
.C2(n_1635),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1672),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1668),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1643),
.B(n_1634),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1666),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1651),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1648),
.B(n_1605),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1666),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1656),
.B(n_1636),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1654),
.B(n_1668),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1657),
.A2(n_1683),
.B1(n_1658),
.B2(n_1654),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1648),
.B(n_1541),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1688),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1665),
.B(n_1636),
.Y(n_1705)
);

NAND2x1_ASAP7_75t_L g1706 ( 
.A(n_1654),
.B(n_1593),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1665),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1648),
.B(n_1629),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1663),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1647),
.B(n_1627),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1655),
.B(n_1622),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1669),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_1600),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1655),
.B(n_1588),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1675),
.B(n_1599),
.Y(n_1716)
);

INVx3_ASAP7_75t_SL g1717 ( 
.A(n_1654),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1644),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1687),
.B(n_1594),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1644),
.B(n_1602),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1663),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1644),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1689),
.A2(n_1654),
.B1(n_1668),
.B2(n_1664),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_1702),
.C(n_1688),
.D(n_1704),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1707),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1705),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1694),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1702),
.A2(n_1664),
.B1(n_1668),
.B2(n_1670),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1709),
.Y(n_1730)
);

INVxp67_ASAP7_75t_SL g1731 ( 
.A(n_1704),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1691),
.A2(n_1675),
.B1(n_1660),
.B2(n_1685),
.C(n_1686),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1709),
.B(n_1661),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1690),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1711),
.A2(n_1677),
.B1(n_1686),
.B2(n_1685),
.C(n_1647),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1696),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1641),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1710),
.B(n_1641),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1694),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1711),
.B(n_1642),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1700),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1694),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1719),
.A2(n_1701),
.B(n_1706),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1719),
.A2(n_1667),
.B1(n_1671),
.B2(n_1662),
.C(n_1583),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1721),
.B(n_1661),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1711),
.B(n_1670),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1716),
.B(n_1646),
.C(n_1679),
.D(n_1681),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1718),
.B(n_1642),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1718),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1713),
.B(n_1650),
.C(n_1676),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1691),
.A2(n_1698),
.B1(n_1712),
.B2(n_1716),
.C(n_1713),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1697),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1701),
.A2(n_1601),
.B1(n_1680),
.B2(n_1676),
.C(n_1645),
.Y(n_1753)
);

OAI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1701),
.A2(n_1676),
.B(n_1677),
.C(n_1652),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1696),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1703),
.B(n_1708),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1722),
.B(n_1642),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1716),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_L g1759 ( 
.A(n_1713),
.B(n_1650),
.C(n_1679),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1721),
.B(n_1659),
.Y(n_1761)
);

NAND3xp33_ASAP7_75t_L g1762 ( 
.A(n_1715),
.B(n_1650),
.C(n_1682),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1725),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1743),
.B(n_1717),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1727),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1739),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1751),
.B(n_1698),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1734),
.Y(n_1768)
);

AND2x4_ASAP7_75t_SL g1769 ( 
.A(n_1740),
.B(n_1698),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1742),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1750),
.B(n_1706),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1754),
.A2(n_1712),
.B(n_1673),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1760),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1731),
.B(n_1699),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1732),
.B(n_1693),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1746),
.B(n_1695),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1736),
.B(n_1695),
.Y(n_1777)
);

INVx4_ASAP7_75t_SL g1778 ( 
.A(n_1758),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1758),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1759),
.A2(n_1674),
.B(n_1678),
.Y(n_1781)
);

INVxp67_ASAP7_75t_SL g1782 ( 
.A(n_1761),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1755),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1724),
.B(n_1650),
.C(n_1715),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1725),
.Y(n_1785)
);

AOI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1749),
.A2(n_1714),
.B(n_1692),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1728),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1723),
.B(n_1715),
.C(n_1649),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1728),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1786),
.Y(n_1790)
);

INVx5_ASAP7_75t_L g1791 ( 
.A(n_1771),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1763),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1786),
.Y(n_1793)
);

AND2x2_ASAP7_75t_SL g1794 ( 
.A(n_1787),
.B(n_1729),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1786),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1767),
.B(n_1733),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1769),
.B(n_1748),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1765),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1730),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1784),
.B(n_1744),
.C(n_1735),
.D(n_1753),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1783),
.B(n_1737),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1778),
.B(n_1693),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1765),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1782),
.B(n_1738),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1787),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1766),
.Y(n_1806)
);

INVx4_ASAP7_75t_L g1807 ( 
.A(n_1778),
.Y(n_1807)
);

AND2x4_ASAP7_75t_SL g1808 ( 
.A(n_1763),
.B(n_1757),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1766),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1776),
.B(n_1778),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1770),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1785),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1782),
.B(n_1733),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1787),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1776),
.B(n_1726),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1770),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1778),
.B(n_1726),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1778),
.B(n_1741),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1767),
.B(n_1745),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1779),
.B(n_1756),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1777),
.B(n_1747),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1779),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1778),
.B(n_1693),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1789),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1774),
.B(n_1762),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1781),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1781),
.Y(n_1827)
);

NOR2x1p5_ASAP7_75t_SL g1828 ( 
.A(n_1805),
.B(n_1768),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1792),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1810),
.B(n_1764),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1792),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1812),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1812),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1798),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1798),
.Y(n_1835)
);

INVx3_ASAP7_75t_SL g1836 ( 
.A(n_1807),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1796),
.B(n_1775),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1810),
.B(n_1780),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1794),
.B(n_1775),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1810),
.B(n_1797),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1794),
.B(n_1780),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1803),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1805),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1800),
.B(n_1764),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1807),
.B(n_1773),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1807),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1805),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1800),
.B(n_1626),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1796),
.B(n_1784),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1807),
.B(n_1789),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1803),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1794),
.B(n_1780),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1801),
.B(n_1708),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1797),
.B(n_1773),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1806),
.Y(n_1855)
);

NAND2x1_ASAP7_75t_L g1856 ( 
.A(n_1824),
.B(n_1802),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1791),
.B(n_1788),
.C(n_1772),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1819),
.B(n_1774),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1808),
.B(n_1789),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1806),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1809),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1814),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1819),
.B(n_1705),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1801),
.B(n_1708),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1821),
.B(n_1785),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1843),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1858),
.B(n_1821),
.Y(n_1867)
);

OAI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1839),
.A2(n_1788),
.B1(n_1791),
.B2(n_1771),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1843),
.Y(n_1869)
);

CKINVDCx16_ASAP7_75t_R g1870 ( 
.A(n_1848),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1862),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1865),
.B(n_1814),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1844),
.B(n_1820),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1848),
.B(n_1626),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1841),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1862),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1844),
.B(n_1802),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1859),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1829),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1859),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1859),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1831),
.B(n_1820),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1836),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1840),
.B(n_1808),
.Y(n_1884)
);

OAI21x1_ASAP7_75t_L g1885 ( 
.A1(n_1856),
.A2(n_1824),
.B(n_1814),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_L g1886 ( 
.A(n_1857),
.B(n_1824),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1832),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1838),
.B(n_1808),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1830),
.B(n_1802),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1830),
.B(n_1802),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1854),
.B(n_1823),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1823),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1886),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1866),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1886),
.A2(n_1837),
.B(n_1852),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1870),
.A2(n_1823),
.B1(n_1850),
.B2(n_1836),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1885),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1866),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1870),
.A2(n_1849),
.B1(n_1791),
.B2(n_1846),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1889),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1869),
.Y(n_1901)
);

O2A1O1Ixp5_ASAP7_75t_L g1902 ( 
.A1(n_1868),
.A2(n_1877),
.B(n_1873),
.C(n_1850),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1869),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1885),
.Y(n_1904)
);

OAI32xp33_ASAP7_75t_L g1905 ( 
.A1(n_1883),
.A2(n_1833),
.A3(n_1824),
.B1(n_1846),
.B2(n_1825),
.Y(n_1905)
);

AOI33xp33_ASAP7_75t_L g1906 ( 
.A1(n_1879),
.A2(n_1834),
.A3(n_1835),
.B1(n_1861),
.B2(n_1860),
.B3(n_1855),
.Y(n_1906)
);

O2A1O1Ixp5_ASAP7_75t_L g1907 ( 
.A1(n_1878),
.A2(n_1850),
.B(n_1846),
.C(n_1880),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1889),
.B(n_1845),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1890),
.A2(n_1823),
.B1(n_1818),
.B2(n_1817),
.Y(n_1909)
);

OAI32xp33_ASAP7_75t_L g1910 ( 
.A1(n_1875),
.A2(n_1825),
.A3(n_1847),
.B1(n_1842),
.B2(n_1851),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1871),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1878),
.B(n_1880),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1871),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1908),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1900),
.B(n_1878),
.Y(n_1915)
);

OAI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1902),
.A2(n_1872),
.B(n_1880),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1908),
.B(n_1881),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1912),
.B(n_1881),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1899),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1893),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1896),
.B(n_1881),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1909),
.B(n_1890),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1897),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1894),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1895),
.B(n_1892),
.Y(n_1925)
);

AOI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1916),
.A2(n_1910),
.B1(n_1905),
.B2(n_1907),
.C(n_1887),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1920),
.A2(n_1905),
.B(n_1910),
.C(n_1919),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1925),
.A2(n_1906),
.B1(n_1867),
.B2(n_1904),
.C(n_1872),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1915),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1917),
.Y(n_1930)
);

O2A1O1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1920),
.A2(n_1913),
.B(n_1911),
.C(n_1898),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1925),
.Y(n_1932)
);

AOI321xp33_ASAP7_75t_L g1933 ( 
.A1(n_1921),
.A2(n_1903),
.A3(n_1901),
.B1(n_1897),
.B2(n_1867),
.C(n_1879),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1914),
.A2(n_1918),
.B(n_1874),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1923),
.A2(n_1887),
.B(n_1876),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_SL g1936 ( 
.A(n_1922),
.B(n_1906),
.C(n_1876),
.Y(n_1936)
);

INVxp67_ASAP7_75t_SL g1937 ( 
.A(n_1932),
.Y(n_1937)
);

OAI221xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1926),
.A2(n_1933),
.B1(n_1927),
.B2(n_1922),
.C(n_1934),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1931),
.Y(n_1939)
);

AOI21xp33_ASAP7_75t_L g1940 ( 
.A1(n_1929),
.A2(n_1930),
.B(n_1924),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1936),
.A2(n_1892),
.B1(n_1891),
.B2(n_1888),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1928),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1935),
.A2(n_1791),
.B1(n_1882),
.B2(n_1891),
.Y(n_1943)
);

NOR4xp25_ASAP7_75t_SL g1944 ( 
.A(n_1928),
.B(n_1828),
.C(n_1847),
.D(n_1791),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1941),
.B(n_1937),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1939),
.B(n_1884),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1942),
.Y(n_1947)
);

AOI32xp33_ASAP7_75t_L g1948 ( 
.A1(n_1943),
.A2(n_1884),
.A3(n_1888),
.B1(n_1818),
.B2(n_1817),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1938),
.B(n_1592),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1940),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1943),
.B(n_1863),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1944),
.B(n_1864),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1947),
.A2(n_1791),
.B1(n_1771),
.B2(n_1815),
.Y(n_1953)
);

XNOR2xp5_ASAP7_75t_L g1954 ( 
.A(n_1946),
.B(n_1853),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1949),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1945),
.Y(n_1956)
);

AOI222xp33_ASAP7_75t_L g1957 ( 
.A1(n_1950),
.A2(n_1791),
.B1(n_1826),
.B2(n_1827),
.C1(n_1795),
.C2(n_1793),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1951),
.A2(n_1771),
.B1(n_1815),
.B2(n_1799),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1956),
.B(n_1952),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1954),
.B(n_1799),
.Y(n_1960)
);

NOR2xp67_ASAP7_75t_L g1961 ( 
.A(n_1955),
.B(n_1948),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1957),
.Y(n_1962)
);

NAND2x1p5_ASAP7_75t_L g1963 ( 
.A(n_1959),
.B(n_1958),
.Y(n_1963)
);

OAI211xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1963),
.A2(n_1962),
.B(n_1960),
.C(n_1961),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_L g1965 ( 
.A(n_1964),
.B(n_1795),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1964),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1965),
.Y(n_1967)
);

AO22x2_ASAP7_75t_L g1968 ( 
.A1(n_1966),
.A2(n_1827),
.B1(n_1826),
.B2(n_1793),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1967),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1968),
.A2(n_1953),
.B1(n_1813),
.B2(n_1804),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1969),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1971),
.A2(n_1970),
.B1(n_1827),
.B2(n_1826),
.Y(n_1972)
);

OA21x2_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1793),
.B(n_1790),
.Y(n_1973)
);

NOR3xp33_ASAP7_75t_SL g1974 ( 
.A(n_1973),
.B(n_1611),
.C(n_1804),
.Y(n_1974)
);

OA22x2_ASAP7_75t_L g1975 ( 
.A1(n_1974),
.A2(n_1795),
.B1(n_1790),
.B2(n_1822),
.Y(n_1975)
);

AOI211xp5_ASAP7_75t_L g1976 ( 
.A1(n_1975),
.A2(n_1816),
.B(n_1822),
.C(n_1811),
.Y(n_1976)
);


endmodule