module fake_netlist_6_1363_n_2726 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_808, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_788, n_325, n_767, n_804, n_329, n_464, n_600, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2726);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_788;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2726;

wire n_992;
wire n_2542;
wire n_1671;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_1371;
wire n_873;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_822;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_1344;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_1663;
wire n_2009;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_1165;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2319;
wire n_2519;
wire n_825;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_890;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_1992;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_931;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2289;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1818;
wire n_1108;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_1900;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_876;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_875;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_1461;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1362;
wire n_1156;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_798),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_167),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_574),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_296),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_311),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_272),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_724),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_766),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_255),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_396),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_785),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_264),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_775),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

CKINVDCx16_ASAP7_75t_R g827 ( 
.A(n_321),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_343),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_328),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_186),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_401),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_463),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_739),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_671),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_485),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_650),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_758),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_466),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_216),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_93),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_85),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_87),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_114),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_223),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_411),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_805),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_407),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_528),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_629),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_480),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_261),
.Y(n_851)
);

BUFx10_ASAP7_75t_L g852 ( 
.A(n_760),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_357),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_687),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_251),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_769),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_429),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_61),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_522),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_551),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_106),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_210),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_5),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_518),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_224),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_161),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_200),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_24),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_113),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_759),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_1),
.Y(n_872)
);

INVxp33_ASAP7_75t_R g873 ( 
.A(n_213),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_793),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_233),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_588),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_367),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_763),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_227),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_213),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_559),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_554),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_177),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_427),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_286),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_647),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_303),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_369),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_613),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_770),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_796),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_686),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_654),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_658),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_495),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_757),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_748),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_263),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_490),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_301),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_562),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_678),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_227),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_79),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_754),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_443),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_158),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_26),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_508),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_46),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_251),
.Y(n_911)
);

BUFx10_ASAP7_75t_L g912 ( 
.A(n_780),
.Y(n_912)
);

BUFx10_ASAP7_75t_L g913 ( 
.A(n_579),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_571),
.Y(n_914)
);

BUFx5_ASAP7_75t_L g915 ( 
.A(n_266),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_346),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_379),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_644),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_640),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_252),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_615),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_572),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_799),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_513),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_8),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_60),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_449),
.Y(n_927)
);

CKINVDCx16_ASAP7_75t_R g928 ( 
.A(n_550),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_433),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_20),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_637),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_215),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_68),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_774),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_66),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_33),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_381),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_54),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_704),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_117),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_139),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_595),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_232),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_27),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_717),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_85),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_468),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_437),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_432),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_290),
.Y(n_950)
);

BUFx10_ASAP7_75t_L g951 ( 
.A(n_106),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_289),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_736),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_777),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_601),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_781),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_576),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_49),
.Y(n_958)
);

INVx4_ASAP7_75t_R g959 ( 
.A(n_794),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_744),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_745),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_90),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_304),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_15),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_265),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_573),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_795),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_484),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_115),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_544),
.Y(n_970)
);

BUFx10_ASAP7_75t_L g971 ( 
.A(n_669),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_477),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_753),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_231),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_812),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_111),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_740),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_404),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_400),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_765),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_589),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_786),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_608),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_619),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_475),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_2),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_585),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_0),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_417),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_782),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_44),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_110),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_389),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_455),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_453),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_163),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_677),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_126),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_778),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_462),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_65),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_247),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_88),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_738),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_132),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_626),
.Y(n_1006)
);

CKINVDCx14_ASAP7_75t_R g1007 ( 
.A(n_170),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_750),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_72),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_764),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_147),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_234),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_402),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_768),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_423),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_742),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_313),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_259),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_60),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_783),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_190),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_309),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_646),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_497),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_534),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_561),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_241),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_182),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_167),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_747),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_483),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_552),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_268),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_465),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_302),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_132),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_351),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_521),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_342),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_165),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_298),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_482),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_174),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_209),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_776),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_674),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_788),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_121),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_335),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_743),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_388),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_121),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_577),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_233),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_703),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_741),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_772),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_71),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_692),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_272),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_706),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_133),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_752),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_761),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_390),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_42),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_751),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_101),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_633),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_376),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_119),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_811),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_3),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_69),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_789),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_632),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_300),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_299),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_605),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_101),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_3),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_266),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_496),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_385),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_116),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_284),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_446),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_697),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_802),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_306),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_749),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_755),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_420),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_458),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_73),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_12),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_163),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_89),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_787),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_806),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_212),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_5),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_801),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_394),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_569),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_504),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_347),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_269),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_331),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_218),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_240),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_171),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_290),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_96),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_242),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_364),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_76),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_612),
.Y(n_1118)
);

BUFx10_ASAP7_75t_L g1119 ( 
.A(n_157),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_702),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_474),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_606),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_767),
.Y(n_1123)
);

CKINVDCx14_ASAP7_75t_R g1124 ( 
.A(n_168),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_110),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_590),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_540),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_610),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_409),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_457),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_655),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_122),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_202),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_712),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_790),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_244),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_578),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_223),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_516),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_737),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_541),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_226),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_141),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_393),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_542),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_792),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_733),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_82),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_501),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_97),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_83),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_104),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_89),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_746),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_19),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_519),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_773),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_112),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_694),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_567),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_318),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_87),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_784),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_235),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_62),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_243),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_293),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_699),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_312),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_425),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_380),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_52),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_498),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_708),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_171),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_635),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_580),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_771),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_698),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_720),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_549),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_27),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_257),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_39),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_689),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_803),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_139),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_791),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_118),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_804),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_797),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_58),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_91),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_412),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_279),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_779),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_254),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_660),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_676),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_156),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_756),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_57),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_183),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_159),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_52),
.Y(n_1205)
);

CKINVDCx16_ASAP7_75t_R g1206 ( 
.A(n_159),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_22),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_247),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_154),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_915),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_813),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1007),
.B(n_800),
.Y(n_1212)
);

CKINVDCx16_ASAP7_75t_R g1213 ( 
.A(n_1021),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_816),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_835),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_1206),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_819),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_915),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_887),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_825),
.B(n_832),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_915),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_915),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_915),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_986),
.Y(n_1224)
);

INVxp33_ASAP7_75t_SL g1225 ( 
.A(n_991),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_893),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_915),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_881),
.B(n_1),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_899),
.B(n_2),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_947),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_880),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_823),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_880),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_880),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_863),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_938),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1073),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_994),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_833),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_855),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1112),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_837),
.Y(n_1242)
);

INVxp33_ASAP7_75t_SL g1243 ( 
.A(n_866),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_838),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_852),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1125),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1124),
.B(n_0),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_999),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_818),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1020),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_869),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_845),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_870),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1032),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_908),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_952),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1054),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_846),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_920),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_933),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_849),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1069),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1072),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_853),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_935),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_857),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_871),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1078),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1093),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1103),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1116),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1138),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_874),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1121),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1142),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_940),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1126),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_877),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_827),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_941),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_928),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_943),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_878),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_884),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_828),
.B(n_876),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_886),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_944),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_962),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_882),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_919),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_891),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_988),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_996),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_951),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1005),
.Y(n_1295)
);

CKINVDCx14_ASAP7_75t_R g1296 ( 
.A(n_1152),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_979),
.B(n_6),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1172),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1036),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_892),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_895),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1048),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1058),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1062),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1081),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1086),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1095),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1108),
.Y(n_1308)
);

INVxp33_ASAP7_75t_SL g1309 ( 
.A(n_814),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1114),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_897),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_900),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_902),
.Y(n_1313)
);

CKINVDCx16_ASAP7_75t_R g1314 ( 
.A(n_951),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_906),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_909),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1092),
.B(n_6),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1132),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1136),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_990),
.B(n_4),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1143),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1150),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_916),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_1119),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_824),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_830),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_918),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1164),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1167),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1175),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_931),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_934),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1187),
.Y(n_1333)
);

INVxp33_ASAP7_75t_L g1334 ( 
.A(n_1189),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_1119),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_937),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1207),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_939),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_990),
.B(n_4),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_942),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1208),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_949),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_815),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_953),
.Y(n_1344)
);

CKINVDCx16_ASAP7_75t_R g1345 ( 
.A(n_852),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_955),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_957),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_960),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_961),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_817),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_831),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_834),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_836),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_847),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_912),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_963),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_848),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_856),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_SL g1359 ( 
.A(n_912),
.Y(n_1359)
);

NOR2xp67_ASAP7_75t_L g1360 ( 
.A(n_1130),
.B(n_7),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_966),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_967),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1320),
.B(n_1130),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1211),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1325),
.B(n_822),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1231),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1233),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1234),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1326),
.B(n_860),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1210),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1343),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1218),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1220),
.A2(n_841),
.B1(n_842),
.B2(n_839),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1221),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1289),
.B(n_922),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1350),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1351),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1319),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1245),
.B(n_981),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1222),
.Y(n_1380)
);

AND2x6_ASAP7_75t_L g1381 ( 
.A(n_1223),
.B(n_1006),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1352),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1353),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1214),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1227),
.Y(n_1385)
);

XNOR2xp5_ASAP7_75t_L g1386 ( 
.A(n_1215),
.B(n_821),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1354),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1345),
.B(n_913),
.Y(n_1388)
);

CKINVDCx8_ASAP7_75t_R g1389 ( 
.A(n_1213),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1321),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1217),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1232),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1239),
.B(n_1076),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1296),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1328),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1219),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1249),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1216),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1357),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1355),
.B(n_1105),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1242),
.Y(n_1401)
);

BUFx8_ASAP7_75t_L g1402 ( 
.A(n_1359),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1358),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1251),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1255),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1259),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1260),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1244),
.B(n_1145),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1252),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1339),
.A2(n_864),
.B(n_859),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1235),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1265),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1276),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1279),
.B(n_913),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1280),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1243),
.A2(n_844),
.B1(n_851),
.B2(n_843),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1282),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1290),
.B(n_1258),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1287),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1288),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1224),
.B(n_888),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1236),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1292),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1293),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1295),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1299),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1302),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1237),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1309),
.B(n_890),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1303),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1281),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1304),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1360),
.A2(n_889),
.B(n_867),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1261),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1224),
.B(n_924),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1305),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1306),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1283),
.B(n_894),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1307),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1308),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1310),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1318),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1264),
.B(n_1178),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1285),
.B(n_948),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1266),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_SL g1446 ( 
.A(n_1294),
.B(n_971),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1322),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1267),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1273),
.B(n_820),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1329),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1330),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1333),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1337),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1278),
.B(n_826),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1341),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1246),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1240),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1284),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1253),
.B(n_1041),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1240),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1300),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1297),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1317),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1334),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1301),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1312),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1257),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1241),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1228),
.B(n_1026),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1316),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1323),
.B(n_829),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1331),
.B(n_850),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_SL g1473 ( 
.A(n_1314),
.B(n_971),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1247),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1332),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1338),
.B(n_854),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1340),
.Y(n_1477)
);

AND2x6_ASAP7_75t_L g1478 ( 
.A(n_1229),
.B(n_1006),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1324),
.B(n_1123),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1390),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1404),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1466),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1444),
.B(n_1344),
.Y(n_1483)
);

AND2x6_ASAP7_75t_L g1484 ( 
.A(n_1458),
.B(n_1006),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1366),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1406),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1378),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1364),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1412),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1410),
.A2(n_901),
.B(n_896),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1478),
.B(n_1346),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1449),
.B(n_1347),
.Y(n_1492)
);

NAND2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1464),
.B(n_1391),
.Y(n_1493)
);

NOR2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1384),
.B(n_858),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1378),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1467),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1395),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1395),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1478),
.B(n_1348),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1462),
.A2(n_1225),
.B1(n_1256),
.B2(n_1253),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1367),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1463),
.A2(n_1256),
.B1(n_1275),
.B2(n_1272),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1421),
.B(n_1349),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1429),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1419),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1368),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1478),
.B(n_1356),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1454),
.B(n_1361),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1379),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1420),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1474),
.A2(n_1298),
.B1(n_1212),
.B2(n_946),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1471),
.B(n_1286),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_1094),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1398),
.B(n_855),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1400),
.B(n_954),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1365),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1423),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1435),
.B(n_1335),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1459),
.B(n_1291),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1424),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1476),
.B(n_1311),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1425),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_L g1523 ( 
.A(n_1467),
.B(n_1002),
.C(n_998),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1370),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1372),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1418),
.B(n_1392),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1401),
.B(n_1313),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1375),
.B(n_1315),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1373),
.B(n_862),
.C(n_861),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1457),
.A2(n_1009),
.B1(n_1018),
.B2(n_875),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1402),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1374),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1393),
.B(n_1144),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1408),
.B(n_1327),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1414),
.B(n_1336),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_SL g1536 ( 
.A(n_1388),
.B(n_1342),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1396),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1405),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1380),
.Y(n_1539)
);

BUFx8_ASAP7_75t_SL g1540 ( 
.A(n_1431),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1427),
.Y(n_1541)
);

INVx5_ASAP7_75t_L g1542 ( 
.A(n_1381),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1430),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1446),
.B(n_1362),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1409),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1385),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1397),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1460),
.A2(n_1071),
.B1(n_1115),
.B2(n_1043),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1410),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1381),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1443),
.B(n_968),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1405),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1475),
.A2(n_1068),
.B1(n_872),
.B2(n_879),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1432),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1369),
.B(n_1226),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1473),
.B(n_1123),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1477),
.B(n_1359),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1434),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1394),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1363),
.B(n_972),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1407),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1445),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1436),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1432),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1439),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1441),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1440),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1413),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1461),
.B(n_1230),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1448),
.B(n_1238),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1441),
.Y(n_1571)
);

XNOR2xp5_ASAP7_75t_L g1572 ( 
.A(n_1386),
.B(n_1248),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1451),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1451),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1416),
.B(n_984),
.Y(n_1575)
);

NOR2x1p5_ASAP7_75t_L g1576 ( 
.A(n_1465),
.B(n_868),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1470),
.B(n_973),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1415),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1411),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1452),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1433),
.A2(n_1153),
.B1(n_1110),
.B2(n_1038),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1438),
.B(n_989),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1469),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1371),
.B(n_983),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1433),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1479),
.B(n_993),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1376),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1422),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1377),
.B(n_985),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1382),
.A2(n_1038),
.B1(n_1141),
.B2(n_1026),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1431),
.B(n_1068),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1428),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1417),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1453),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1483),
.B(n_1383),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1504),
.B(n_1250),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1492),
.B(n_1387),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1531),
.B(n_1468),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1481),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1516),
.A2(n_1262),
.B1(n_1263),
.B2(n_1254),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1528),
.B(n_1456),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1482),
.B(n_1389),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1508),
.B(n_1399),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1513),
.B(n_1403),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1511),
.B(n_885),
.C(n_883),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1533),
.B(n_905),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1551),
.B(n_914),
.Y(n_1608)
);

INVx8_ASAP7_75t_L g1609 ( 
.A(n_1537),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1503),
.B(n_1268),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1524),
.B(n_917),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1486),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1496),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1482),
.B(n_1426),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1512),
.B(n_1269),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1553),
.B(n_903),
.C(n_898),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1549),
.A2(n_1010),
.B1(n_1049),
.B2(n_982),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1489),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1480),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1521),
.B(n_1270),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1555),
.B(n_1271),
.Y(n_1621)
);

O2A1O1Ixp5_ASAP7_75t_L g1622 ( 
.A1(n_1549),
.A2(n_1585),
.B(n_1490),
.C(n_1510),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1534),
.B(n_1274),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1581),
.A2(n_1277),
.B1(n_1100),
.B2(n_1135),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1500),
.B(n_1386),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1525),
.B(n_921),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1532),
.B(n_923),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1539),
.B(n_927),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1505),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1491),
.B(n_987),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1571),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1529),
.B(n_907),
.C(n_904),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1518),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1499),
.B(n_1507),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1488),
.B(n_1437),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1546),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1558),
.B(n_997),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1585),
.A2(n_1447),
.B(n_1442),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1517),
.B(n_929),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1520),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1522),
.A2(n_1064),
.B1(n_956),
.B2(n_970),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1515),
.A2(n_1004),
.B1(n_1008),
.B2(n_1000),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1547),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1541),
.B(n_1543),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1575),
.A2(n_1455),
.B(n_1450),
.C(n_975),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1563),
.B(n_945),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1565),
.A2(n_978),
.B1(n_980),
.B2(n_977),
.Y(n_1647)
);

INVx8_ASAP7_75t_L g1648 ( 
.A(n_1540),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1490),
.A2(n_1017),
.B(n_995),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1577),
.B(n_873),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1576),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1562),
.B(n_1013),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1567),
.B(n_1023),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1561),
.Y(n_1654)
);

NOR3xp33_ASAP7_75t_L g1655 ( 
.A(n_1519),
.B(n_911),
.C(n_910),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1579),
.B(n_840),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1580),
.B(n_1024),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1526),
.B(n_926),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1514),
.B(n_930),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1530),
.A2(n_1159),
.B1(n_1088),
.B2(n_1051),
.C(n_1047),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1588),
.B(n_865),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1591),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1594),
.B(n_1045),
.Y(n_1663)
);

NAND2xp33_ASAP7_75t_L g1664 ( 
.A(n_1542),
.B(n_1014),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1514),
.B(n_936),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1515),
.B(n_1015),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1592),
.B(n_925),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1593),
.B(n_1578),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1559),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1568),
.B(n_1046),
.Y(n_1670)
);

NOR2xp67_ASAP7_75t_L g1671 ( 
.A(n_1545),
.B(n_1016),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1584),
.B(n_1050),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1583),
.B(n_1196),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1589),
.B(n_1059),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_L g1675 ( 
.A(n_1557),
.B(n_1022),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1587),
.B(n_1198),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1497),
.B(n_1063),
.Y(n_1677)
);

NAND2xp33_ASAP7_75t_L g1678 ( 
.A(n_1542),
.B(n_1025),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1501),
.B(n_1075),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1506),
.B(n_1079),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1556),
.A2(n_1523),
.B1(n_1502),
.B2(n_1582),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1485),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1493),
.B(n_1030),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1487),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1495),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1498),
.Y(n_1686)
);

NAND2xp33_ASAP7_75t_L g1687 ( 
.A(n_1542),
.B(n_1031),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1538),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1586),
.B(n_950),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1560),
.B(n_1087),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1566),
.B(n_932),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1574),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1484),
.B(n_1089),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1550),
.B(n_1191),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1484),
.B(n_1091),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1550),
.B(n_1194),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_L g1697 ( 
.A(n_1550),
.B(n_1034),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1569),
.B(n_1027),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1552),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1554),
.B(n_1066),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1484),
.B(n_1099),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1564),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1573),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1509),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1548),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1590),
.B(n_1104),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1494),
.B(n_1106),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1591),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1535),
.B(n_1109),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1536),
.A2(n_1035),
.B1(n_1039),
.B2(n_1037),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1572),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1544),
.B(n_1042),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1570),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1572),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1527),
.B(n_1082),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1531),
.B(n_1053),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1483),
.B(n_1127),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1480),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1496),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1549),
.A2(n_1131),
.B1(n_1156),
.B2(n_1129),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1481),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1481),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1496),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1571),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1483),
.B(n_1163),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1483),
.B(n_1174),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1481),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1516),
.B(n_1055),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1481),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1481),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1516),
.B(n_1056),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1481),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1480),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1483),
.A2(n_1061),
.B1(n_1065),
.B2(n_1057),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1483),
.B(n_1185),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1504),
.B(n_958),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1488),
.B(n_1067),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1483),
.B(n_1199),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1481),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1558),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1516),
.B(n_1070),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1504),
.B(n_1101),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1504),
.A2(n_1201),
.B1(n_1083),
.B2(n_1084),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1483),
.B(n_1381),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1480),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1481),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1481),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1516),
.B(n_1077),
.Y(n_1748)
);

NAND2xp33_ASAP7_75t_L g1749 ( 
.A(n_1491),
.B(n_1090),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1483),
.B(n_1107),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1483),
.B(n_1118),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1483),
.B(n_1120),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1607),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1719),
.Y(n_1754)
);

AOI21xp33_ASAP7_75t_L g1755 ( 
.A1(n_1717),
.A2(n_965),
.B(n_964),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1725),
.A2(n_1162),
.B(n_1200),
.C(n_959),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1599),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1649),
.A2(n_1038),
.B(n_1026),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1597),
.B(n_1603),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1638),
.A2(n_1141),
.B(n_1128),
.Y(n_1760)
);

OAI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1622),
.A2(n_295),
.B(n_294),
.Y(n_1761)
);

OAI321xp33_ASAP7_75t_L g1762 ( 
.A1(n_1726),
.A2(n_1141),
.A3(n_992),
.B1(n_974),
.B2(n_1001),
.C(n_976),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1607),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1634),
.A2(n_1134),
.B(n_1122),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1619),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1595),
.B(n_1137),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1735),
.A2(n_1140),
.B1(n_1146),
.B2(n_1139),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1656),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1600),
.B(n_1003),
.C(n_969),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1644),
.A2(n_1149),
.B(n_1147),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1718),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1604),
.A2(n_1157),
.B(n_1154),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1733),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1738),
.B(n_1740),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1750),
.B(n_1160),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1607),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1613),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1668),
.A2(n_1168),
.B(n_1161),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1650),
.A2(n_1170),
.B1(n_1171),
.B2(n_1169),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1624),
.A2(n_1705),
.B(n_1709),
.C(n_1660),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1612),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_L g1782 ( 
.A(n_1744),
.B(n_1173),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1176),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1752),
.B(n_1177),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1631),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1608),
.A2(n_1180),
.B(n_1179),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1615),
.B(n_1011),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1596),
.B(n_1012),
.Y(n_1788)
);

AOI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1690),
.A2(n_1186),
.B(n_1181),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1609),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1623),
.B(n_1019),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1742),
.B(n_1028),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1745),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1672),
.A2(n_1190),
.B(n_1188),
.Y(n_1794)
);

OAI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1720),
.A2(n_1197),
.B(n_1195),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_L g1796 ( 
.A1(n_1736),
.A2(n_1658),
.B(n_1681),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1617),
.A2(n_1033),
.B1(n_1040),
.B2(n_1029),
.Y(n_1797)
);

NOR2x2_ASAP7_75t_L g1798 ( 
.A(n_1598),
.B(n_1044),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1618),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1674),
.A2(n_1060),
.B(n_1052),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1636),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1643),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1723),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1635),
.B(n_1074),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1629),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1606),
.B(n_1080),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1640),
.A2(n_1165),
.B(n_1158),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1630),
.A2(n_1096),
.B(n_1085),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1721),
.B(n_1097),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1722),
.B(n_1098),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1727),
.Y(n_1811)
);

AOI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1639),
.A2(n_305),
.B(n_297),
.Y(n_1812)
);

AO21x1_ASAP7_75t_L g1813 ( 
.A1(n_1689),
.A2(n_7),
.B(n_8),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1729),
.Y(n_1814)
);

O2A1O1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1707),
.A2(n_1646),
.B(n_1657),
.C(n_1653),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1730),
.A2(n_1111),
.B(n_1113),
.C(n_1102),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1732),
.B(n_1117),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1631),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1631),
.Y(n_1819)
);

CKINVDCx10_ASAP7_75t_R g1820 ( 
.A(n_1598),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1739),
.A2(n_1148),
.B(n_1133),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1746),
.A2(n_1155),
.B(n_1151),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1698),
.B(n_1166),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1747),
.A2(n_1183),
.B(n_1182),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1601),
.B(n_1184),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1642),
.A2(n_1193),
.B1(n_1202),
.B2(n_1192),
.Y(n_1826)
);

NAND2x1p5_ASAP7_75t_L g1827 ( 
.A(n_1724),
.B(n_307),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1692),
.B(n_1203),
.Y(n_1828)
);

OR2x2_ASAP7_75t_SL g1829 ( 
.A(n_1625),
.B(n_1204),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1663),
.A2(n_1209),
.B(n_1205),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1666),
.A2(n_310),
.B(n_308),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1633),
.A2(n_1614),
.B1(n_1734),
.B2(n_1632),
.Y(n_1832)
);

INVx8_ASAP7_75t_L g1833 ( 
.A(n_1609),
.Y(n_1833)
);

AOI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1611),
.A2(n_315),
.B(n_314),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1737),
.B(n_316),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_R g1836 ( 
.A(n_1711),
.B(n_317),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1691),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1675),
.B(n_319),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1621),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1682),
.Y(n_1840)
);

O2A1O1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1749),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1654),
.B(n_1679),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1680),
.B(n_9),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1661),
.B(n_320),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1724),
.Y(n_1845)
);

NOR3xp33_ASAP7_75t_L g1846 ( 
.A(n_1620),
.B(n_10),
.C(n_11),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1715),
.A2(n_323),
.B1(n_324),
.B2(n_322),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1626),
.A2(n_326),
.B(n_325),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_R g1849 ( 
.A(n_1651),
.B(n_327),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1673),
.A2(n_330),
.B(n_329),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1714),
.B(n_12),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1627),
.B(n_13),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1724),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1628),
.B(n_13),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1670),
.B(n_14),
.Y(n_1855)
);

BUFx4f_ASAP7_75t_L g1856 ( 
.A(n_1648),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1712),
.A2(n_333),
.B(n_332),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1728),
.A2(n_336),
.B(n_334),
.Y(n_1858)
);

OAI321xp33_ASAP7_75t_L g1859 ( 
.A1(n_1616),
.A2(n_16),
.A3(n_18),
.B1(n_14),
.B2(n_15),
.C(n_17),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1671),
.B(n_16),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1667),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1648),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1700),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1645),
.A2(n_338),
.B(n_337),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1743),
.B(n_1688),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1669),
.B(n_17),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1731),
.A2(n_340),
.B(n_339),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1741),
.A2(n_344),
.B(n_341),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1713),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1748),
.A2(n_348),
.B(n_345),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1686),
.B(n_18),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1685),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1684),
.B(n_19),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1699),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1637),
.B(n_20),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1704),
.B(n_349),
.Y(n_1876)
);

AOI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1676),
.A2(n_352),
.B(n_350),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1702),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1677),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1605),
.A2(n_354),
.B(n_353),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1652),
.B(n_21),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1683),
.A2(n_1678),
.B(n_1664),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1647),
.B(n_21),
.Y(n_1883)
);

O2A1O1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1706),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1710),
.A2(n_356),
.B(n_355),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1641),
.B(n_23),
.Y(n_1886)
);

OAI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1655),
.A2(n_25),
.B(n_26),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_L g1888 ( 
.A(n_1610),
.B(n_25),
.C(n_28),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1602),
.B(n_1703),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1708),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1890)
);

NAND3xp33_ASAP7_75t_SL g1891 ( 
.A(n_1659),
.B(n_29),
.C(n_30),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1665),
.B(n_31),
.C(n_32),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1687),
.A2(n_359),
.B(n_358),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1694),
.B(n_31),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1696),
.A2(n_361),
.B(n_360),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1662),
.B(n_32),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1697),
.A2(n_363),
.B(n_362),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1693),
.A2(n_1701),
.B(n_1695),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1716),
.Y(n_1899)
);

O2A1O1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1717),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1900)
);

NOR2xp67_ASAP7_75t_L g1901 ( 
.A(n_1740),
.B(n_365),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1597),
.B(n_366),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1619),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1692),
.Y(n_1904)
);

BUFx12f_ASAP7_75t_L g1905 ( 
.A(n_1598),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1607),
.Y(n_1906)
);

OAI321xp33_ASAP7_75t_L g1907 ( 
.A1(n_1717),
.A2(n_36),
.A3(n_38),
.B1(n_34),
.B2(n_35),
.C(n_37),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_R g1908 ( 
.A(n_1740),
.B(n_368),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1622),
.A2(n_371),
.B(n_370),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1597),
.B(n_36),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1649),
.A2(n_373),
.B(n_372),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1597),
.B(n_37),
.Y(n_1912)
);

INVx8_ASAP7_75t_L g1913 ( 
.A(n_1609),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1597),
.B(n_38),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1597),
.B(n_39),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1597),
.B(n_40),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1599),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1649),
.A2(n_375),
.B(n_374),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1649),
.A2(n_378),
.B(n_377),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1649),
.A2(n_383),
.B(n_382),
.Y(n_1920)
);

AO21x1_ASAP7_75t_L g1921 ( 
.A1(n_1717),
.A2(n_40),
.B(n_41),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1602),
.B(n_384),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1717),
.A2(n_387),
.B1(n_391),
.B2(n_386),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1649),
.A2(n_395),
.B(n_392),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1649),
.A2(n_398),
.B(n_397),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1597),
.A2(n_403),
.B1(n_405),
.B2(n_399),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1597),
.B(n_406),
.Y(n_1927)
);

O2A1O1Ixp5_ASAP7_75t_L g1928 ( 
.A1(n_1717),
.A2(n_410),
.B(n_413),
.C(n_408),
.Y(n_1928)
);

NAND2x1p5_ASAP7_75t_L g1929 ( 
.A(n_1904),
.B(n_414),
.Y(n_1929)
);

O2A1O1Ixp33_ASAP7_75t_SL g1930 ( 
.A1(n_1902),
.A2(n_416),
.B(n_418),
.C(n_415),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1759),
.A2(n_421),
.B(n_419),
.Y(n_1931)
);

AO21x1_ASAP7_75t_L g1932 ( 
.A1(n_1909),
.A2(n_41),
.B(n_42),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1763),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1815),
.A2(n_1882),
.B(n_1842),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1862),
.B(n_422),
.Y(n_1935)
);

AOI21x1_ASAP7_75t_L g1936 ( 
.A1(n_1758),
.A2(n_426),
.B(n_424),
.Y(n_1936)
);

INVx5_ASAP7_75t_L g1937 ( 
.A(n_1763),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1787),
.B(n_43),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1775),
.A2(n_430),
.B(n_428),
.Y(n_1939)
);

OAI21xp33_ASAP7_75t_SL g1940 ( 
.A1(n_1910),
.A2(n_43),
.B(n_44),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1796),
.A2(n_434),
.B1(n_435),
.B2(n_431),
.Y(n_1941)
);

BUFx3_ASAP7_75t_L g1942 ( 
.A(n_1833),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1790),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1774),
.B(n_436),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1791),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1788),
.A2(n_442),
.B1(n_444),
.B2(n_441),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1826),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.C(n_48),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1833),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1765),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1754),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1863),
.B(n_445),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1792),
.B(n_45),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1823),
.B(n_47),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1766),
.B(n_1803),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1879),
.B(n_447),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1771),
.Y(n_1956)
);

OAI21xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1912),
.A2(n_48),
.B(n_49),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1913),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_R g1959 ( 
.A(n_1913),
.B(n_1856),
.Y(n_1959)
);

NAND3xp33_ASAP7_75t_SL g1960 ( 
.A(n_1769),
.B(n_50),
.C(n_51),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1914),
.B(n_448),
.Y(n_1961)
);

BUFx8_ASAP7_75t_L g1962 ( 
.A(n_1905),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1879),
.B(n_450),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_R g1964 ( 
.A(n_1789),
.B(n_451),
.Y(n_1964)
);

O2A1O1Ixp5_ASAP7_75t_L g1965 ( 
.A1(n_1784),
.A2(n_454),
.B(n_456),
.C(n_452),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1839),
.B(n_50),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1777),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1837),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1828),
.Y(n_1969)
);

A2O1A1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1780),
.A2(n_54),
.B(n_51),
.C(n_53),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1869),
.B(n_459),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1915),
.B(n_53),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1916),
.B(n_460),
.Y(n_1973)
);

INVx5_ASAP7_75t_L g1974 ( 
.A(n_1776),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1776),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_R g1976 ( 
.A(n_1820),
.B(n_461),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1757),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_SL g1978 ( 
.A1(n_1829),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1768),
.B(n_464),
.Y(n_1979)
);

O2A1O1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1887),
.A2(n_58),
.B(n_55),
.C(n_56),
.Y(n_1980)
);

INVxp67_ASAP7_75t_L g1981 ( 
.A(n_1851),
.Y(n_1981)
);

BUFx12f_ASAP7_75t_L g1982 ( 
.A(n_1785),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1781),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1806),
.B(n_59),
.Y(n_1984)
);

O2A1O1Ixp5_ASAP7_75t_L g1985 ( 
.A1(n_1885),
.A2(n_1864),
.B(n_1783),
.C(n_1860),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1799),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1865),
.A2(n_469),
.B1(n_470),
.B2(n_467),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1861),
.B(n_471),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1911),
.A2(n_1925),
.B(n_1924),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1805),
.B(n_1811),
.Y(n_1990)
);

CKINVDCx8_ASAP7_75t_R g1991 ( 
.A(n_1785),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1818),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1814),
.A2(n_473),
.B1(n_476),
.B2(n_472),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1917),
.A2(n_479),
.B1(n_481),
.B2(n_478),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1875),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1761),
.A2(n_487),
.B(n_486),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1836),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1832),
.B(n_488),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1840),
.B(n_63),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1918),
.A2(n_491),
.B(n_489),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1818),
.Y(n_2001)
);

BUFx3_ASAP7_75t_L g2002 ( 
.A(n_1819),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1819),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1773),
.B(n_63),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1872),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1919),
.A2(n_1920),
.B(n_1898),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1901),
.B(n_492),
.Y(n_2007)
);

INVx8_ASAP7_75t_L g2008 ( 
.A(n_1845),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1755),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1881),
.B(n_493),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1793),
.B(n_64),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1801),
.B(n_67),
.Y(n_2012)
);

INVx4_ASAP7_75t_L g2013 ( 
.A(n_1845),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1782),
.A2(n_499),
.B(n_494),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1802),
.Y(n_2015)
);

NOR3xp33_ASAP7_75t_L g2016 ( 
.A(n_1891),
.B(n_1762),
.C(n_1892),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1927),
.A2(n_502),
.B(n_500),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1846),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1804),
.B(n_70),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1903),
.B(n_70),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1807),
.B(n_71),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1844),
.A2(n_505),
.B(n_503),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1848),
.A2(n_507),
.B(n_506),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1908),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1896),
.B(n_72),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_R g2026 ( 
.A(n_1753),
.B(n_509),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1928),
.A2(n_511),
.B(n_510),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_R g2028 ( 
.A(n_1853),
.B(n_512),
.Y(n_2028)
);

OAI21xp33_ASAP7_75t_L g2029 ( 
.A1(n_1795),
.A2(n_1824),
.B(n_1866),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1830),
.B(n_73),
.Y(n_2030)
);

NAND3xp33_ASAP7_75t_SL g2031 ( 
.A(n_1888),
.B(n_74),
.C(n_75),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1838),
.A2(n_515),
.B(n_514),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1906),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1878),
.Y(n_2034)
);

AOI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1835),
.A2(n_1868),
.B(n_1857),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1873),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1889),
.A2(n_520),
.B(n_517),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1906),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1874),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1899),
.B(n_74),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1876),
.Y(n_2041)
);

NAND3xp33_ASAP7_75t_L g2042 ( 
.A(n_1779),
.B(n_75),
.C(n_76),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1756),
.B(n_523),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1880),
.A2(n_525),
.B(n_524),
.Y(n_2044)
);

INVx4_ASAP7_75t_L g2045 ( 
.A(n_1827),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1849),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1977),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1954),
.B(n_1825),
.Y(n_2048)
);

OAI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1996),
.A2(n_1877),
.B(n_1834),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1983),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1982),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_2006),
.A2(n_1897),
.B(n_1893),
.Y(n_2052)
);

INVx4_ASAP7_75t_L g2053 ( 
.A(n_1937),
.Y(n_2053)
);

NAND2x1p5_ASAP7_75t_L g2054 ( 
.A(n_1937),
.B(n_1922),
.Y(n_2054)
);

OAI22x1_ASAP7_75t_L g2055 ( 
.A1(n_1938),
.A2(n_1953),
.B1(n_2019),
.B2(n_2042),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1989),
.A2(n_1895),
.B(n_1831),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1986),
.Y(n_2057)
);

NAND2x1p5_ASAP7_75t_L g2058 ( 
.A(n_1937),
.B(n_1847),
.Y(n_2058)
);

AO31x2_ASAP7_75t_L g2059 ( 
.A1(n_1932),
.A2(n_1813),
.A3(n_1921),
.B(n_1923),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1934),
.A2(n_1812),
.B(n_1858),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1950),
.Y(n_2061)
);

A2O1A1Ixp33_ASAP7_75t_L g2062 ( 
.A1(n_2029),
.A2(n_1841),
.B(n_1808),
.C(n_1800),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_2035),
.A2(n_1870),
.B(n_1867),
.Y(n_2063)
);

AO31x2_ASAP7_75t_L g2064 ( 
.A1(n_2023),
.A2(n_1816),
.A3(n_1843),
.B(n_1852),
.Y(n_2064)
);

OAI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2030),
.A2(n_1883),
.B1(n_1894),
.B2(n_1907),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1990),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2005),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2036),
.B(n_1809),
.Y(n_2068)
);

INVx2_ASAP7_75t_SL g2069 ( 
.A(n_2008),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1985),
.A2(n_1850),
.B(n_1760),
.Y(n_2070)
);

AO21x1_ASAP7_75t_L g2071 ( 
.A1(n_1998),
.A2(n_2044),
.B(n_2021),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2027),
.A2(n_2000),
.B(n_2007),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2014),
.A2(n_1855),
.B(n_1854),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_1936),
.A2(n_1871),
.B(n_1764),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_2008),
.B(n_1886),
.Y(n_2075)
);

INVx3_ASAP7_75t_SL g2076 ( 
.A(n_1948),
.Y(n_2076)
);

AOI221x1_ASAP7_75t_L g2077 ( 
.A1(n_2016),
.A2(n_1890),
.B1(n_1767),
.B2(n_1772),
.C(n_1786),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1967),
.B(n_1810),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1968),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_1974),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2034),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1961),
.A2(n_1770),
.B(n_1794),
.Y(n_2082)
);

OAI21x1_ASAP7_75t_L g2083 ( 
.A1(n_1965),
.A2(n_2017),
.B(n_2037),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1973),
.A2(n_1817),
.B(n_1926),
.Y(n_2084)
);

NAND2x1p5_ASAP7_75t_L g2085 ( 
.A(n_1974),
.B(n_1821),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1984),
.B(n_1822),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_L g2087 ( 
.A1(n_1939),
.A2(n_1884),
.B(n_1778),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_1991),
.Y(n_2088)
);

INVx3_ASAP7_75t_L g2089 ( 
.A(n_1974),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1975),
.Y(n_2090)
);

OAI22x1_ASAP7_75t_L g2091 ( 
.A1(n_1966),
.A2(n_1859),
.B1(n_1798),
.B2(n_1900),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1959),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1952),
.B(n_1797),
.Y(n_2093)
);

AO32x2_ASAP7_75t_L g2094 ( 
.A1(n_1978),
.A2(n_79),
.A3(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_2094)
);

OR2x6_ASAP7_75t_L g2095 ( 
.A(n_1942),
.B(n_1969),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_2001),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_1981),
.B(n_77),
.Y(n_2097)
);

O2A1O1Ixp33_ASAP7_75t_L g2098 ( 
.A1(n_2031),
.A2(n_81),
.B(n_78),
.C(n_80),
.Y(n_2098)
);

OA21x2_ASAP7_75t_L g2099 ( 
.A1(n_2043),
.A2(n_527),
.B(n_526),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1972),
.B(n_81),
.Y(n_2100)
);

AO31x2_ASAP7_75t_L g2101 ( 
.A1(n_1970),
.A2(n_530),
.A3(n_531),
.B(n_529),
.Y(n_2101)
);

A2O1A1Ixp33_ASAP7_75t_L g2102 ( 
.A1(n_1980),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1931),
.A2(n_533),
.B(n_532),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_SL g2104 ( 
.A(n_1997),
.B(n_84),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_2002),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_2022),
.A2(n_536),
.B(n_535),
.Y(n_2106)
);

AOI21x1_ASAP7_75t_L g2107 ( 
.A1(n_2010),
.A2(n_810),
.B(n_538),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1949),
.Y(n_2108)
);

A2O1A1Ixp33_ASAP7_75t_L g2109 ( 
.A1(n_2009),
.A2(n_90),
.B(n_86),
.C(n_88),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_2033),
.Y(n_2110)
);

OA21x2_ASAP7_75t_L g2111 ( 
.A1(n_2004),
.A2(n_2012),
.B(n_2011),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1944),
.A2(n_539),
.B(n_537),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_L g2113 ( 
.A1(n_2032),
.A2(n_2020),
.B(n_1987),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1956),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2015),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2039),
.Y(n_2116)
);

AOI221x1_ASAP7_75t_L g2117 ( 
.A1(n_1960),
.A2(n_92),
.B1(n_86),
.B2(n_91),
.C(n_93),
.Y(n_2117)
);

INVx4_ASAP7_75t_L g2118 ( 
.A(n_2033),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2041),
.A2(n_545),
.B(n_543),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1999),
.Y(n_2120)
);

OAI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_2040),
.A2(n_547),
.B(n_546),
.Y(n_2121)
);

AOI21xp5_ASAP7_75t_L g2122 ( 
.A1(n_1979),
.A2(n_553),
.B(n_548),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_1943),
.Y(n_2123)
);

OAI21x1_ASAP7_75t_L g2124 ( 
.A1(n_1941),
.A2(n_556),
.B(n_555),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_1988),
.A2(n_558),
.B(n_557),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2025),
.B(n_92),
.Y(n_2126)
);

AO32x2_ASAP7_75t_L g2127 ( 
.A1(n_1993),
.A2(n_96),
.A3(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1971),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_L g2129 ( 
.A1(n_1951),
.A2(n_563),
.B(n_560),
.Y(n_2129)
);

INVx5_ASAP7_75t_L g2130 ( 
.A(n_2038),
.Y(n_2130)
);

AO31x2_ASAP7_75t_L g2131 ( 
.A1(n_1994),
.A2(n_565),
.A3(n_566),
.B(n_564),
.Y(n_2131)
);

BUFx12f_ASAP7_75t_L g2132 ( 
.A(n_1962),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2038),
.Y(n_2133)
);

OA21x2_ASAP7_75t_L g2134 ( 
.A1(n_1946),
.A2(n_570),
.B(n_568),
.Y(n_2134)
);

OAI21x1_ASAP7_75t_L g2135 ( 
.A1(n_1929),
.A2(n_581),
.B(n_575),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_2046),
.B(n_94),
.Y(n_2136)
);

AOI221xp5_ASAP7_75t_L g2137 ( 
.A1(n_2018),
.A2(n_99),
.B1(n_95),
.B2(n_98),
.C(n_100),
.Y(n_2137)
);

CKINVDCx20_ASAP7_75t_R g2138 ( 
.A(n_1958),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_SL g2139 ( 
.A1(n_2048),
.A2(n_1940),
.B1(n_1957),
.B2(n_1976),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2061),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2066),
.B(n_2024),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_2079),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2050),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_2055),
.A2(n_1947),
.B1(n_1995),
.B2(n_2045),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_SL g2145 ( 
.A1(n_2137),
.A2(n_1945),
.B(n_1955),
.Y(n_2145)
);

OAI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2117),
.A2(n_1933),
.B1(n_2013),
.B2(n_2003),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_SL g2147 ( 
.A1(n_2098),
.A2(n_1963),
.B(n_1935),
.Y(n_2147)
);

CKINVDCx20_ASAP7_75t_R g2148 ( 
.A(n_2138),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2057),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_2091),
.A2(n_1964),
.B1(n_2028),
.B2(n_2026),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_2047),
.Y(n_2151)
);

BUFx10_ASAP7_75t_L g2152 ( 
.A(n_2051),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_2065),
.A2(n_1992),
.B1(n_1930),
.B2(n_100),
.Y(n_2153)
);

OAI22xp33_ASAP7_75t_L g2154 ( 
.A1(n_2068),
.A2(n_102),
.B1(n_98),
.B2(n_99),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2120),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2155)
);

BUFx10_ASAP7_75t_L g2156 ( 
.A(n_2051),
.Y(n_2156)
);

BUFx12f_ASAP7_75t_L g2157 ( 
.A(n_2132),
.Y(n_2157)
);

BUFx10_ASAP7_75t_L g2158 ( 
.A(n_2092),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_2130),
.Y(n_2159)
);

BUFx12f_ASAP7_75t_L g2160 ( 
.A(n_2118),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2071),
.A2(n_107),
.B1(n_103),
.B2(n_105),
.Y(n_2161)
);

CKINVDCx6p67_ASAP7_75t_R g2162 ( 
.A(n_2130),
.Y(n_2162)
);

OAI22xp33_ASAP7_75t_L g2163 ( 
.A1(n_2093),
.A2(n_108),
.B1(n_105),
.B2(n_107),
.Y(n_2163)
);

AOI22xp33_ASAP7_75t_SL g2164 ( 
.A1(n_2121),
.A2(n_111),
.B1(n_108),
.B2(n_109),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2067),
.Y(n_2165)
);

NAND2x1p5_ASAP7_75t_L g2166 ( 
.A(n_2053),
.B(n_582),
.Y(n_2166)
);

BUFx8_ASAP7_75t_SL g2167 ( 
.A(n_2105),
.Y(n_2167)
);

AOI22xp33_ASAP7_75t_SL g2168 ( 
.A1(n_2100),
.A2(n_113),
.B1(n_109),
.B2(n_112),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2081),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_2088),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2126),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_2110),
.Y(n_2172)
);

BUFx2_ASAP7_75t_L g2173 ( 
.A(n_2133),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_SL g2174 ( 
.A1(n_2086),
.A2(n_2058),
.B1(n_2134),
.B2(n_2084),
.Y(n_2174)
);

CKINVDCx11_ASAP7_75t_R g2175 ( 
.A(n_2076),
.Y(n_2175)
);

INVx1_ASAP7_75t_SL g2176 ( 
.A(n_2123),
.Y(n_2176)
);

INVx8_ASAP7_75t_L g2177 ( 
.A(n_2095),
.Y(n_2177)
);

OAI22x1_ASAP7_75t_SL g2178 ( 
.A1(n_2090),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_2095),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_SL g2180 ( 
.A1(n_2124),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_SL g2181 ( 
.A1(n_2072),
.A2(n_2128),
.B1(n_2112),
.B2(n_2075),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2108),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2114),
.Y(n_2183)
);

OAI21xp33_ASAP7_75t_SL g2184 ( 
.A1(n_2129),
.A2(n_584),
.B(n_583),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_SL g2185 ( 
.A1(n_2075),
.A2(n_124),
.B1(n_120),
.B2(n_123),
.Y(n_2185)
);

OAI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_2078),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2115),
.Y(n_2187)
);

AOI22xp33_ASAP7_75t_L g2188 ( 
.A1(n_2104),
.A2(n_2136),
.B1(n_2111),
.B2(n_2085),
.Y(n_2188)
);

BUFx12f_ASAP7_75t_L g2189 ( 
.A(n_2069),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2116),
.B(n_125),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_2089),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_SL g2192 ( 
.A1(n_2056),
.A2(n_2122),
.B1(n_2125),
.B2(n_2094),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2127),
.Y(n_2193)
);

BUFx3_ASAP7_75t_L g2194 ( 
.A(n_2080),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2107),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2097),
.B(n_127),
.Y(n_2196)
);

BUFx10_ASAP7_75t_L g2197 ( 
.A(n_2096),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2094),
.B(n_127),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2054),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_2199)
);

NAND2x1p5_ASAP7_75t_L g2200 ( 
.A(n_2135),
.B(n_586),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2109),
.B(n_128),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2106),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2127),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_2102),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_2204)
);

CKINVDCx11_ASAP7_75t_R g2205 ( 
.A(n_2077),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2101),
.Y(n_2206)
);

BUFx2_ASAP7_75t_L g2207 ( 
.A(n_2059),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_2119),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2062),
.B(n_131),
.Y(n_2209)
);

INVx4_ASAP7_75t_L g2210 ( 
.A(n_2099),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2103),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2142),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2143),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2140),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2201),
.B(n_2059),
.Y(n_2215)
);

BUFx2_ASAP7_75t_L g2216 ( 
.A(n_2206),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2165),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2151),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2151),
.B(n_2064),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_2207),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2207),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2182),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_2193),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2169),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2183),
.Y(n_2225)
);

OAI21x1_ASAP7_75t_L g2226 ( 
.A1(n_2211),
.A2(n_2060),
.B(n_2052),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2187),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2149),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2139),
.B(n_2101),
.Y(n_2229)
);

BUFx2_ASAP7_75t_L g2230 ( 
.A(n_2203),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_2173),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_2172),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2150),
.A2(n_2073),
.B1(n_2082),
.B2(n_2070),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2190),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2209),
.Y(n_2235)
);

NAND2x1_ASAP7_75t_L g2236 ( 
.A(n_2210),
.B(n_2113),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2141),
.B(n_2064),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2198),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2197),
.Y(n_2239)
);

BUFx2_ASAP7_75t_L g2240 ( 
.A(n_2202),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2205),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2195),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2188),
.B(n_2131),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2174),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_2167),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_2172),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2194),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2168),
.B(n_2131),
.Y(n_2248)
);

AO21x2_ASAP7_75t_L g2249 ( 
.A1(n_2204),
.A2(n_2074),
.B(n_2049),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2145),
.A2(n_2087),
.B(n_2083),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2144),
.B(n_587),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_2148),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2196),
.Y(n_2253)
);

BUFx3_ASAP7_75t_L g2254 ( 
.A(n_2160),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2177),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2177),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2181),
.Y(n_2257)
);

OAI21x1_ASAP7_75t_L g2258 ( 
.A1(n_2200),
.A2(n_2063),
.B(n_592),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_2162),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2185),
.B(n_591),
.Y(n_2260)
);

AO21x2_ASAP7_75t_L g2261 ( 
.A1(n_2146),
.A2(n_133),
.B(n_134),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2163),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_2159),
.Y(n_2263)
);

OAI21x1_ASAP7_75t_L g2264 ( 
.A1(n_2153),
.A2(n_2161),
.B(n_2166),
.Y(n_2264)
);

INVx2_ASAP7_75t_SL g2265 ( 
.A(n_2152),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2154),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2186),
.Y(n_2267)
);

BUFx6f_ASAP7_75t_L g2268 ( 
.A(n_2170),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2171),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_2191),
.B(n_593),
.Y(n_2270)
);

INVx5_ASAP7_75t_L g2271 ( 
.A(n_2189),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2192),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2208),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2179),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2170),
.B(n_2176),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_2175),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2147),
.B(n_134),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2199),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_2158),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2156),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2180),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_2155),
.B(n_594),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2164),
.B(n_135),
.Y(n_2283)
);

OR2x2_ASAP7_75t_L g2284 ( 
.A(n_2238),
.B(n_135),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2212),
.B(n_596),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2215),
.B(n_136),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_SL g2287 ( 
.A(n_2245),
.B(n_2157),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_2281),
.A2(n_2184),
.B1(n_2178),
.B2(n_138),
.Y(n_2288)
);

NAND4xp25_ASAP7_75t_L g2289 ( 
.A(n_2283),
.B(n_138),
.C(n_136),
.D(n_137),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_2231),
.B(n_597),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2282),
.A2(n_141),
.B1(n_137),
.B2(n_140),
.Y(n_2291)
);

OR2x6_ASAP7_75t_L g2292 ( 
.A(n_2273),
.B(n_598),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2224),
.Y(n_2293)
);

OAI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2233),
.A2(n_600),
.B(n_599),
.Y(n_2294)
);

NOR2x1_ASAP7_75t_SL g2295 ( 
.A(n_2261),
.B(n_602),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2235),
.B(n_140),
.Y(n_2296)
);

BUFx5_ASAP7_75t_L g2297 ( 
.A(n_2242),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2253),
.B(n_142),
.Y(n_2298)
);

OAI21x1_ASAP7_75t_L g2299 ( 
.A1(n_2226),
.A2(n_604),
.B(n_603),
.Y(n_2299)
);

A2O1A1Ixp33_ASAP7_75t_L g2300 ( 
.A1(n_2264),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_SL g2301 ( 
.A(n_2276),
.B(n_2252),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2218),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2272),
.B(n_143),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2214),
.B(n_144),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2225),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2221),
.Y(n_2306)
);

AO21x2_ASAP7_75t_L g2307 ( 
.A1(n_2250),
.A2(n_145),
.B(n_146),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2217),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2275),
.B(n_607),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2221),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_2232),
.Y(n_2311)
);

AO21x2_ASAP7_75t_L g2312 ( 
.A1(n_2243),
.A2(n_145),
.B(n_146),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2220),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2234),
.B(n_147),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2228),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2282),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2219),
.B(n_148),
.Y(n_2317)
);

OAI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2251),
.A2(n_611),
.B(n_609),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2229),
.B(n_149),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2220),
.Y(n_2320)
);

OR2x2_ASAP7_75t_L g2321 ( 
.A(n_2237),
.B(n_150),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2222),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2227),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2275),
.B(n_614),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2223),
.B(n_151),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2223),
.B(n_151),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2244),
.B(n_152),
.Y(n_2327)
);

OA21x2_ASAP7_75t_L g2328 ( 
.A1(n_2257),
.A2(n_152),
.B(n_153),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2230),
.Y(n_2329)
);

OR2x6_ASAP7_75t_L g2330 ( 
.A(n_2276),
.B(n_616),
.Y(n_2330)
);

AOI22xp33_ASAP7_75t_L g2331 ( 
.A1(n_2241),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2274),
.B(n_155),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2213),
.Y(n_2333)
);

O2A1O1Ixp33_ASAP7_75t_SL g2334 ( 
.A1(n_2277),
.A2(n_2269),
.B(n_2266),
.C(n_2262),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_2230),
.B(n_156),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2216),
.B(n_157),
.Y(n_2336)
);

INVx1_ASAP7_75t_SL g2337 ( 
.A(n_2247),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2239),
.B(n_158),
.Y(n_2338)
);

OAI21x1_ASAP7_75t_L g2339 ( 
.A1(n_2236),
.A2(n_618),
.B(n_617),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2248),
.B(n_160),
.Y(n_2340)
);

NOR2x1_ASAP7_75t_SL g2341 ( 
.A(n_2249),
.B(n_620),
.Y(n_2341)
);

INVx4_ASAP7_75t_L g2342 ( 
.A(n_2232),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2216),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_2240),
.B(n_160),
.Y(n_2344)
);

OAI21x1_ASAP7_75t_SL g2345 ( 
.A1(n_2278),
.A2(n_161),
.B(n_162),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2240),
.Y(n_2346)
);

AOI22xp33_ASAP7_75t_L g2347 ( 
.A1(n_2289),
.A2(n_2267),
.B1(n_2260),
.B2(n_2279),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2293),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2305),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2306),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2310),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2302),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2313),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2337),
.B(n_2255),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_2311),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2329),
.B(n_2346),
.Y(n_2356)
);

OAI222xp33_ASAP7_75t_L g2357 ( 
.A1(n_2291),
.A2(n_2271),
.B1(n_2256),
.B2(n_2236),
.C1(n_2270),
.C2(n_2280),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2320),
.B(n_2268),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2343),
.B(n_2258),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2315),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2308),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2322),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2323),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2319),
.B(n_2268),
.Y(n_2364)
);

INVxp67_ASAP7_75t_L g2365 ( 
.A(n_2311),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2333),
.Y(n_2366)
);

INVxp67_ASAP7_75t_SL g2367 ( 
.A(n_2297),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2297),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2340),
.B(n_2265),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2297),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2297),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2336),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2286),
.B(n_2271),
.Y(n_2373)
);

AOI22xp33_ASAP7_75t_SL g2374 ( 
.A1(n_2295),
.A2(n_2271),
.B1(n_2270),
.B2(n_2259),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2344),
.Y(n_2375)
);

OAI22xp5_ASAP7_75t_SL g2376 ( 
.A1(n_2288),
.A2(n_2254),
.B1(n_2246),
.B2(n_2263),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2325),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2317),
.B(n_2246),
.Y(n_2378)
);

INVxp67_ASAP7_75t_SL g2379 ( 
.A(n_2326),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2342),
.B(n_162),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_2335),
.B(n_2321),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2338),
.B(n_164),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2312),
.B(n_164),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2284),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2307),
.B(n_165),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2290),
.B(n_166),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2334),
.B(n_166),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2298),
.B(n_168),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2348),
.Y(n_2389)
);

AO21x2_ASAP7_75t_L g2390 ( 
.A1(n_2367),
.A2(n_2341),
.B(n_2300),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2349),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2378),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2379),
.B(n_2327),
.Y(n_2393)
);

INVx1_ASAP7_75t_SL g2394 ( 
.A(n_2354),
.Y(n_2394)
);

OAI221xp5_ASAP7_75t_L g2395 ( 
.A1(n_2347),
.A2(n_2316),
.B1(n_2331),
.B2(n_2318),
.C(n_2294),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2381),
.B(n_2301),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_2356),
.B(n_2314),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2381),
.B(n_2287),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2355),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2356),
.B(n_2296),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_2375),
.B(n_2304),
.Y(n_2401)
);

NAND4xp25_ASAP7_75t_L g2402 ( 
.A(n_2385),
.B(n_2303),
.C(n_2332),
.D(n_2285),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2358),
.B(n_2328),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2350),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2360),
.B(n_2292),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2372),
.B(n_2292),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2373),
.B(n_2330),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2352),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2351),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2376),
.A2(n_2330),
.B1(n_2345),
.B2(n_2309),
.Y(n_2410)
);

AO21x2_ASAP7_75t_L g2411 ( 
.A1(n_2385),
.A2(n_2299),
.B(n_2339),
.Y(n_2411)
);

OAI31xp33_ASAP7_75t_L g2412 ( 
.A1(n_2376),
.A2(n_2324),
.A3(n_172),
.B(n_169),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2363),
.Y(n_2413)
);

AOI221xp5_ASAP7_75t_L g2414 ( 
.A1(n_2387),
.A2(n_172),
.B1(n_169),
.B2(n_170),
.C(n_173),
.Y(n_2414)
);

INVx3_ASAP7_75t_L g2415 ( 
.A(n_2361),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2377),
.B(n_173),
.Y(n_2416)
);

NAND4xp25_ASAP7_75t_L g2417 ( 
.A(n_2387),
.B(n_176),
.C(n_174),
.D(n_175),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2366),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2353),
.B(n_175),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2384),
.B(n_176),
.Y(n_2420)
);

OAI33xp33_ASAP7_75t_L g2421 ( 
.A1(n_2359),
.A2(n_177),
.A3(n_178),
.B1(n_179),
.B2(n_180),
.B3(n_181),
.Y(n_2421)
);

OR2x6_ASAP7_75t_L g2422 ( 
.A(n_2383),
.B(n_178),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2362),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2359),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2368),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2370),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2364),
.B(n_179),
.Y(n_2427)
);

NAND4xp25_ASAP7_75t_L g2428 ( 
.A(n_2383),
.B(n_182),
.C(n_180),
.D(n_181),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2371),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2369),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2365),
.B(n_183),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2380),
.B(n_184),
.Y(n_2432)
);

INVx4_ASAP7_75t_L g2433 ( 
.A(n_2386),
.Y(n_2433)
);

AOI33xp33_ASAP7_75t_L g2434 ( 
.A1(n_2388),
.A2(n_2374),
.A3(n_2382),
.B1(n_2386),
.B2(n_187),
.B3(n_188),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2374),
.B(n_184),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2357),
.Y(n_2436)
);

BUFx3_ASAP7_75t_L g2437 ( 
.A(n_2357),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2381),
.B(n_185),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2360),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2394),
.B(n_185),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2397),
.B(n_186),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2429),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2403),
.B(n_187),
.Y(n_2443)
);

AND2x4_ASAP7_75t_SL g2444 ( 
.A(n_2399),
.B(n_188),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2392),
.B(n_189),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2439),
.B(n_189),
.Y(n_2446)
);

AND2x4_ASAP7_75t_L g2447 ( 
.A(n_2398),
.B(n_190),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2430),
.B(n_191),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2396),
.B(n_191),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2429),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2400),
.B(n_192),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2424),
.B(n_192),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2406),
.B(n_193),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2409),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2409),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2436),
.B(n_2413),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2405),
.B(n_193),
.Y(n_2457)
);

OAI33xp33_ASAP7_75t_L g2458 ( 
.A1(n_2417),
.A2(n_2436),
.A3(n_2428),
.B1(n_2389),
.B2(n_2404),
.B3(n_2393),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2391),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2418),
.B(n_194),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2425),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2408),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2423),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2415),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2405),
.B(n_194),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2415),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2401),
.B(n_195),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2426),
.Y(n_2468)
);

INVx3_ASAP7_75t_SL g2469 ( 
.A(n_2422),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2419),
.Y(n_2470)
);

NAND2x1p5_ASAP7_75t_L g2471 ( 
.A(n_2433),
.B(n_195),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2437),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2416),
.Y(n_2473)
);

OR2x2_ASAP7_75t_L g2474 ( 
.A(n_2411),
.B(n_196),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2433),
.B(n_196),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2420),
.Y(n_2476)
);

HB1xp67_ASAP7_75t_L g2477 ( 
.A(n_2390),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2399),
.Y(n_2478)
);

OR2x2_ASAP7_75t_L g2479 ( 
.A(n_2402),
.B(n_197),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2438),
.B(n_197),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_R g2481 ( 
.A(n_2435),
.B(n_198),
.Y(n_2481)
);

INVxp67_ASAP7_75t_L g2482 ( 
.A(n_2432),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2407),
.B(n_198),
.Y(n_2483)
);

HB1xp67_ASAP7_75t_L g2484 ( 
.A(n_2422),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2399),
.B(n_199),
.Y(n_2485)
);

BUFx3_ASAP7_75t_L g2486 ( 
.A(n_2431),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2427),
.B(n_199),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2454),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2472),
.B(n_2434),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2472),
.B(n_2414),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2478),
.B(n_2410),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2455),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2456),
.B(n_2412),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2459),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2462),
.Y(n_2495)
);

NOR2xp67_ASAP7_75t_L g2496 ( 
.A(n_2477),
.B(n_2395),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2443),
.B(n_200),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2463),
.Y(n_2498)
);

NAND2x1_ASAP7_75t_SL g2499 ( 
.A(n_2469),
.B(n_2421),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2470),
.B(n_201),
.Y(n_2500)
);

INVx2_ASAP7_75t_SL g2501 ( 
.A(n_2484),
.Y(n_2501)
);

HB1xp67_ASAP7_75t_L g2502 ( 
.A(n_2474),
.Y(n_2502)
);

INVx1_ASAP7_75t_SL g2503 ( 
.A(n_2444),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2470),
.B(n_201),
.Y(n_2504)
);

NAND2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2446),
.B(n_202),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2468),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2468),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2473),
.B(n_203),
.Y(n_2508)
);

BUFx3_ASAP7_75t_L g2509 ( 
.A(n_2447),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2461),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2476),
.B(n_203),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2464),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2441),
.B(n_204),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2464),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2466),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2486),
.B(n_204),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2452),
.B(n_205),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2442),
.B(n_2450),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2466),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2460),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2440),
.Y(n_2521)
);

NOR2x1_ASAP7_75t_L g2522 ( 
.A(n_2451),
.B(n_205),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2448),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2457),
.B(n_2465),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2447),
.B(n_206),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2453),
.B(n_206),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2445),
.Y(n_2527)
);

OR2x2_ASAP7_75t_L g2528 ( 
.A(n_2479),
.B(n_207),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2475),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2449),
.B(n_2483),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2482),
.B(n_207),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2506),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2491),
.B(n_2485),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2509),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_2496),
.B(n_2481),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2488),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2492),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2501),
.B(n_2502),
.Y(n_2538)
);

OR2x2_ASAP7_75t_L g2539 ( 
.A(n_2520),
.B(n_2467),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2494),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2489),
.B(n_2487),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2490),
.B(n_2480),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2529),
.B(n_2471),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2495),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2507),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2498),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2493),
.B(n_2499),
.Y(n_2547)
);

OR2x2_ASAP7_75t_L g2548 ( 
.A(n_2521),
.B(n_2458),
.Y(n_2548)
);

OR2x2_ASAP7_75t_L g2549 ( 
.A(n_2510),
.B(n_208),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2499),
.B(n_2527),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2518),
.B(n_208),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2512),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2523),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2553)
);

INVxp67_ASAP7_75t_SL g2554 ( 
.A(n_2522),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2514),
.Y(n_2555)
);

INVx1_ASAP7_75t_SL g2556 ( 
.A(n_2503),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2528),
.B(n_211),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2500),
.B(n_212),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2524),
.B(n_214),
.Y(n_2559)
);

INVxp33_ASAP7_75t_L g2560 ( 
.A(n_2530),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2504),
.B(n_214),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2532),
.Y(n_2562)
);

OAI211xp5_ASAP7_75t_L g2563 ( 
.A1(n_2535),
.A2(n_2517),
.B(n_2513),
.C(n_2497),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2532),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2556),
.B(n_2525),
.Y(n_2565)
);

OAI32xp33_ASAP7_75t_L g2566 ( 
.A1(n_2547),
.A2(n_2505),
.A3(n_2511),
.B1(n_2508),
.B2(n_2515),
.Y(n_2566)
);

AOI21xp33_ASAP7_75t_L g2567 ( 
.A1(n_2548),
.A2(n_2519),
.B(n_2531),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2552),
.Y(n_2568)
);

XOR2x2_ASAP7_75t_SL g2569 ( 
.A(n_2550),
.B(n_2525),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2534),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2555),
.Y(n_2571)
);

NAND3xp33_ASAP7_75t_L g2572 ( 
.A(n_2554),
.B(n_2516),
.C(n_2526),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2533),
.B(n_215),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2542),
.A2(n_216),
.B(n_217),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2543),
.Y(n_2575)
);

INVx1_ASAP7_75t_SL g2576 ( 
.A(n_2559),
.Y(n_2576)
);

OR2x2_ASAP7_75t_L g2577 ( 
.A(n_2538),
.B(n_217),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2545),
.Y(n_2578)
);

OAI322xp33_ASAP7_75t_L g2579 ( 
.A1(n_2553),
.A2(n_218),
.A3(n_219),
.B1(n_220),
.B2(n_221),
.C1(n_222),
.C2(n_224),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2541),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2560),
.B(n_222),
.Y(n_2581)
);

AOI221xp5_ASAP7_75t_L g2582 ( 
.A1(n_2546),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.C(n_229),
.Y(n_2582)
);

NAND3x1_ASAP7_75t_L g2583 ( 
.A(n_2558),
.B(n_225),
.C(n_228),
.Y(n_2583)
);

AOI221xp5_ASAP7_75t_L g2584 ( 
.A1(n_2540),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.C(n_232),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2536),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2551),
.B(n_230),
.Y(n_2586)
);

OAI321xp33_ASAP7_75t_L g2587 ( 
.A1(n_2544),
.A2(n_234),
.A3(n_235),
.B1(n_236),
.B2(n_237),
.C(n_238),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2539),
.B(n_236),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2537),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2562),
.Y(n_2590)
);

AOI21xp33_ASAP7_75t_L g2591 ( 
.A1(n_2566),
.A2(n_2549),
.B(n_2557),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2564),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2574),
.B(n_2561),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2565),
.B(n_237),
.Y(n_2594)
);

O2A1O1Ixp33_ASAP7_75t_L g2595 ( 
.A1(n_2567),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2568),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2576),
.B(n_239),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2570),
.B(n_241),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2583),
.B(n_242),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2571),
.Y(n_2600)
);

XNOR2x1_ASAP7_75t_L g2601 ( 
.A(n_2580),
.B(n_243),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2575),
.B(n_244),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2581),
.B(n_245),
.Y(n_2603)
);

NOR3xp33_ASAP7_75t_L g2604 ( 
.A(n_2563),
.B(n_245),
.C(n_246),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2572),
.B(n_2580),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2577),
.A2(n_249),
.B1(n_246),
.B2(n_248),
.Y(n_2606)
);

INVx1_ASAP7_75t_SL g2607 ( 
.A(n_2586),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2569),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2588),
.B(n_248),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2582),
.A2(n_2584),
.B1(n_2579),
.B2(n_2585),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2589),
.A2(n_252),
.B1(n_249),
.B2(n_250),
.Y(n_2611)
);

INVx1_ASAP7_75t_SL g2612 ( 
.A(n_2573),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_SL g2613 ( 
.A1(n_2587),
.A2(n_254),
.B1(n_250),
.B2(n_253),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2578),
.Y(n_2614)
);

XNOR2xp5_ASAP7_75t_L g2615 ( 
.A(n_2572),
.B(n_253),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2562),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2574),
.B(n_255),
.Y(n_2617)
);

OAI222xp33_ASAP7_75t_L g2618 ( 
.A1(n_2580),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.C1(n_259),
.C2(n_260),
.Y(n_2618)
);

AOI31xp33_ASAP7_75t_L g2619 ( 
.A1(n_2567),
.A2(n_260),
.A3(n_256),
.B(n_258),
.Y(n_2619)
);

AOI322xp5_ASAP7_75t_L g2620 ( 
.A1(n_2567),
.A2(n_261),
.A3(n_262),
.B1(n_263),
.B2(n_264),
.C1(n_265),
.C2(n_267),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2565),
.B(n_262),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2574),
.B(n_267),
.Y(n_2622)
);

INVxp67_ASAP7_75t_L g2623 ( 
.A(n_2565),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2597),
.Y(n_2624)
);

INVxp67_ASAP7_75t_SL g2625 ( 
.A(n_2599),
.Y(n_2625)
);

INVx1_ASAP7_75t_SL g2626 ( 
.A(n_2607),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2604),
.B(n_268),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2598),
.Y(n_2628)
);

INVx2_ASAP7_75t_SL g2629 ( 
.A(n_2602),
.Y(n_2629)
);

NOR3xp33_ASAP7_75t_L g2630 ( 
.A(n_2623),
.B(n_269),
.C(n_270),
.Y(n_2630)
);

OAI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2605),
.A2(n_270),
.B(n_271),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2593),
.A2(n_271),
.B(n_273),
.Y(n_2632)
);

OR2x2_ASAP7_75t_L g2633 ( 
.A(n_2612),
.B(n_273),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2608),
.B(n_274),
.Y(n_2634)
);

NOR3xp33_ASAP7_75t_L g2635 ( 
.A(n_2591),
.B(n_274),
.C(n_275),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2603),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2621),
.B(n_275),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2594),
.B(n_276),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2590),
.Y(n_2639)
);

XNOR2xp5_ASAP7_75t_L g2640 ( 
.A(n_2615),
.B(n_276),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2601),
.B(n_2619),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2592),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2620),
.B(n_2610),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2617),
.B(n_277),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2622),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2609),
.B(n_277),
.Y(n_2646)
);

AOI21xp33_ASAP7_75t_SL g2647 ( 
.A1(n_2613),
.A2(n_278),
.B(n_279),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2616),
.Y(n_2648)
);

AOI211x1_ASAP7_75t_L g2649 ( 
.A1(n_2643),
.A2(n_2618),
.B(n_2596),
.C(n_2614),
.Y(n_2649)
);

INVxp67_ASAP7_75t_SL g2650 ( 
.A(n_2640),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2626),
.B(n_2600),
.Y(n_2651)
);

INVxp67_ASAP7_75t_L g2652 ( 
.A(n_2625),
.Y(n_2652)
);

NOR3xp33_ASAP7_75t_L g2653 ( 
.A(n_2635),
.B(n_2595),
.C(n_2613),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2629),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2641),
.B(n_2606),
.Y(n_2655)
);

INVxp67_ASAP7_75t_SL g2656 ( 
.A(n_2633),
.Y(n_2656)
);

INVx1_ASAP7_75t_SL g2657 ( 
.A(n_2638),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2624),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2637),
.Y(n_2659)
);

INVxp67_ASAP7_75t_SL g2660 ( 
.A(n_2634),
.Y(n_2660)
);

NAND4xp25_ASAP7_75t_L g2661 ( 
.A(n_2645),
.B(n_2636),
.C(n_2632),
.D(n_2628),
.Y(n_2661)
);

AOI221xp5_ASAP7_75t_L g2662 ( 
.A1(n_2647),
.A2(n_2611),
.B1(n_280),
.B2(n_281),
.C(n_282),
.Y(n_2662)
);

NAND4xp25_ASAP7_75t_L g2663 ( 
.A(n_2631),
.B(n_281),
.C(n_278),
.D(n_280),
.Y(n_2663)
);

NAND5xp2_ASAP7_75t_L g2664 ( 
.A(n_2639),
.B(n_282),
.C(n_283),
.D(n_284),
.E(n_285),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2630),
.B(n_283),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2646),
.Y(n_2666)
);

NOR3xp33_ASAP7_75t_L g2667 ( 
.A(n_2627),
.B(n_285),
.C(n_286),
.Y(n_2667)
);

AOI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2644),
.A2(n_287),
.B(n_288),
.Y(n_2668)
);

NAND4xp75_ASAP7_75t_L g2669 ( 
.A(n_2642),
.B(n_287),
.C(n_288),
.D(n_289),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2648),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2647),
.B(n_291),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2647),
.B(n_291),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_L g2673 ( 
.A(n_2641),
.B(n_292),
.Y(n_2673)
);

AOI221xp5_ASAP7_75t_L g2674 ( 
.A1(n_2643),
.A2(n_292),
.B1(n_293),
.B2(n_621),
.C(n_622),
.Y(n_2674)
);

CKINVDCx6p67_ASAP7_75t_R g2675 ( 
.A(n_2626),
.Y(n_2675)
);

NOR3x1_ASAP7_75t_L g2676 ( 
.A(n_2643),
.B(n_623),
.C(n_624),
.Y(n_2676)
);

NOR3xp33_ASAP7_75t_L g2677 ( 
.A(n_2635),
.B(n_625),
.C(n_627),
.Y(n_2677)
);

OAI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2635),
.A2(n_628),
.B(n_630),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2624),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2647),
.B(n_631),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2626),
.B(n_634),
.Y(n_2681)
);

AOI211xp5_ASAP7_75t_L g2682 ( 
.A1(n_2653),
.A2(n_636),
.B(n_638),
.C(n_639),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2675),
.Y(n_2683)
);

CKINVDCx20_ASAP7_75t_R g2684 ( 
.A(n_2657),
.Y(n_2684)
);

AOI221xp5_ASAP7_75t_L g2685 ( 
.A1(n_2649),
.A2(n_641),
.B1(n_642),
.B2(n_643),
.C(n_645),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2650),
.A2(n_648),
.B1(n_649),
.B2(n_651),
.Y(n_2686)
);

NAND4xp25_ASAP7_75t_L g2687 ( 
.A(n_2655),
.B(n_652),
.C(n_653),
.D(n_656),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2656),
.B(n_809),
.Y(n_2688)
);

NAND4xp25_ASAP7_75t_L g2689 ( 
.A(n_2661),
.B(n_657),
.C(n_659),
.D(n_661),
.Y(n_2689)
);

OAI211xp5_ASAP7_75t_L g2690 ( 
.A1(n_2662),
.A2(n_662),
.B(n_663),
.C(n_664),
.Y(n_2690)
);

AOI211xp5_ASAP7_75t_L g2691 ( 
.A1(n_2672),
.A2(n_665),
.B(n_666),
.C(n_667),
.Y(n_2691)
);

AOI322xp5_ASAP7_75t_L g2692 ( 
.A1(n_2673),
.A2(n_668),
.A3(n_670),
.B1(n_672),
.B2(n_673),
.C1(n_675),
.C2(n_679),
.Y(n_2692)
);

AOI221xp5_ASAP7_75t_L g2693 ( 
.A1(n_2652),
.A2(n_680),
.B1(n_681),
.B2(n_682),
.C(n_683),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2654),
.A2(n_684),
.B1(n_685),
.B2(n_688),
.Y(n_2694)
);

NAND4xp25_ASAP7_75t_L g2695 ( 
.A(n_2651),
.B(n_690),
.C(n_691),
.D(n_693),
.Y(n_2695)
);

OAI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2674),
.A2(n_2671),
.B1(n_2660),
.B2(n_2666),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2668),
.B(n_808),
.Y(n_2697)
);

NOR2x1_ASAP7_75t_L g2698 ( 
.A(n_2669),
.B(n_696),
.Y(n_2698)
);

NAND4xp75_ASAP7_75t_L g2699 ( 
.A(n_2676),
.B(n_807),
.C(n_701),
.D(n_705),
.Y(n_2699)
);

AOI322xp5_ASAP7_75t_L g2700 ( 
.A1(n_2667),
.A2(n_700),
.A3(n_707),
.B1(n_709),
.B2(n_710),
.C1(n_711),
.C2(n_713),
.Y(n_2700)
);

INVx1_ASAP7_75t_SL g2701 ( 
.A(n_2681),
.Y(n_2701)
);

AOI21xp33_ASAP7_75t_SL g2702 ( 
.A1(n_2683),
.A2(n_2665),
.B(n_2658),
.Y(n_2702)
);

NAND3xp33_ASAP7_75t_L g2703 ( 
.A(n_2685),
.B(n_2679),
.C(n_2677),
.Y(n_2703)
);

NOR3xp33_ASAP7_75t_L g2704 ( 
.A(n_2696),
.B(n_2659),
.C(n_2663),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2684),
.Y(n_2705)
);

NAND3xp33_ASAP7_75t_L g2706 ( 
.A(n_2698),
.B(n_2670),
.C(n_2678),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2701),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2697),
.A2(n_2680),
.B(n_2664),
.Y(n_2708)
);

AND3x1_ASAP7_75t_L g2709 ( 
.A(n_2691),
.B(n_714),
.C(n_715),
.Y(n_2709)
);

NAND4xp75_ASAP7_75t_L g2710 ( 
.A(n_2688),
.B(n_716),
.C(n_718),
.D(n_719),
.Y(n_2710)
);

NAND5xp2_ASAP7_75t_L g2711 ( 
.A(n_2690),
.B(n_721),
.C(n_722),
.D(n_723),
.E(n_725),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2705),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2707),
.B(n_2699),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2710),
.Y(n_2714)
);

NAND4xp75_ASAP7_75t_L g2715 ( 
.A(n_2708),
.B(n_2686),
.C(n_2693),
.D(n_2700),
.Y(n_2715)
);

NAND4xp75_ASAP7_75t_L g2716 ( 
.A(n_2712),
.B(n_2709),
.C(n_2702),
.D(n_2704),
.Y(n_2716)
);

INVx4_ASAP7_75t_L g2717 ( 
.A(n_2716),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2717),
.A2(n_2706),
.B1(n_2703),
.B2(n_2714),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2718),
.B(n_2713),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2719),
.A2(n_2715),
.B1(n_2689),
.B2(n_2695),
.Y(n_2720)
);

OAI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2720),
.A2(n_2682),
.B(n_2687),
.Y(n_2721)
);

OAI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2721),
.A2(n_2694),
.B(n_2692),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2722),
.B(n_2711),
.Y(n_2723)
);

AOI22x1_ASAP7_75t_L g2724 ( 
.A1(n_2723),
.A2(n_726),
.B1(n_727),
.B2(n_728),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2724),
.A2(n_729),
.B1(n_730),
.B2(n_731),
.Y(n_2725)
);

AOI211xp5_ASAP7_75t_L g2726 ( 
.A1(n_2725),
.A2(n_732),
.B(n_734),
.C(n_735),
.Y(n_2726)
);


endmodule