module real_jpeg_28703_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_0),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_0),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_0),
.A2(n_26),
.B1(n_48),
.B2(n_50),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_1),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_169),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_169),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_169),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_2),
.B(n_48),
.Y(n_86)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_2),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_4),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_95),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_95),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_4),
.A2(n_48),
.B1(n_50),
.B2(n_95),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_6),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_28),
.B(n_32),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_6),
.B(n_30),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_6),
.A2(n_54),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_6),
.B(n_54),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_69),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_6),
.A2(n_85),
.B1(n_89),
.B2(n_251),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_6),
.A2(n_31),
.B(n_267),
.Y(n_266)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_127),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_9),
.A2(n_48),
.B1(n_50),
.B2(n_127),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_127),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_50),
.A3(n_54),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_11),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_12),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_174)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_15),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_158),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_158),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_15),
.A2(n_48),
.B1(n_50),
.B2(n_158),
.Y(n_245)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_17),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_97),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_17),
.A2(n_54),
.B1(n_55),
.B2(n_97),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_17),
.A2(n_48),
.B1(n_50),
.B2(n_97),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_335),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_77),
.B(n_331),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_21),
.B(n_37),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_21),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_23),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_25),
.A2(n_34),
.B(n_167),
.C(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_27),
.A2(n_30),
.B1(n_94),
.B2(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_27),
.A2(n_30),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_27),
.A2(n_30),
.B1(n_126),
.B2(n_198),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_27),
.A2(n_30),
.B(n_35),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_31),
.A2(n_62),
.B(n_64),
.C(n_67),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_65),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g275 ( 
.A1(n_31),
.A2(n_55),
.A3(n_65),
.B1(n_268),
.B2(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_32),
.B(n_167),
.Y(n_268)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_70),
.C(n_72),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_38),
.A2(n_39),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_40),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_42),
.A2(n_74),
.B1(n_76),
.B2(n_96),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_46),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_46),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_46),
.A2(n_58),
.B1(n_136),
.B2(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_47),
.A2(n_52),
.B1(n_57),
.B2(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_47),
.A2(n_52),
.B1(n_103),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_47),
.A2(n_52),
.B1(n_122),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_47),
.A2(n_52),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_47),
.A2(n_52),
.B1(n_225),
.B2(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_47),
.B(n_167),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_47),
.A2(n_52),
.B1(n_163),
.B2(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_48),
.B(n_51),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_48),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_54),
.B(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_58),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_69),
.B1(n_112),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_60),
.A2(n_69),
.B1(n_157),
.B2(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_60),
.A2(n_69),
.B1(n_124),
.B2(n_201),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_67),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_67),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_61),
.A2(n_67),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_61),
.A2(n_67),
.B1(n_159),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_61),
.A2(n_67),
.B1(n_181),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_65),
.Y(n_277)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_70),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_76),
.B1(n_93),
.B2(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_74),
.A2(n_76),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_324),
.B(n_330),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_139),
.A3(n_148),
.B1(n_322),
.B2(n_323),
.C(n_341),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_128),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_80),
.B(n_128),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_109),
.C(n_116),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_81),
.B(n_109),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_98),
.B1(n_99),
.B2(n_108),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_92),
.B(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_83),
.A2(n_84),
.B1(n_100),
.B2(n_101),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_90),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_87),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_85),
.A2(n_87),
.B1(n_120),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_85),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_85),
.A2(n_89),
.B1(n_245),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_85),
.A2(n_87),
.B1(n_239),
.B2(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_86),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_86),
.A2(n_88),
.B1(n_174),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_86),
.A2(n_88),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g240 ( 
.A(n_88),
.Y(n_240)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_104),
.A2(n_107),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_104),
.A2(n_107),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_114),
.B(n_115),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_114),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_129),
.CI(n_138),
.CON(n_128),
.SN(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_129),
.C(n_138),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_116),
.A2(n_117),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.C(n_125),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_118),
.B(n_123),
.CI(n_125),
.CON(n_305),
.SN(n_305)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_121),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_128),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_137),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_131),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_133),
.C(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_131),
.B(n_146),
.C(n_147),
.Y(n_325)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_140),
.B(n_141),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_303),
.A3(n_311),
.B1(n_316),
.B2(n_321),
.C(n_342),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_203),
.C(n_215),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_185),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_185),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_170),
.C(n_177),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_152),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_165),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_160),
.B2(n_161),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_161),
.C(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_170),
.A2(n_177),
.B1(n_178),
.B2(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_170),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_173),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_179),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_182),
.B(n_184),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_183),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_192),
.C(n_193),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_190),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_202),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_199),
.C(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_204),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_205),
.B(n_206),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_208),
.B(n_209),
.C(n_214),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_297),
.B(n_302),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_283),
.B(n_296),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_261),
.B(n_282),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_241),
.B(n_260),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_220),
.B(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_235),
.C(n_237),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_236),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_248),
.B(n_259),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_247),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_253),
.B(n_258),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_250),
.B(n_252),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_274),
.B1(n_280),
.B2(n_281),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_264)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_273),
.C(n_281),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_271),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_274),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_292),
.C(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_305),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_312),
.A2(n_317),
.B(n_320),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule