module real_jpeg_33526_n_5 (n_4, n_0, n_1, n_2, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_5;

wire n_17;
wire n_12;
wire n_8;
wire n_18;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire n_6;
wire n_7;
wire n_16;
wire n_13;
wire n_9;

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_16),
.Y(n_15)
);

BUFx2_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_13),
.Y(n_12)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g5 ( 
.A1(n_6),
.A2(n_10),
.B1(n_17),
.B2(n_18),
.Y(n_5)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g6 ( 
.A1(n_7),
.A2(n_8),
.B(n_9),
.Y(n_6)
);

NAND2xp33_ASAP7_75t_SL g9 ( 
.A(n_7),
.B(n_8),
.Y(n_9)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g10 ( 
.A1(n_11),
.A2(n_14),
.B(n_15),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);


endmodule