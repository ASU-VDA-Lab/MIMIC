module real_jpeg_6732_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_0),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_0),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_0),
.A2(n_184),
.B1(n_254),
.B2(n_257),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_0),
.A2(n_89),
.B1(n_91),
.B2(n_184),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_0),
.A2(n_184),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_2),
.A2(n_63),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_2),
.A2(n_63),
.B1(n_363),
.B2(n_384),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_2),
.A2(n_63),
.B1(n_322),
.B2(n_434),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_3),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_3),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_3),
.Y(n_221)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_3),
.Y(n_242)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_4),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_4),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_4),
.Y(n_357)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_4),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_5),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_93),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_5),
.A2(n_93),
.B1(n_276),
.B2(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_5),
.A2(n_93),
.B1(n_159),
.B2(n_284),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_6),
.A2(n_56),
.B1(n_187),
.B2(n_310),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_6),
.A2(n_56),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_6),
.A2(n_56),
.B1(n_396),
.B2(n_399),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_7),
.A2(n_149),
.B1(n_152),
.B2(n_155),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_7),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_7),
.B(n_170),
.C(n_174),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_7),
.B(n_78),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_7),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_7),
.B(n_123),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_11),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_11),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_11),
.A2(n_162),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_11),
.A2(n_162),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_11),
.A2(n_162),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_13),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_13),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_98),
.B1(n_110),
.B2(n_125),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_13),
.A2(n_98),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_14),
.Y(n_120)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_14),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_15),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_15),
.A2(n_125),
.B1(n_275),
.B2(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_15),
.A2(n_275),
.B1(n_389),
.B2(n_392),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g448 ( 
.A1(n_15),
.A2(n_275),
.B1(n_403),
.B2(n_449),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_16),
.A2(n_168),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_16),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_16),
.A2(n_207),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_16),
.A2(n_207),
.B1(n_282),
.B2(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_16),
.A2(n_60),
.B1(n_207),
.B2(n_403),
.Y(n_422)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_525),
.B(n_528),
.Y(n_25)
);

AO21x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_138),
.B(n_524),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_136),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_28),
.B(n_136),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_127),
.C(n_133),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_29),
.A2(n_30),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_64),
.C(n_99),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_31),
.B(n_512),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_32),
.A2(n_57),
.B1(n_59),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_32),
.A2(n_57),
.B1(n_128),
.B2(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_32),
.A2(n_354),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_32),
.A2(n_41),
.B1(n_401),
.B2(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_32),
.A2(n_50),
.B1(n_57),
.B2(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_33),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_33),
.B(n_355),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_33),
.A2(n_58),
.B(n_527),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_36),
.Y(n_330)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_41),
.B(n_155),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_42),
.Y(n_332)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_45),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_45),
.Y(n_391)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_46),
.Y(n_303)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_48),
.Y(n_394)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_57),
.A2(n_422),
.B(n_450),
.Y(n_460)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_58),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_58),
.B(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_64),
.A2(n_99),
.B1(n_100),
.B2(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_64),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_65),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_65),
.A2(n_94),
.B1(n_300),
.B2(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_65),
.A2(n_94),
.B1(n_388),
.B2(n_395),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_65),
.A2(n_88),
.B1(n_94),
.B2(n_501),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_71),
.Y(n_263)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_77),
.Y(n_268)
);

INVx6_ASAP7_75t_L g436 ( 
.A(n_77),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_78),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g423 ( 
.A1(n_78),
.A2(n_134),
.B1(n_305),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_78),
.A2(n_134),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_80),
.Y(n_286)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_84),
.Y(n_384)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_86),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_86),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_86),
.Y(n_363)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_91),
.A2(n_155),
.B(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_94),
.B(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_94),
.A2(n_300),
.B(n_304),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_99),
.A2(n_100),
.B1(n_499),
.B2(n_500),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_99),
.B(n_496),
.C(n_499),
.Y(n_507)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_122),
.B(n_124),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_148),
.B(n_156),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_101),
.A2(n_122),
.B1(n_206),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_101),
.A2(n_156),
.B(n_253),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_101),
.A2(n_122),
.B1(n_362),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_102),
.B(n_157),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_102),
.A2(n_123),
.B1(n_382),
.B2(n_385),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_102),
.A2(n_123),
.B1(n_385),
.B2(n_410),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_102),
.A2(n_123),
.B1(n_410),
.B2(n_439),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_103)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_104),
.Y(n_383)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_107),
.Y(n_257)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_112),
.A2(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_118),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_118),
.Y(n_276)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_120),
.Y(n_345)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_120),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_122),
.A2(n_211),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_124),
.Y(n_439)
);

INVx5_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_127),
.B(n_133),
.Y(n_521)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_132),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_134),
.A2(n_260),
.B(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_134),
.B(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_134),
.A2(n_264),
.B(n_463),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_136),
.B(n_526),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_136),
.B(n_526),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_137),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_518),
.B(n_523),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_489),
.B(n_515),
.Y(n_139)
);

OAI311xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_366),
.A3(n_465),
.B1(n_483),
.C1(n_484),
.Y(n_140)
);

AOI21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_315),
.B(n_365),
.Y(n_141)
);

AO21x1_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_291),
.B(n_314),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_247),
.B(n_290),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_214),
.B(n_246),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_179),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_146),
.B(n_179),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_165),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_147),
.A2(n_165),
.B1(n_166),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_155),
.A2(n_189),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_155),
.B(n_334),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_155),
.A2(n_326),
.B(n_333),
.Y(n_352)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_177),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_203),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_180),
.B(n_204),
.C(n_213),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_189),
.B(n_197),
.Y(n_180)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_189),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_189),
.A2(n_372),
.B1(n_375),
.B2(n_377),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_189),
.A2(n_230),
.B(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_200),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_190),
.A2(n_272),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_190),
.A2(n_340),
.B1(n_418),
.B2(n_419),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_198),
.Y(n_338)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_201),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_235),
.B(n_245),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_223),
.B(n_234),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_221),
.Y(n_376)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_221),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_233),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_233),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_232),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_226),
.Y(n_311)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_227),
.Y(n_380)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_232),
.A2(n_271),
.B(n_277),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_243),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_243),
.Y(n_245)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_249),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_269),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_258),
.B2(n_259),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_258),
.C(n_269),
.Y(n_292)
);

INVx3_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI32xp33_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_281),
.A3(n_283),
.B1(n_285),
.B2(n_287),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_280),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_293),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_298),
.B2(n_313),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_297),
.C(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_306),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_307),
.C(n_308),
.Y(n_346)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_303),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_303),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_316),
.B(n_317),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_349),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_318)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_335),
.B2(n_336),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_321),
.B(n_335),
.Y(n_461)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_325),
.A3(n_330),
.B1(n_331),
.B2(n_333),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_346),
.B(n_347),
.C(n_349),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_358),
.B2(n_364),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_350),
.B(n_359),
.C(n_361),
.Y(n_474)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_360),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_451),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_SL g484 ( 
.A1(n_367),
.A2(n_451),
.B(n_485),
.C(n_488),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_425),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_368),
.B(n_425),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_407),
.C(n_413),
.Y(n_368)
);

FAx1_ASAP7_75t_SL g464 ( 
.A(n_369),
.B(n_407),
.CI(n_413),
.CON(n_464),
.SN(n_464)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_386),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_370),
.B(n_387),
.C(n_400),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_381),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_371),
.B(n_381),
.Y(n_457)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_400),
.Y(n_386)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_409),
.B(n_411),
.Y(n_443)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_411),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_412),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_411),
.A2(n_443),
.B(n_446),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_420),
.C(n_423),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_415),
.B(n_417),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_420),
.A2(n_421),
.B1(n_423),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_423),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_426),
.B(n_429),
.C(n_441),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_441),
.B2(n_442),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_437),
.B(n_440),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_438),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_440),
.B(n_494),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_492),
.C(n_494),
.Y(n_514)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_464),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_464),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_457),
.C(n_458),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_454),
.B1(n_457),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_457),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_476),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.C(n_462),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_460),
.B1(n_462),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_464),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_478),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_486),
.B(n_487),
.Y(n_485)
);

NOR2x1_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_475),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_475),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.C(n_474),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_481),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_473),
.B1(n_474),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_480),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_504),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_503),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_503),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_496),
.B1(n_498),
.B2(n_502),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_495),
.A2(n_496),
.B1(n_510),
.B2(n_511),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_506),
.C(n_510),
.Y(n_522)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_498),
.Y(n_502)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_514),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_514),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_522),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_522),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_521),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule