module real_jpeg_30046_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_244;
wire n_179;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_65),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_79),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_2),
.A2(n_26),
.B1(n_33),
.B2(n_79),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_40),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_40),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_6),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_60),
.B(n_61),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_7),
.B(n_38),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_38),
.B(n_42),
.C(n_182),
.D(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_7),
.B(n_70),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_7),
.A2(n_25),
.B(n_195),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_62),
.B(n_73),
.C(n_114),
.D(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_7),
.B(n_62),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_54),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_48),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_11),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_12),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_121)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_26),
.Y(n_183)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_115),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_21),
.B(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_88),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_22),
.B(n_80),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_52),
.C(n_66),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_24),
.B(n_36),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_25),
.A2(n_34),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_25),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_25),
.A2(n_84),
.B(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_25),
.A2(n_105),
.B1(n_107),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_25),
.B(n_197),
.Y(n_210)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_29),
.B(n_99),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_31),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_33),
.A2(n_39),
.A3(n_44),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_33),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_37),
.A2(n_49),
.B(n_148),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_43),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_38),
.A2(n_61),
.A3(n_223),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_39),
.B(n_76),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_41),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_42),
.A2(n_46),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_42),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_42),
.A2(n_46),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_49),
.B(n_150),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_49),
.A2(n_148),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_49),
.B(n_99),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_59),
.B(n_99),
.C(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_57),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_58),
.B(n_95),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_64),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_72),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_69),
.B1(n_110),
.B2(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_78),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_69),
.A2(n_72),
.B(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_70),
.A2(n_73),
.B1(n_112),
.B2(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_76),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_86),
.Y(n_125)
);

INVx5_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_83),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_83),
.A2(n_210),
.B(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_88),
.A2(n_89),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.C(n_108),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_91),
.B1(n_108),
.B2(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_93),
.B(n_99),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_103),
.A2(n_106),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_107),
.A2(n_202),
.B(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B(n_113),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_135),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_134),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_174),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_160),
.B(n_173),
.Y(n_139)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_157),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_145),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.C(n_154),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_147),
.B1(n_154),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_161),
.B(n_163),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_168),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_164),
.B(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_168),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_169),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_172),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_171),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_250),
.C(n_251),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_245),
.B(n_249),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_234),
.B(n_244),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_218),
.B(n_233),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_198),
.B(n_217),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_180),
.B(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_184),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_192),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_194),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_205),
.B(n_216),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_204),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_215),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_219),
.B(n_220),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_224),
.C(n_227),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_230),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);


endmodule