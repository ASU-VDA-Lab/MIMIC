module fake_aes_9957_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
OA21x2_ASAP7_75t_L g12 ( .A1(n_0), .A2(n_10), .B(n_5), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_0), .Y(n_17) );
OR2x6_ASAP7_75t_L g18 ( .A(n_15), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_13), .B(n_1), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_15), .B(n_2), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
OAI21xp5_ASAP7_75t_L g22 ( .A1(n_17), .A2(n_14), .B(n_13), .Y(n_22) );
A2O1A1Ixp33_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_13), .B(n_14), .C(n_16), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_11), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_21), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_21), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_16), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_11), .B1(n_13), .B2(n_19), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_28), .B(n_27), .Y(n_30) );
AOI211xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_13), .B(n_12), .C(n_5), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_28), .B(n_2), .Y(n_32) );
OAI211xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_12), .B(n_6), .C(n_3), .Y(n_33) );
NOR2x1p5_ASAP7_75t_L g34 ( .A(n_30), .B(n_12), .Y(n_34) );
NOR3xp33_ASAP7_75t_L g35 ( .A(n_31), .B(n_12), .C(n_6), .Y(n_35) );
INVxp67_ASAP7_75t_SL g36 ( .A(n_34), .Y(n_36) );
XNOR2xp5_ASAP7_75t_L g37 ( .A(n_35), .B(n_12), .Y(n_37) );
AOI21xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_33), .B(n_12), .Y(n_38) );
AOI22xp33_ASAP7_75t_SL g39 ( .A1(n_38), .A2(n_36), .B1(n_37), .B2(n_8), .Y(n_39) );
endmodule