module fake_jpeg_11041_n_449 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_449);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_449;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_58),
.B(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_28),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_60),
.B(n_69),
.Y(n_136)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_64),
.B(n_85),
.Y(n_123)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_28),
.B(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_72),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_92),
.Y(n_139)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_11),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_10),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_35),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_89),
.Y(n_147)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_35),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_34),
.B(n_9),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_98),
.Y(n_149)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_101),
.B(n_103),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_32),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_37),
.B(n_0),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_111),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_37),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_108),
.Y(n_168)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_38),
.B(n_0),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_35),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_113),
.Y(n_171)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_1),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_43),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_115),
.B(n_1),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_40),
.B1(n_42),
.B2(n_31),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_118),
.A2(n_124),
.B(n_141),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_42),
.B1(n_55),
.B2(n_43),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_119),
.A2(n_153),
.B1(n_175),
.B2(n_184),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_56),
.A2(n_42),
.B1(n_53),
.B2(n_26),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_25),
.C(n_47),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_143),
.C(n_146),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_64),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_140),
.A2(n_144),
.B1(n_151),
.B2(n_158),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_56),
.A2(n_26),
.B1(n_53),
.B2(n_43),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_85),
.B(n_24),
.C(n_47),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_26),
.B1(n_53),
.B2(n_55),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_58),
.B(n_41),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_145),
.B(n_148),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_99),
.A2(n_32),
.B(n_41),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_39),
.B1(n_49),
.B2(n_50),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_91),
.A2(n_55),
.B1(n_48),
.B2(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_50),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_154),
.B(n_155),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_101),
.B(n_49),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_52),
.C(n_27),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_185),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_176),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_93),
.A2(n_48),
.B1(n_52),
.B2(n_21),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_67),
.B(n_29),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_179),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_101),
.B(n_29),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_102),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_98),
.B(n_1),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_112),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_118),
.B1(n_184),
.B2(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_3),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_194),
.B(n_195),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_4),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_90),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_196),
.B(n_207),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_144),
.A2(n_114),
.B1(n_70),
.B2(n_71),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_197),
.A2(n_209),
.B1(n_219),
.B2(n_243),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_164),
.A2(n_102),
.B1(n_62),
.B2(n_74),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_4),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_200),
.B(n_203),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_57),
.B1(n_59),
.B2(n_77),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_202),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_128),
.B(n_5),
.Y(n_203)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_5),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_205),
.B(n_206),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_80),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_133),
.B(n_22),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_136),
.A2(n_22),
.B(n_135),
.C(n_147),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_208),
.B(n_211),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_126),
.A2(n_22),
.B1(n_181),
.B2(n_187),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_210),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_22),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_135),
.A2(n_22),
.B1(n_119),
.B2(n_150),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_212),
.A2(n_239),
.B1(n_247),
.B2(n_196),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_240),
.B1(n_189),
.B2(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_214),
.B(n_224),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_141),
.B(n_153),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_216),
.A2(n_233),
.B(n_201),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_126),
.A2(n_187),
.B1(n_157),
.B2(n_134),
.Y(n_219)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_117),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_173),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_117),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_227),
.B(n_229),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_120),
.B(n_116),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_129),
.B(n_186),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_235),
.Y(n_268)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_127),
.Y(n_231)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_120),
.B(n_116),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_127),
.B(n_137),
.Y(n_233)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_150),
.B(n_174),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_121),
.Y(n_237)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_131),
.Y(n_238)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_169),
.B(n_159),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_131),
.A2(n_182),
.B1(n_174),
.B2(n_170),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_122),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_244),
.B1(n_248),
.B2(n_210),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_132),
.B(n_161),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_245),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_170),
.A2(n_182),
.B1(n_152),
.B2(n_122),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_161),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_246),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_167),
.B(n_180),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_253),
.A2(n_265),
.B1(n_288),
.B2(n_236),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_276),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_193),
.A2(n_197),
.B1(n_248),
.B2(n_188),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_274),
.B1(n_286),
.B2(n_226),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_191),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_258),
.B(n_261),
.Y(n_323)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_211),
.A3(n_215),
.B1(n_194),
.B2(n_191),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_260),
.A2(n_283),
.B(n_277),
.C(n_267),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_192),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_218),
.B1(n_193),
.B2(n_198),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_267),
.B(n_289),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_204),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_269),
.B(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_201),
.A2(n_195),
.B1(n_205),
.B2(n_235),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_221),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_219),
.A2(n_209),
.B1(n_224),
.B2(n_243),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_218),
.A2(n_240),
.B1(n_223),
.B2(n_238),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_233),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_220),
.B(n_239),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_290),
.B(n_289),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_231),
.C(n_222),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_301),
.C(n_303),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_242),
.B(n_246),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_258),
.B(n_249),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_251),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_309),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_245),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_305),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_300),
.A2(n_270),
.B1(n_261),
.B2(n_279),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_242),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_234),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_304),
.B(n_300),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_225),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_250),
.B(n_190),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_321),
.Y(n_346)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_308),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_312),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_314),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_328),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_237),
.B1(n_241),
.B2(n_244),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_322),
.B1(n_284),
.B2(n_294),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_264),
.A2(n_217),
.B(n_253),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_294),
.B(n_266),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_283),
.B(n_277),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_324),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_273),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_270),
.A2(n_252),
.B1(n_287),
.B2(n_262),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_288),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_321),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_329),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_322),
.A2(n_290),
.B1(n_287),
.B2(n_262),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_343),
.B1(n_347),
.B2(n_352),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_307),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_356),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_318),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_345),
.A2(n_350),
.B1(n_297),
.B2(n_309),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_304),
.A2(n_282),
.B1(n_271),
.B2(n_284),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_310),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_257),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_349),
.B(n_295),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_257),
.C(n_266),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_339),
.C(n_296),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_317),
.A2(n_282),
.B1(n_259),
.B2(n_263),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_285),
.B(n_263),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_353),
.B(n_325),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_369),
.Y(n_380)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

BUFx2_ASAP7_75t_SL g383 ( 
.A(n_358),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_336),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_375),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_363),
.C(n_370),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_305),
.C(n_299),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_315),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_364),
.B(n_367),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_348),
.B1(n_333),
.B2(n_335),
.Y(n_381)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_315),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_318),
.B1(n_303),
.B2(n_326),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_373),
.B1(n_345),
.B2(n_350),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_323),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_312),
.C(n_324),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_372),
.C(n_351),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_319),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_343),
.A2(n_310),
.B1(n_298),
.B2(n_306),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_353),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_377),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_356),
.B(n_311),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_340),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_394),
.B1(n_360),
.B2(n_355),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_378),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_334),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_388),
.C(n_389),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_374),
.B1(n_359),
.B2(n_375),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_340),
.C(n_346),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_341),
.B(n_302),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_338),
.C(n_354),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_392),
.C(n_395),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_338),
.C(n_354),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_365),
.A2(n_352),
.B1(n_330),
.B2(n_337),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_370),
.C(n_357),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g421 ( 
.A(n_397),
.B(n_400),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_386),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_402),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_396),
.A2(n_360),
.B1(n_368),
.B2(n_373),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_379),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_393),
.B(n_355),
.Y(n_403)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_394),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_407),
.Y(n_413)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_337),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_408),
.A2(n_390),
.B(n_383),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_409),
.A2(n_392),
.B(n_395),
.Y(n_420)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_384),
.Y(n_410)
);

BUFx24_ASAP7_75t_SL g417 ( 
.A(n_410),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_398),
.B(n_380),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_406),
.Y(n_424)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_419),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_379),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_406),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_422),
.A2(n_380),
.B(n_382),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_412),
.Y(n_423)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_414),
.C(n_388),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_415),
.A2(n_400),
.B1(n_397),
.B2(n_408),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_425),
.B(n_427),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_403),
.Y(n_426)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_421),
.A2(n_402),
.B1(n_407),
.B2(n_405),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_421),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_430),
.B(n_433),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_417),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_425),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_436),
.A2(n_423),
.B(n_429),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_437),
.A2(n_440),
.B(n_432),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_438),
.B(n_439),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_434),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_431),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_443),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_441),
.A2(n_427),
.B(n_416),
.Y(n_444)
);

A2O1A1O1Ixp25_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_328),
.B(n_331),
.C(n_313),
.D(n_316),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_446),
.A2(n_442),
.B(n_327),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_445),
.C(n_327),
.Y(n_448)
);

BUFx24_ASAP7_75t_SL g449 ( 
.A(n_448),
.Y(n_449)
);


endmodule