module fake_jpeg_29887_n_390 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_28),
.Y(n_82)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_0),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_30),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_17),
.B1(n_28),
.B2(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_93),
.B1(n_65),
.B2(n_42),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_82),
.B(n_25),
.Y(n_145)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_17),
.B1(n_34),
.B2(n_20),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_20),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_43),
.C(n_57),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_32),
.B1(n_37),
.B2(n_31),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_45),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_40),
.A2(n_37),
.B1(n_36),
.B2(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_36),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_33),
.B1(n_23),
.B2(n_2),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_33),
.B1(n_23),
.B2(n_2),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_52),
.B1(n_65),
.B2(n_40),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_33),
.B1(n_30),
.B2(n_25),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_48),
.B1(n_58),
.B2(n_47),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_76),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_110),
.Y(n_159)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_76),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx2_ASAP7_75t_SL g162 ( 
.A(n_112),
.Y(n_162)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_117),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_51),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_48),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_48),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_129),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_53),
.B(n_49),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_131),
.C(n_133),
.Y(n_160)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_30),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_103),
.B1(n_90),
.B2(n_89),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_42),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_62),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_138),
.C(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_62),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_137),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_69),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_3),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_63),
.B1(n_58),
.B2(n_30),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_144),
.B1(n_83),
.B2(n_73),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_25),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_25),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_123),
.C(n_131),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_4),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_4),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_120),
.B1(n_130),
.B2(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_169),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_90),
.B1(n_100),
.B2(n_89),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_166),
.B1(n_136),
.B2(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_173),
.Y(n_196)
);

BUFx24_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_163),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_123),
.A2(n_91),
.B1(n_102),
.B2(n_77),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_91),
.B1(n_77),
.B2(n_70),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_115),
.B(n_119),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_81),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_134),
.A2(n_73),
.B(n_81),
.C(n_79),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_188),
.A2(n_167),
.B1(n_5),
.B2(n_6),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_193),
.B(n_202),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_115),
.B1(n_129),
.B2(n_145),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_200),
.B1(n_216),
.B2(n_171),
.Y(n_231)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_192),
.B(n_114),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_127),
.B(n_117),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_160),
.A2(n_131),
.B(n_118),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_213),
.B(n_152),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_112),
.B1(n_113),
.B2(n_139),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_199),
.Y(n_228)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_133),
.B1(n_147),
.B2(n_108),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_204),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_112),
.B1(n_128),
.B2(n_79),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_143),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_138),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_132),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_210),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_151),
.B(n_112),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_126),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_110),
.B(n_107),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_126),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_164),
.Y(n_245)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_217),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_121),
.B1(n_114),
.B2(n_6),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_181),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_224),
.C(n_226),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_181),
.C(n_175),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_153),
.B1(n_148),
.B2(n_155),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_225),
.A2(n_237),
.B1(n_244),
.B2(n_188),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_174),
.C(n_148),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_249),
.B1(n_217),
.B2(n_209),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_183),
.B(n_161),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_235),
.B(n_241),
.Y(n_276)
);

OA21x2_ASAP7_75t_SL g234 ( 
.A1(n_193),
.A2(n_211),
.B(n_206),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_234),
.B(n_187),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_177),
.B1(n_154),
.B2(n_171),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_177),
.C(n_154),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_239),
.C(n_247),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_163),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_163),
.B(n_179),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_SL g242 ( 
.A(n_190),
.B(n_163),
.C(n_167),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_242),
.A2(n_197),
.B(n_215),
.C(n_203),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_179),
.B1(n_156),
.B2(n_164),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_248),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_199),
.Y(n_247)
);

OAI22x1_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_167),
.B1(n_5),
.B2(n_7),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_216),
.B1(n_185),
.B2(n_196),
.Y(n_263)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_271),
.B1(n_274),
.B2(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_213),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_281),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_200),
.B1(n_204),
.B2(n_208),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_267),
.B1(n_231),
.B2(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_275),
.B1(n_280),
.B2(n_283),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_196),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_198),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_269),
.Y(n_307)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_185),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_228),
.B(n_247),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_270),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_186),
.Y(n_273)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_184),
.B(n_220),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_184),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_279),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_191),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_223),
.B(n_4),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_9),
.Y(n_305)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_285),
.A2(n_294),
.B1(n_295),
.B2(n_303),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_225),
.B1(n_237),
.B2(n_254),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_299),
.B1(n_301),
.B2(n_275),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_239),
.C(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_304),
.C(n_11),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_250),
.B1(n_246),
.B2(n_245),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_250),
.B1(n_246),
.B2(n_242),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_302),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_224),
.B1(n_238),
.B2(n_251),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_276),
.A2(n_244),
.B1(n_241),
.B2(n_8),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_5),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_8),
.C(n_9),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_282),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_283),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_312),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_281),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_316),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_291),
.A2(n_277),
.B1(n_273),
.B2(n_275),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_315),
.A2(n_323),
.B1(n_306),
.B2(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_288),
.B(n_301),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_318),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_275),
.B(n_262),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_320),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_293),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_268),
.B1(n_266),
.B2(n_255),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_324),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_285),
.A2(n_258),
.B1(n_260),
.B2(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_259),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_259),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_328),
.B1(n_306),
.B2(n_308),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_11),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_286),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_302),
.C(n_305),
.Y(n_329)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_329),
.B(n_337),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_313),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_290),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_334),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_299),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_297),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_322),
.Y(n_346)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_311),
.B(n_293),
.CI(n_294),
.CON(n_339),
.SN(n_339)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_340),
.A2(n_320),
.B1(n_312),
.B2(n_327),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_344),
.B(n_328),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_342),
.Y(n_348)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_331),
.A2(n_313),
.B1(n_318),
.B2(n_316),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_355),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_352),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_338),
.A2(n_319),
.B(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_351),
.B(n_340),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_330),
.Y(n_353)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_353),
.Y(n_367)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_332),
.Y(n_363)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_360),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_364),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_334),
.C(n_333),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_353),
.B(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_366),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_336),
.C(n_339),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_356),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

AOI31xp33_ASAP7_75t_L g380 ( 
.A1(n_372),
.A2(n_373),
.A3(n_358),
.B(n_298),
.Y(n_380)
);

AOI32xp33_ASAP7_75t_SL g373 ( 
.A1(n_358),
.A2(n_332),
.A3(n_351),
.B1(n_347),
.B2(n_349),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_374),
.A2(n_376),
.B(n_367),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_368),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_359),
.A2(n_350),
.B(n_314),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_378),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g379 ( 
.A(n_369),
.B(n_361),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_381),
.C(n_372),
.Y(n_383)
);

OAI322xp33_ASAP7_75t_L g384 ( 
.A1(n_380),
.A2(n_373),
.A3(n_371),
.B1(n_296),
.B2(n_326),
.C1(n_329),
.C2(n_337),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_370),
.A2(n_298),
.B(n_296),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_377),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_384),
.A2(n_321),
.B1(n_12),
.B2(n_13),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_385),
.A2(n_386),
.B(n_382),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_388),
.A2(n_13),
.B(n_14),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_14),
.Y(n_390)
);


endmodule