module real_jpeg_5861_n_32 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_29, n_191, n_10, n_31, n_9, n_186, n_12, n_24, n_189, n_187, n_6, n_190, n_28, n_192, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_193, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_184, n_30, n_16, n_15, n_13, n_32);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_29;
input n_191;
input n_10;
input n_31;
input n_9;
input n_186;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_28;
input n_192;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_193;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_0),
.B(n_106),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_1),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_2),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_61),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_4),
.B(n_74),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_5),
.B(n_126),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_6),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_7),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_9),
.B(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_10),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_11),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_64),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_12),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_12),
.B(n_168),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_13),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_14),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_15),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_16),
.B(n_53),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_16),
.A2(n_50),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_17),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_19),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_20),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_21),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_23),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_23),
.B(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_24),
.B(n_110),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_28),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_83),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_30),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_30),
.B(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_179),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_42),
.B(n_177),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_36),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_41),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_176),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_44),
.B(n_50),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_49),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_49),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_50),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_175),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_163),
.B(n_172),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_143),
.B(n_157),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_78),
.B(n_131),
.C(n_140),
.Y(n_58)
);

NOR4xp25_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.C(n_69),
.D(n_73),
.Y(n_59)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_76),
.B(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_125),
.B(n_130),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_118),
.B(n_124),
.Y(n_79)
);

AO221x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_92),
.B1(n_115),
.B2(n_116),
.C(n_117),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_98),
.B(n_114),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_109),
.B(n_113),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B(n_108),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_123),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B(n_137),
.C(n_138),
.D(n_139),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.C(n_153),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_153),
.B(n_158),
.C(n_161),
.D(n_162),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_184),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_185),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_186),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_187),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_188),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_189),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_190),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_191),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_192),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_193),
.Y(n_127)
);


endmodule