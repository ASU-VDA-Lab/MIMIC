module real_jpeg_25713_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVxp67_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_0),
.B(n_26),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_0),
.B(n_63),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_42),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_28),
.Y(n_203)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_28),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_7),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_8),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_8),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_63),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_28),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_8),
.B(n_46),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_8),
.B(n_130),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_10),
.B(n_46),
.Y(n_141)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_12),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_63),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_13),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_14),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_42),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_14),
.B(n_26),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_14),
.B(n_46),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_14),
.B(n_28),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_14),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_46),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_16),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_16),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_46),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_16),
.B(n_42),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_16),
.B(n_28),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_16),
.B(n_38),
.Y(n_195)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_145),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_94),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_21),
.A2(n_22),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_49),
.C(n_58),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.C(n_40),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_24),
.B(n_229),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_24),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_27),
.CI(n_30),
.CON(n_24),
.SN(n_24)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_25),
.B(n_27),
.C(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_40),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.C(n_45),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_41),
.B(n_44),
.CI(n_45),
.CON(n_216),
.SN(n_216)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_50),
.B(n_54),
.C(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_66),
.C(n_67),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_69),
.B(n_201),
.Y(n_200)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_73),
.B(n_94),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.C(n_83),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_74),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_82),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_81),
.Y(n_82)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_96),
.C(n_97),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_83),
.B(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.C(n_92),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_84),
.A2(n_85),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_140),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_102),
.CI(n_105),
.CON(n_98),
.SN(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_143),
.B2(n_144),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_135),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_134),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_234),
.C(n_235),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_222),
.C(n_223),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_210),
.C(n_211),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_173),
.C(n_184),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_163),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_158),
.C(n_163),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_153),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_161),
.C(n_162),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_171),
.C(n_172),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_183),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_178),
.B1(n_183),
.B2(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_206),
.C(n_207),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.C(n_198),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_191),
.C(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_218),
.C(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_216),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.C(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);


endmodule