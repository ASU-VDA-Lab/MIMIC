module fake_jpeg_14789_n_62 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_7),
.B(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_40),
.C(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_10),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_6),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_26),
.B(n_13),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_12),
.B1(n_23),
.B2(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_53),
.B1(n_48),
.B2(n_15),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_49),
.C(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_45),
.B1(n_54),
.B2(n_43),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_54),
.B(n_17),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_11),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);


endmodule