module fake_jpeg_5216_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_44),
.B1(n_56),
.B2(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_59),
.B1(n_45),
.B2(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_51),
.B1(n_62),
.B2(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_63),
.B1(n_55),
.B2(n_12),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_52),
.B1(n_46),
.B2(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_81),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_82)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_79),
.Y(n_85)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_76),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_73),
.B(n_74),
.C(n_15),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_86),
.B(n_90),
.C(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_92),
.B(n_95),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_94),
.B1(n_10),
.B2(n_17),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_9),
.B(n_18),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_20),
.C(n_21),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_22),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_23),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_24),
.B(n_26),
.C(n_34),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_37),
.C(n_39),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_42),
.Y(n_107)
);


endmodule