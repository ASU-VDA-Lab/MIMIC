module fake_jpeg_12078_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_35),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_5),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_12),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_3),
.Y(n_96)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_49),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_69),
.B1(n_65),
.B2(n_62),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_94),
.B1(n_78),
.B2(n_74),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_91),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_69),
.B1(n_59),
.B2(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_49),
.B1(n_53),
.B2(n_63),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_84),
.B(n_98),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_55),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_102),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_50),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_53),
.B1(n_63),
.B2(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_116),
.B1(n_118),
.B2(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_55),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_6),
.B(n_8),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_48),
.B(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_117),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_53),
.B1(n_66),
.B2(n_64),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_70),
.C(n_26),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_138),
.C(n_31),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_3),
.C(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_126),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_6),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_136),
.B1(n_125),
.B2(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_21),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_13),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_28),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_23),
.B(n_27),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_29),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_126),
.B(n_139),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_154),
.C(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_141),
.B1(n_147),
.B2(n_144),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_138),
.C(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_121),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_159),
.A3(n_155),
.B1(n_161),
.B2(n_134),
.C1(n_40),
.C2(n_41),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_159),
.C(n_167),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_134),
.CI(n_33),
.CON(n_170),
.SN(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_32),
.C(n_34),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_172)
);


endmodule