module fake_jpeg_6244_n_289 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_14),
.B1(n_24),
.B2(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_13),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_46),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_16),
.B1(n_22),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_14),
.B1(n_32),
.B2(n_31),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_37),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_14),
.B1(n_24),
.B2(n_17),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_34),
.B1(n_28),
.B2(n_37),
.Y(n_71)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_75),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_67),
.B1(n_77),
.B2(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_54),
.B1(n_45),
.B2(n_50),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_81),
.B1(n_29),
.B2(n_18),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_28),
.B1(n_22),
.B2(n_29),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_22),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_62),
.C(n_20),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_38),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_40),
.B1(n_32),
.B2(n_35),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_42),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_30),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_70),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_102),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_30),
.C(n_17),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_63),
.Y(n_112)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_102),
.B1(n_87),
.B2(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_65),
.B1(n_66),
.B2(n_64),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_118),
.B1(n_97),
.B2(n_93),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_71),
.B(n_80),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_128),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_71),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_122),
.B(n_20),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_64),
.C(n_80),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_113),
.C(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_121),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_68),
.C(n_78),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_125),
.B1(n_91),
.B2(n_85),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_41),
.B1(n_51),
.B2(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_81),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_27),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_52),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_59),
.B1(n_68),
.B2(n_79),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_78),
.C(n_53),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_46),
.B1(n_79),
.B2(n_93),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_118),
.B1(n_79),
.B2(n_59),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_149),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_123),
.C(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_122),
.B(n_23),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_89),
.Y(n_154)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_109),
.B(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_124),
.B(n_127),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_165),
.B(n_173),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_124),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_161),
.C(n_171),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_107),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_15),
.B(n_21),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_146),
.B1(n_143),
.B2(n_136),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_101),
.B1(n_116),
.B2(n_47),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_172),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_137),
.C(n_152),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_47),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_134),
.B1(n_132),
.B2(n_138),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_58),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_115),
.C(n_15),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_192),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_133),
.C(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_141),
.B1(n_145),
.B2(n_140),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_195),
.B(n_205),
.C(n_167),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_104),
.B1(n_129),
.B2(n_101),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_15),
.C(n_17),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_96),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_20),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_72),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_101),
.B1(n_116),
.B2(n_115),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_199),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_202),
.C(n_163),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_201),
.B1(n_179),
.B2(n_163),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_21),
.B1(n_23),
.B2(n_52),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_161),
.C(n_171),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_52),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_175),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_216),
.C(n_223),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_177),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_204),
.Y(n_228)
);

AO221x1_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_156),
.B1(n_203),
.B2(n_198),
.C(n_98),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_157),
.C(n_162),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_162),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_26),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_175),
.B(n_165),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_220),
.B(n_57),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_169),
.B(n_168),
.C(n_157),
.D(n_164),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_8),
.Y(n_245)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_156),
.C(n_160),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_25),
.C(n_26),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_23),
.B1(n_21),
.B2(n_72),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_196),
.B1(n_194),
.B2(n_186),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_186),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_210),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_200),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_241),
.B(n_244),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_209),
.B1(n_187),
.B2(n_212),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_234),
.B1(n_207),
.B2(n_221),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_197),
.B1(n_201),
.B2(n_191),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_242),
.C(n_223),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_26),
.CI(n_1),
.CON(n_237),
.SN(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_206),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_0),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_245),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_98),
.B(n_83),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_105),
.C(n_83),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_233),
.C(n_228),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_222),
.C(n_225),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_8),
.B(n_13),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_214),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_253),
.B(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_208),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_210),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_237),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_236),
.B1(n_232),
.B2(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_69),
.C(n_1),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_240),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_234),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_264),
.B(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_246),
.B(n_240),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_270),
.C(n_12),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_239),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_237),
.C(n_238),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_267),
.A2(n_246),
.B1(n_256),
.B2(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.C(n_276),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_247),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_277),
.A2(n_9),
.B(n_2),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_273),
.C2(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_280),
.B(n_282),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_275),
.C2(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_6),
.Y(n_287)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_281),
.B(n_5),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_287),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_285),
.Y(n_289)
);


endmodule