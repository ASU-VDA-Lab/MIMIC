module real_jpeg_11536_n_20 (n_17, n_8, n_0, n_93, n_2, n_91, n_10, n_9, n_12, n_92, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_93;
input n_2;
input n_91;
input n_10;
input n_9;
input n_12;
input n_92;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_0),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI221xp5_ASAP7_75t_L g40 ( 
.A1(n_0),
.A2(n_8),
.B1(n_28),
.B2(n_41),
.C(n_42),
.Y(n_40)
);

AOI221xp5_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_1),
.B1(n_28),
.B2(n_43),
.C(n_44),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_18),
.B1(n_28),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_4),
.B1(n_28),
.B2(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_0),
.B(n_9),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_0),
.A2(n_49),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_91),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_52),
.B1(n_58),
.B2(n_69),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_9),
.B(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_9),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_10),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_12),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_92),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_93),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_22),
.B1(n_23),
.B2(n_50),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_19),
.A2(n_50),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_51),
.B1(n_76),
.B2(n_79),
.C(n_88),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR5xp2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.C(n_46),
.D(n_47),
.E(n_49),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_34),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_31),
.C(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_33),
.Y(n_85)
);

NOR5xp2_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_40),
.C(n_47),
.D(n_82),
.E(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_37),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_70),
.B(n_74),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_75),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_60),
.B(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B(n_68),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_85),
.Y(n_87)
);


endmodule