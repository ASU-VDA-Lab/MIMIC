module real_jpeg_13117_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_2),
.A2(n_46),
.B1(n_60),
.B2(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_2),
.A2(n_29),
.B1(n_36),
.B2(n_46),
.Y(n_144)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_4),
.A2(n_53),
.B1(n_60),
.B2(n_64),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_60),
.B1(n_64),
.B2(n_71),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_71),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_71),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_8),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_8),
.A2(n_60),
.B1(n_64),
.B2(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_103),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_103),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_69),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_60),
.B1(n_64),
.B2(n_69),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_69),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_12),
.A2(n_60),
.B1(n_64),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_80),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_80),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_13),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_13),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_13),
.A2(n_66),
.B(n_163),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_154),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_13),
.A2(n_44),
.B(n_49),
.C(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_13),
.B(n_110),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_13),
.B(n_33),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_13),
.B(n_54),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_64),
.B(n_74),
.C(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_14),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_14),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_15),
.A2(n_60),
.B1(n_64),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_15),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_15),
.A2(n_66),
.B1(n_67),
.B2(n_136),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_136),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_136),
.Y(n_210)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_104),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_22),
.B(n_104),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_88),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_23),
.B(n_82),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_57),
.C(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_28),
.A2(n_33),
.B(n_38),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_28),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_28),
.A2(n_33),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_28),
.A2(n_33),
.B1(n_143),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_28),
.A2(n_33),
.B1(n_94),
.B2(n_144),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_28),
.A2(n_33),
.B1(n_157),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_28),
.A2(n_33),
.B1(n_154),
.B2(n_210),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_28),
.A2(n_33),
.B1(n_203),
.B2(n_210),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_29),
.B(n_212),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_32),
.A2(n_35),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_32),
.A2(n_92),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_36),
.A2(n_50),
.B(n_154),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_43),
.A2(n_51),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_45),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_44),
.B(n_77),
.Y(n_155)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_45),
.A2(n_64),
.A3(n_76),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_47),
.A2(n_54),
.B1(n_86),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_47),
.A2(n_54),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_54),
.B1(n_97),
.B2(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_47),
.A2(n_54),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_47),
.A2(n_54),
.B1(n_189),
.B2(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_51),
.A2(n_98),
.B1(n_147),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_72),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_58),
.A2(n_59),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_60),
.B(n_154),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_60),
.A2(n_63),
.A3(n_66),
.B1(n_164),
.B2(n_178),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_62),
.B(n_64),
.Y(n_178)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_67),
.B(n_154),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_73),
.A2(n_78),
.B1(n_138),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_74),
.A2(n_110),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_74),
.A2(n_110),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_78),
.A2(n_135),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_84),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_85),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_88),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.C(n_101),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_89),
.A2(n_90),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_91),
.B(n_95),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_99),
.B(n_101),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_100),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_102),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_124),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_113),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_267),
.B(n_271),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_254),
.B(n_255),
.C(n_266),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_238),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_181),
.B(n_237),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_158),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_131),
.B(n_158),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_145),
.C(n_149),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_132),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_140),
.C(n_142),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_141),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_172),
.B2(n_180),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_159),
.B(n_173),
.C(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_161),
.B(n_167),
.C(n_171),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_179),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_174),
.B(n_177),
.Y(n_253)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_231),
.B(n_236),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_219),
.B(n_230),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_199),
.B(n_218),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_185),
.B(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_195),
.C(n_197),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_207),
.B(n_217),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_205),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_213),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_221),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_240),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_243),
.C(n_244),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_249),
.C(n_253),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_264),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);


endmodule