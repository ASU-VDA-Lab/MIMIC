module fake_jpeg_29016_n_341 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_341);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_45),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_0),
.B(n_1),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_2),
.C(n_4),
.Y(n_74)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_51),
.B(n_41),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_57),
.Y(n_78)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_84),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_25),
.B1(n_43),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_96),
.B1(n_98),
.B2(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_31),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_30),
.B1(n_42),
.B2(n_40),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_85),
.A2(n_93),
.B1(n_108),
.B2(n_6),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_91),
.B(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_95),
.B(n_103),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_59),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_70),
.B(n_39),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_38),
.B1(n_44),
.B2(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_35),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_6),
.Y(n_152)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_28),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_78),
.B(n_10),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_53),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_21),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_142),
.C(n_156),
.Y(n_181)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_144),
.Y(n_172)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_28),
.B1(n_26),
.B2(n_21),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_88),
.A2(n_26),
.B1(n_65),
.B2(n_66),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_143),
.B1(n_90),
.B2(n_87),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_89),
.B(n_69),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_88),
.A2(n_64),
.B1(n_68),
.B2(n_49),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_82),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_152),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_99),
.B1(n_108),
.B2(n_77),
.Y(n_159)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_154),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_73),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_7),
.C(n_8),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_163),
.B1(n_167),
.B2(n_169),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_159),
.A2(n_161),
.B1(n_164),
.B2(n_128),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_99),
.B1(n_112),
.B2(n_75),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_112),
.B1(n_76),
.B2(n_75),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_76),
.B1(n_106),
.B2(n_111),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_165),
.A2(n_180),
.B(n_184),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_111),
.B1(n_114),
.B2(n_11),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_114),
.B1(n_10),
.B2(n_11),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_182),
.B1(n_185),
.B2(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_9),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_17),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_156),
.Y(n_193)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_12),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_177),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_130),
.B(n_15),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_15),
.B1(n_16),
.B2(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_142),
.B1(n_126),
.B2(n_124),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_186),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_195),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_118),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_142),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_208),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_210),
.B1(n_191),
.B2(n_170),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_120),
.B(n_147),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_220),
.B(n_159),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_132),
.C(n_138),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_153),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_146),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_131),
.B1(n_134),
.B2(n_137),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_131),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_178),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_221),
.B(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_181),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_214),
.A2(n_159),
.B(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_159),
.B(n_157),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_181),
.B(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_183),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_224),
.B(n_227),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_187),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_240),
.C(n_211),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_243),
.B(n_249),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_157),
.B(n_187),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_201),
.B1(n_218),
.B2(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_250),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_206),
.A2(n_191),
.B(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_245),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_243),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_200),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_261),
.C(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_264),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_205),
.B1(n_220),
.B2(n_217),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_271),
.B(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_207),
.C(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_207),
.C(n_193),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_199),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_270),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_210),
.B1(n_201),
.B2(n_223),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_244),
.B1(n_223),
.B2(n_238),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_214),
.C(n_204),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_232),
.C(n_247),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_194),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_227),
.A2(n_208),
.B(n_222),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_224),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_279),
.C(n_281),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_268),
.B(n_259),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_265),
.B1(n_258),
.B2(n_228),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_196),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_221),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_231),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.C(n_289),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_231),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_196),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_189),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_233),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_271),
.B(n_272),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_293),
.A2(n_294),
.B(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_267),
.B1(n_262),
.B2(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_277),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_268),
.B1(n_260),
.B2(n_262),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_234),
.B1(n_230),
.B2(n_239),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_260),
.C(n_258),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_285),
.C(n_279),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_281),
.B1(n_232),
.B2(n_228),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_233),
.B(n_246),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_306),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_283),
.Y(n_305)
);

XOR2x2_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_303),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_307),
.B(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_280),
.C(n_289),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_290),
.C(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_323),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_293),
.B(n_298),
.C(n_294),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_297),
.B(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_295),
.B(n_291),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_306),
.B(n_310),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_318),
.A2(n_301),
.B(n_314),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_311),
.C(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_282),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_329),
.B(n_324),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_322),
.C(n_320),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_327),
.C(n_324),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_316),
.B(n_311),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_304),
.B(n_234),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_230),
.B(n_250),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_337),
.B(n_216),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_336),
.Y(n_341)
);


endmodule