module real_jpeg_13743_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_3),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_3),
.B(n_34),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_26),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_45),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_28),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_5),
.B(n_34),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_41),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_6),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_45),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_6),
.B(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_7),
.B(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_7),
.B(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_41),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_7),
.B(n_70),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_10),
.B(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_10),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_10),
.B(n_28),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_11),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_11),
.B(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_11),
.B(n_62),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_11),
.B(n_41),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_13),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_13),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_45),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_28),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_13),
.B(n_34),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_13),
.B(n_62),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_13),
.B(n_41),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_14),
.B(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_41),
.Y(n_132)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_19),
.B(n_111),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.C(n_98),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_20),
.B(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_57),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_22),
.B(n_36),
.C(n_57),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_27),
.B(n_30),
.C(n_33),
.Y(n_122)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_47),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_39),
.B(n_43),
.C(n_47),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_40),
.B(n_56),
.Y(n_212)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.C(n_52),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_52),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_56),
.B(n_63),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.C(n_71),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_58),
.A2(n_59),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_59),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_61),
.CI(n_65),
.CON(n_59),
.SN(n_59)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_61),
.C(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_63),
.B(n_95),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_66),
.B(n_71),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_67),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.C(n_77),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_74),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_75),
.B(n_95),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_76),
.B(n_91),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_77),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_78),
.A2(n_79),
.B1(n_98),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_88),
.C(n_97),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_83),
.C(n_86),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_83),
.A2(n_85),
.B1(n_105),
.B2(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_97),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_90),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_91),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.C(n_110),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_102),
.CI(n_110),
.CON(n_147),
.SN(n_147)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.C(n_108),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_103),
.A2(n_104),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_105),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_140),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_124),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_139),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_138),
.B(n_181),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_167),
.B(n_248),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_164),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_145),
.B(n_164),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_152),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_146),
.A2(n_147),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_147),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_246)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_158),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_154),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_157),
.B(n_158),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_162),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_242),
.B(n_247),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_227),
.B(n_241),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_197),
.B(n_226),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_183),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_171),
.B(n_183),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_180),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_223),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.CI(n_175),
.CON(n_172),
.SN(n_172)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_196),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_189),
.C(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_193),
.C(n_194),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_220),
.B(n_225),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_210),
.B(n_219),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_208),
.C(n_209),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_214),
.B(n_218),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_229),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_235),
.C(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);


endmodule