module real_jpeg_11677_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_45),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_3),
.B(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_3),
.B(n_72),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_3),
.B(n_76),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_4),
.B(n_45),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_4),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_4),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_76),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_7),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_7),
.B(n_53),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_8),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_8),
.B(n_30),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_45),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_8),
.B(n_62),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_8),
.B(n_26),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_12),
.B(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_13),
.B(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_30),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_45),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_13),
.B(n_62),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_13),
.B(n_26),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_13),
.B(n_72),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_13),
.B(n_76),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_13),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_14),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_14),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_62),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_14),
.B(n_76),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_14),
.B(n_53),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_26),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_53),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_15),
.B(n_30),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_169),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_167),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_19),
.B(n_130),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.C(n_100),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_20),
.B(n_85),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_64),
.B2(n_65),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_21),
.B(n_66),
.C(n_78),
.Y(n_166)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_41),
.C(n_58),
.Y(n_134)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_25),
.B(n_29),
.C(n_32),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g187 ( 
.A(n_26),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_33),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_33),
.B(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_37),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_37),
.B(n_121),
.Y(n_258)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_56),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_44),
.B(n_52),
.C(n_54),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_45),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_48),
.A2(n_54),
.B1(n_107),
.B2(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_50),
.B(n_109),
.Y(n_290)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_68),
.C(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_52),
.A2(n_55),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_52),
.B(n_260),
.Y(n_270)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_107),
.C(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_61),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_63),
.B(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_75),
.C(n_77),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_70),
.A2(n_71),
.B1(n_181),
.B2(n_182),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_71),
.B(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_73),
.B(n_125),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_73),
.B(n_109),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_77),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_83),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_82),
.A2(n_83),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_82),
.A2(n_83),
.B1(n_97),
.B2(n_117),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_83),
.B(n_97),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.C(n_95),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_86),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_90),
.B(n_95),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.C(n_94),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_93),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_93),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_93),
.A2(n_163),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_94),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.C(n_98),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_100),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_114),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_105),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_108),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_114),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_126),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_115),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_119),
.A2(n_120),
.B(n_123),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_121),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_125),
.B(n_187),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_126),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.C(n_129),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_128),
.CI(n_129),
.CON(n_179),
.SN(n_179)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_166),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_146),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_144),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_155),
.B2(n_156),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_165),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_161),
.A2(n_162),
.B1(n_184),
.B2(n_185),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_184),
.C(n_186),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_197),
.B(n_328),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_195),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_171),
.B(n_195),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_174),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_188),
.C(n_191),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_183),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_178),
.A2(n_179),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_179),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_180),
.B(n_183),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_186),
.B(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_245),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_222),
.B(n_244),
.Y(n_199)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_200),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_220),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_220),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_208),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.C(n_219),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_212),
.CI(n_219),
.CON(n_228),
.SN(n_228)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_217),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_213),
.A2(n_214),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_223),
.B(n_226),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_233),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_227),
.A2(n_228),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_228),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.Y(n_324)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_238),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_235),
.B(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_237),
.B(n_238),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_326),
.C(n_327),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_320),
.B(n_325),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_305),
.B(n_319),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_275),
.B(n_304),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_262),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_250),
.B(n_262),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.C(n_259),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_301),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.CI(n_254),
.CON(n_251),
.SN(n_251)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_257),
.B(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_274),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_268),
.C(n_274),
.Y(n_306)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_298),
.B(n_303),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_288),
.B(n_297),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_292),
.B(n_296),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_306),
.B(n_307),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_313),
.C(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);


endmodule