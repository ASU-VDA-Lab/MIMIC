module fake_jpeg_25317_n_221 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_221);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_10),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_10),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_14),
.B(n_17),
.C(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_11),
.Y(n_52)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_30),
.B1(n_18),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_50),
.B1(n_11),
.B2(n_15),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_54),
.B1(n_36),
.B2(n_18),
.Y(n_59)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_47),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_57),
.B1(n_36),
.B2(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_24),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_29),
.B(n_16),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_23),
.B1(n_22),
.B2(n_31),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_11),
.B1(n_21),
.B2(n_16),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_61),
.B1(n_65),
.B2(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_62),
.B1(n_44),
.B2(n_41),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_57),
.B1(n_43),
.B2(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_66),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_9),
.C(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_12),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_21),
.B1(n_15),
.B2(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_64),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_58),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_43),
.B1(n_46),
.B2(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_62),
.B1(n_60),
.B2(n_74),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_50),
.B(n_55),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_95),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_22),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_51),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_44),
.B1(n_41),
.B2(n_51),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_76),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_106),
.Y(n_137)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_109),
.B(n_111),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_68),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_61),
.Y(n_109)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_83),
.B1(n_38),
.B2(n_37),
.Y(n_135)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_85),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

NAND2x1_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

INVxp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_97),
.B1(n_51),
.B2(n_82),
.Y(n_133)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_126),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_84),
.CI(n_79),
.CON(n_126),
.SN(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_84),
.B1(n_80),
.B2(n_87),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_79),
.C(n_87),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_88),
.C(n_84),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_145),
.B1(n_100),
.B2(n_119),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_101),
.C(n_106),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_146),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_37),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_118),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_38),
.B1(n_2),
.B2(n_3),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_114),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_38),
.B1(n_0),
.B2(n_4),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_100),
.B1(n_109),
.B2(n_102),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_4),
.C(n_5),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_134),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_156),
.B(n_157),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_115),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_129),
.B(n_117),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_172),
.B(n_140),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_158),
.B(n_152),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_138),
.C(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_149),
.C(n_154),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_135),
.B1(n_142),
.B2(n_122),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_150),
.B1(n_107),
.B2(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_157),
.B1(n_151),
.B2(n_126),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_185),
.B(n_188),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_129),
.B(n_107),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_154),
.C(n_98),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_176),
.C(n_134),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_166),
.B(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_173),
.C(n_143),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_165),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_194),
.C(n_177),
.Y(n_202)
);

AO221x1_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_123),
.B1(n_168),
.B2(n_167),
.C(n_178),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_112),
.B(n_4),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_169),
.C(n_146),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_186),
.C(n_98),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_198),
.A2(n_187),
.B(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_181),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_202),
.C(n_205),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_204),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_7),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_190),
.CI(n_195),
.CON(n_206),
.SN(n_206)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_7),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_192),
.C(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_211),
.B(n_0),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_9),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_213),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_0),
.A3(n_206),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_216),
.C(n_214),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_210),
.B(n_209),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_0),
.Y(n_221)
);


endmodule