module fake_jpeg_29127_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_0),
.B(n_1),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_3),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_46),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_48),
.B1(n_44),
.B2(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_82)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_38),
.C(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_35),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_23),
.C(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_22),
.C(n_34),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_96),
.B(n_11),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_12),
.B1(n_15),
.B2(n_18),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_9),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_76),
.B1(n_84),
.B2(n_16),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_101),
.B1(n_96),
.B2(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_86),
.C(n_97),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_102),
.B(n_92),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.C(n_106),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_107),
.B1(n_104),
.B2(n_90),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_19),
.A3(n_24),
.B1(n_27),
.B2(n_28),
.C1(n_30),
.C2(n_31),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_33),
.Y(n_114)
);


endmodule