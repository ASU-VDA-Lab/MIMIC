module fake_jpeg_6946_n_328 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_23),
.B1(n_22),
.B2(n_16),
.Y(n_45)
);

CKINVDCx9p33_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_16),
.B1(n_21),
.B2(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_35),
.B(n_18),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_43),
.B(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_33),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_22),
.B1(n_23),
.B2(n_46),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_81),
.B1(n_85),
.B2(n_93),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_39),
.C(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_22),
.B1(n_23),
.B2(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_47),
.B1(n_55),
.B2(n_39),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_40),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_100),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_35),
.B1(n_17),
.B2(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_37),
.B1(n_33),
.B2(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_107),
.Y(n_130)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_34),
.B(n_29),
.C(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_81),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_121),
.Y(n_144)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_21),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_123),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_84),
.C(n_92),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_145),
.C(n_110),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_83),
.B1(n_89),
.B2(n_92),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_132),
.B1(n_140),
.B2(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_131),
.Y(n_151)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_89),
.B1(n_84),
.B2(n_79),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_95),
.B(n_80),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_149),
.C(n_121),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_141),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_85),
.B1(n_61),
.B2(n_65),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_86),
.B1(n_93),
.B2(n_61),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_26),
.B(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_155),
.C(n_125),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_118),
.C(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_111),
.B1(n_107),
.B2(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_135),
.B1(n_107),
.B2(n_87),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_170),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_108),
.B(n_122),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_162),
.B(n_19),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_122),
.B1(n_108),
.B2(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_99),
.B1(n_19),
.B2(n_32),
.Y(n_201)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_146),
.B1(n_128),
.B2(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_177),
.B(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_147),
.B1(n_82),
.B2(n_26),
.Y(n_187)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_182),
.C(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_138),
.C(n_144),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_147),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_64),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_58),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_87),
.B1(n_91),
.B2(n_58),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_91),
.B1(n_58),
.B2(n_99),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_50),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_201),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_36),
.C(n_37),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_159),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_99),
.B1(n_19),
.B2(n_37),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_202),
.B1(n_152),
.B2(n_165),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_161),
.C(n_158),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_177),
.B1(n_156),
.B2(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_75),
.C(n_74),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_24),
.C(n_32),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_167),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_215),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_214),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_212),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_151),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_169),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_24),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_11),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_66),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_11),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_221),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_63),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_226),
.B1(n_200),
.B2(n_180),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_0),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_205),
.C(n_203),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_187),
.B1(n_14),
.B2(n_32),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_205),
.B1(n_193),
.B2(n_191),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_215),
.C(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_188),
.B1(n_196),
.B2(n_193),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_212),
.B1(n_14),
.B2(n_24),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_182),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_227),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_225),
.B(n_224),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_211),
.B(n_217),
.C(n_208),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_247),
.A2(n_211),
.B(n_217),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_75),
.B1(n_74),
.B2(n_59),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_211),
.A2(n_207),
.B1(n_225),
.B2(n_206),
.Y(n_249)
);

XOR2x1_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_0),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_252),
.B(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_262),
.B(n_264),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_260),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_232),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_265),
.B(n_267),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_0),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_27),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_14),
.B1(n_24),
.B2(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_249),
.C(n_239),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_27),
.CI(n_1),
.CON(n_266),
.SN(n_266)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_241),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_242),
.C(n_233),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_272),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_233),
.B(n_251),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_258),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_244),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_244),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_275),
.C(n_280),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_231),
.B1(n_246),
.B2(n_12),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_278),
.B1(n_273),
.B2(n_270),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_64),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_283),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g278 ( 
.A(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_27),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_264),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_285),
.B(n_290),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_262),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_250),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_266),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_4),
.Y(n_304)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_271),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_303),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.C(n_305),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_2),
.C(n_3),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_304),
.B1(n_5),
.B2(n_6),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_3),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_4),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_301),
.A2(n_297),
.B1(n_298),
.B2(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_286),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_5),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_313),
.C(n_6),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_7),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_6),
.B(n_7),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_315),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_314),
.B(n_8),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_320),
.A2(n_321),
.B(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_316),
.Y(n_323)
);

AO21x1_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_7),
.B(n_9),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_9),
.B(n_10),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_10),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_10),
.Y(n_328)
);


endmodule