module fake_jpeg_22979_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_41)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.Y(n_49)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_52),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_30),
.B1(n_16),
.B2(n_20),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_50),
.A3(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_30),
.B1(n_16),
.B2(n_24),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_25),
.B1(n_18),
.B2(n_20),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_15),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_29),
.B1(n_17),
.B2(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_66),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_55),
.B(n_49),
.C(n_56),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_1),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_1),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_52),
.A3(n_47),
.B1(n_13),
.B2(n_9),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_1),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_46),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_3),
.C(n_4),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_41),
.B1(n_48),
.B2(n_43),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_89),
.B1(n_58),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_41),
.B1(n_44),
.B2(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_87),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_54),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_62),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_99),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_67),
.C(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_104),
.B(n_78),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVxp33_ASAP7_75t_SL g125 ( 
.A(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_78),
.B1(n_77),
.B2(n_80),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_98),
.B1(n_97),
.B2(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_115),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_82),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_60),
.C(n_69),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_124),
.C(n_87),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_68),
.B(n_48),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_90),
.B(n_73),
.C(n_59),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_101),
.B1(n_95),
.B2(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_92),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_108),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_116),
.C(n_112),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_120),
.CI(n_113),
.CON(n_138),
.SN(n_138)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_45),
.B1(n_76),
.B2(n_60),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_123),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_76),
.B1(n_47),
.B2(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_118),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_130),
.B(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_135),
.B(n_132),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_115),
.C(n_124),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.C(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_79),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_133),
.CI(n_130),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_135),
.B(n_111),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_140),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_159),
.A2(n_160),
.B(n_4),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_145),
.B1(n_150),
.B2(n_152),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_13),
.C(n_14),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_154),
.B(n_150),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_166),
.B(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

OAI221xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_138),
.B1(n_154),
.B2(n_12),
.C(n_10),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.C(n_6),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_14),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_171),
.B(n_6),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_7),
.Y(n_173)
);


endmodule