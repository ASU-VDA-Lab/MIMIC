module fake_jpeg_23680_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_49),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_16),
.B1(n_23),
.B2(n_22),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_47),
.B1(n_30),
.B2(n_34),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_23),
.B1(n_19),
.B2(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_20),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_23),
.B(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_63),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_37),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_16),
.B1(n_21),
.B2(n_33),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_16),
.B1(n_21),
.B2(n_26),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_79),
.B1(n_80),
.B2(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_37),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_36),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_77),
.C(n_78),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_87),
.B1(n_44),
.B2(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_83),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_89),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_17),
.B(n_25),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_44),
.A2(n_24),
.B1(n_18),
.B2(n_17),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_32),
.B1(n_28),
.B2(n_20),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_66),
.B1(n_69),
.B2(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_68),
.B1(n_25),
.B2(n_17),
.Y(n_141)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_56),
.B(n_45),
.C(n_18),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_84),
.B1(n_82),
.B2(n_87),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_45),
.B1(n_56),
.B2(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_103),
.B1(n_70),
.B2(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_51),
.B1(n_24),
.B2(n_18),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_51),
.C(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_114),
.Y(n_125)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_117),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_27),
.C(n_24),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_71),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_63),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_98),
.B1(n_126),
.B2(n_101),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_118),
.A2(n_70),
.B1(n_89),
.B2(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_123),
.B1(n_140),
.B2(n_141),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_61),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_137),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_61),
.B(n_58),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_132),
.B(n_99),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_61),
.B(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_18),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_138),
.Y(n_149)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_27),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_81),
.B1(n_62),
.B2(n_68),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_25),
.B1(n_68),
.B2(n_2),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_102),
.B1(n_112),
.B2(n_96),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_0),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_106),
.Y(n_157)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_9),
.B(n_14),
.C(n_13),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_103),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_167),
.B1(n_128),
.B2(n_139),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_99),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_169),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_98),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_170),
.C(n_122),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_112),
.B(n_101),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_160),
.B(n_122),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_171),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_119),
.B(n_122),
.C(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_166),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_109),
.B1(n_101),
.B2(n_111),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_172),
.B1(n_142),
.B2(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_98),
.B1(n_94),
.B2(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_175),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_107),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_100),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_98),
.B1(n_114),
.B2(n_108),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_108),
.C(n_104),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_178),
.B1(n_198),
.B2(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_125),
.B1(n_119),
.B2(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_181),
.B(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_188),
.B1(n_192),
.B2(n_199),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_197),
.C(n_170),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_191),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_137),
.B1(n_134),
.B2(n_3),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_134),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_179),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_9),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_150),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_210),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_199),
.B1(n_149),
.B2(n_198),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_156),
.C(n_175),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_165),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_147),
.B(n_162),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_183),
.B(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_174),
.B1(n_162),
.B2(n_147),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_215),
.B1(n_177),
.B2(n_178),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_169),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_197),
.C(n_196),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_162),
.B1(n_168),
.B2(n_163),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_233),
.B(n_208),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_229),
.B1(n_231),
.B2(n_12),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_184),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_200),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_211),
.C(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_187),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_157),
.C(n_149),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_230),
.C(n_201),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_166),
.C(n_152),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_11),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_204),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_245),
.C(n_246),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_207),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_242),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_205),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_222),
.B1(n_234),
.B2(n_231),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_208),
.C(n_11),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_1),
.C(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_219),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_251),
.B(n_10),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_222),
.C(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_232),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_246),
.CI(n_224),
.CON(n_262),
.SN(n_262)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_260),
.B(n_262),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_244),
.B1(n_221),
.B2(n_237),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_249),
.B1(n_256),
.B2(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_242),
.B1(n_238),
.B2(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_256),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_264),
.A2(n_249),
.B(n_15),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_10),
.B(n_13),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_250),
.A3(n_14),
.B1(n_15),
.B2(n_10),
.C1(n_13),
.C2(n_5),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_269),
.B(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_262),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_258),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_274),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_262),
.B(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_270),
.Y(n_276)
);

AOI31xp33_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_273),
.A3(n_6),
.B(n_7),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_6),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_277),
.B(n_6),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_7),
.Y(n_281)
);


endmodule