module fake_jpeg_32_n_221 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_13),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_16),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_1),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_68),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_73),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_57),
.B1(n_73),
.B2(n_63),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_105)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_77),
.B1(n_57),
.B2(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_80),
.B1(n_71),
.B2(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_77),
.B1(n_63),
.B2(n_62),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_88),
.B1(n_87),
.B2(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_76),
.B1(n_97),
.B2(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_70),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_117),
.B1(n_76),
.B2(n_64),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_1),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_69),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_141),
.B1(n_105),
.B2(n_114),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_60),
.C(n_61),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_143),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_79),
.B(n_75),
.C(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_140),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_94),
.B(n_78),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_2),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_146),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_155),
.B1(n_157),
.B2(n_151),
.Y(n_172)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_2),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_154),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_78),
.B1(n_4),
.B2(n_6),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_3),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_164),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_78),
.B1(n_6),
.B2(n_7),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_30),
.C(n_52),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_166),
.C(n_31),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_131),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_167),
.B(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_29),
.C(n_51),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_152),
.B(n_145),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_171),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_158),
.B(n_163),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_175),
.B1(n_186),
.B2(n_11),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_4),
.B(n_7),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_174),
.Y(n_190)
);

AO21x2_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_54),
.B(n_26),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_50),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.C(n_173),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_25),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_23),
.B(n_47),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_22),
.B(n_46),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_192),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_195),
.B1(n_197),
.B2(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_11),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_175),
.B1(n_185),
.B2(n_179),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_177),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_201),
.C(n_45),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_175),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_21),
.C(n_38),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_35),
.B(n_49),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_205),
.B1(n_193),
.B2(n_191),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_33),
.B1(n_43),
.B2(n_39),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_187),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_202),
.B1(n_208),
.B2(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_12),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_212),
.C(n_34),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_37),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_14),
.B(n_15),
.Y(n_220)
);

XOR2x2_ASAP7_75t_R g221 ( 
.A(n_220),
.B(n_16),
.Y(n_221)
);


endmodule