module fake_jpeg_27043_n_166 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_5),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_14),
.B1(n_17),
.B2(n_11),
.Y(n_31)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_23),
.B1(n_25),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_12),
.B1(n_18),
.B2(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_22),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_14),
.B1(n_18),
.B2(n_21),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_28),
.B1(n_34),
.B2(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_30),
.B1(n_35),
.B2(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_33),
.Y(n_60)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_62),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_44),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_35),
.C(n_36),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_45),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_36),
.B1(n_28),
.B2(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_58),
.B1(n_74),
.B2(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_78),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_48),
.B1(n_39),
.B2(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_76),
.B1(n_57),
.B2(n_24),
.Y(n_82)
);

OAI22x1_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_42),
.B1(n_16),
.B2(n_13),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_43),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_56),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_81),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_53),
.B1(n_64),
.B2(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_53),
.B(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_66),
.C(n_68),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_98),
.C(n_81),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_66),
.C(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_67),
.C(n_72),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_116),
.B1(n_92),
.B2(n_24),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_79),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_107),
.C(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_115),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_72),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_83),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.C(n_114),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_84),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_24),
.C(n_29),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_21),
.A3(n_37),
.B1(n_12),
.B2(n_13),
.C1(n_16),
.C2(n_20),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_92),
.B1(n_97),
.B2(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_17),
.B1(n_27),
.B2(n_13),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_126),
.B1(n_27),
.B2(n_16),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.C(n_8),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_6),
.B(n_7),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_29),
.C(n_26),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_127),
.C(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_27),
.B1(n_13),
.B2(n_10),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_29),
.C(n_26),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_26),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_134),
.C(n_123),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_9),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_132),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_29),
.C(n_26),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_29),
.C(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_127),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_37),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_137),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_122),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_125),
.C(n_117),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_145),
.B(n_134),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_7),
.B(n_6),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_0),
.B(n_1),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_129),
.B(n_133),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_0),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_2),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_15),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_15),
.B(n_3),
.C(n_4),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_157),
.B1(n_148),
.B2(n_4),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_3),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_3),
.B1(n_4),
.B2(n_15),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_162),
.B(n_151),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_15),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_163),
.Y(n_166)
);


endmodule