module fake_jpeg_20422_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx13_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

AO22x1_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_6),
.B1(n_1),
.B2(n_5),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_5),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_13),
.B1(n_9),
.B2(n_7),
.Y(n_19)
);

AND2x4_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_32),
.B(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_24),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.C(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.C(n_33),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_35),
.B(n_29),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_40),
.Y(n_45)
);


endmodule