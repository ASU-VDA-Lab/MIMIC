module fake_jpeg_23578_n_163 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_36),
.Y(n_48)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_66),
.B1(n_34),
.B2(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_55),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.C(n_36),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_30),
.B1(n_22),
.B2(n_31),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_36),
.B(n_19),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_34),
.A2(n_30),
.B1(n_22),
.B2(n_31),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_86),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_27),
.Y(n_95)
);

AOI222xp33_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.C1(n_29),
.C2(n_27),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_93),
.B(n_67),
.C(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_18),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_60),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_91),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_33),
.B1(n_43),
.B2(n_35),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_21),
.B(n_25),
.C(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_107),
.B(n_69),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_1),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_113),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_33),
.B1(n_43),
.B2(n_19),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_102),
.B(n_111),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_1),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_114),
.B1(n_86),
.B2(n_75),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_4),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_4),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx10_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_102),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_129),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_76),
.B(n_71),
.C(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_126),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_125),
.B1(n_96),
.B2(n_130),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_85),
.B1(n_75),
.B2(n_89),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_90),
.B(n_9),
.C(n_8),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_88),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_81),
.B(n_90),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_122),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_138),
.B(n_134),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_142),
.B(n_137),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_145),
.C(n_144),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_145),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_156),
.A3(n_155),
.B1(n_150),
.B2(n_144),
.C1(n_118),
.C2(n_132),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_118),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_141),
.B(n_109),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_97),
.B(n_9),
.Y(n_161)
);

OAI21x1_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_8),
.B(n_11),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_13),
.Y(n_163)
);


endmodule