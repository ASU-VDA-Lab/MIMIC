module fake_jpeg_25266_n_235 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_19),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_30),
.B1(n_18),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_46),
.B1(n_53),
.B2(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_16),
.B1(n_19),
.B2(n_30),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_59),
.B1(n_15),
.B2(n_39),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_39),
.B1(n_35),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_54),
.B1(n_40),
.B2(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_33),
.B2(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_17),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_54),
.Y(n_107)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_72),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_84),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_36),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_79),
.C(n_54),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_75),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_25),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_83),
.B1(n_56),
.B2(n_47),
.Y(n_106)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_38),
.C(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_25),
.B1(n_20),
.B2(n_15),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_51),
.B1(n_61),
.B2(n_55),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_15),
.B1(n_20),
.B2(n_39),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_94),
.Y(n_121)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_69),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_102),
.B(n_106),
.Y(n_110)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_63),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_64),
.B1(n_65),
.B2(n_76),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_45),
.B(n_58),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_112),
.B1(n_127),
.B2(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_74),
.B1(n_81),
.B2(n_66),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_115),
.C(n_126),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_65),
.C(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_122),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_73),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_62),
.B(n_53),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_102),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_129),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_62),
.C(n_45),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_88),
.B(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_137),
.B(n_140),
.Y(n_158)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_85),
.B1(n_92),
.B2(n_89),
.C(n_106),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_145),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_87),
.B1(n_90),
.B2(n_105),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_90),
.B(n_99),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_99),
.B1(n_97),
.B2(n_89),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_112),
.B1(n_129),
.B2(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_99),
.B(n_91),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_143),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_39),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_132),
.C(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_86),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_109),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_78),
.B(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_148),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_119),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_94),
.B(n_101),
.Y(n_151)
);

BUFx12f_ASAP7_75t_SL g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_157),
.B1(n_169),
.B2(n_148),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_119),
.B1(n_108),
.B2(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_162),
.Y(n_171)
);

XOR2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_136),
.B1(n_143),
.B2(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_167),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_139),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_108),
.B1(n_61),
.B2(n_55),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_132),
.C(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_178),
.C(n_179),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_140),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_175),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_137),
.B(n_138),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_161),
.B(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_133),
.C(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_185),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_169),
.B1(n_152),
.B2(n_109),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_157),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_153),
.B1(n_161),
.B2(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_176),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_169),
.B1(n_167),
.B2(n_94),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_169),
.B1(n_101),
.B2(n_98),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_178),
.C(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_205),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_175),
.B(n_174),
.C(n_185),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_196),
.B1(n_198),
.B2(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_44),
.C(n_78),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_1),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_210),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_188),
.C(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_216),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_52),
.C(n_3),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_207),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_207),
.B1(n_204),
.B2(n_202),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_2),
.B(n_4),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_213),
.B(n_209),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_226),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_214),
.B(n_3),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_227),
.C(n_222),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_2),
.B(n_4),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_6),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_6),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_52),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_9),
.B(n_10),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_232),
.B1(n_12),
.B2(n_11),
.C(n_47),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_234),
.B(n_12),
.CI(n_208),
.CON(n_235),
.SN(n_235)
);


endmodule