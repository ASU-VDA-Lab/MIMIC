module fake_jpeg_26852_n_310 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_20),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_41),
.C(n_34),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_16),
.C(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_26),
.B1(n_17),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_30),
.B1(n_17),
.B2(n_21),
.Y(n_64)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

AO22x2_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_36),
.B1(n_30),
.B2(n_37),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_47),
.B1(n_32),
.B2(n_34),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_35),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_59),
.B(n_67),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_61),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_26),
.B1(n_15),
.B2(n_27),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_27),
.B1(n_15),
.B2(n_25),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_68),
.Y(n_93)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_30),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_70),
.Y(n_96)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_40),
.B(n_17),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_80),
.B(n_88),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_26),
.B1(n_51),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_75),
.B1(n_63),
.B2(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_40),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_69),
.B1(n_53),
.B2(n_97),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_47),
.B1(n_34),
.B2(n_32),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_94),
.B1(n_100),
.B2(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_42),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_34),
.B1(n_37),
.B2(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_65),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_55),
.C(n_56),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_104),
.B(n_107),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_106),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_55),
.B(n_72),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_99),
.B(n_96),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_114),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_120),
.B1(n_37),
.B2(n_28),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_98),
.B1(n_84),
.B2(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_113),
.B(n_125),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_87),
.B(n_92),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_79),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_56),
.C(n_37),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_90),
.C(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_117),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_73),
.B1(n_71),
.B2(n_54),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_102),
.B1(n_43),
.B2(n_105),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_87),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_122),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_126),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_31),
.B1(n_35),
.B2(n_33),
.Y(n_124)
);

AO21x2_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_42),
.B(n_85),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_31),
.B(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_140),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_141),
.B1(n_155),
.B2(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_139),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_149),
.C(n_33),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_24),
.B(n_1),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_84),
.B1(n_76),
.B2(n_57),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_142),
.B1(n_157),
.B2(n_29),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

XNOR2x1_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_113),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_76),
.B1(n_62),
.B2(n_54),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_148),
.B1(n_117),
.B2(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_109),
.B1(n_28),
.B2(n_65),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_96),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_151),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_85),
.C(n_33),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_19),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_14),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_28),
.B1(n_21),
.B2(n_70),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_106),
.B(n_27),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_161),
.A2(n_178),
.B(n_179),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_163),
.A2(n_168),
.B1(n_172),
.B2(n_183),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_181),
.C(n_184),
.Y(n_206)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_176),
.B1(n_187),
.B2(n_146),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_21),
.B1(n_28),
.B2(n_16),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_175),
.B1(n_149),
.B2(n_157),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_109),
.B1(n_22),
.B2(n_20),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_171),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_20),
.B1(n_18),
.B2(n_22),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_133),
.Y(n_199)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_31),
.B1(n_24),
.B2(n_20),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_185),
.B1(n_192),
.B2(n_4),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_132),
.B(n_131),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_29),
.C(n_22),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_19),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_24),
.B1(n_18),
.B2(n_14),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_188),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_0),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_154),
.B1(n_138),
.B2(n_155),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_137),
.B1(n_129),
.B2(n_148),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_166),
.B1(n_176),
.B2(n_174),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_202),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_200),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_150),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_127),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_211),
.B1(n_216),
.B2(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_0),
.CI(n_1),
.CON(n_205),
.SN(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_170),
.B(n_2),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_2),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_213),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_163),
.B1(n_168),
.B2(n_172),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_225),
.B1(n_226),
.B2(n_232),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_233),
.B1(n_6),
.B2(n_7),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_162),
.B1(n_191),
.B2(n_175),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_199),
.C(n_181),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_238),
.C(n_209),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_185),
.B1(n_177),
.B2(n_160),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_160),
.B1(n_183),
.B2(n_173),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_213),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_4),
.C(n_5),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_214),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_222),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_193),
.C(n_217),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_252),
.C(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_255),
.B1(n_232),
.B2(n_224),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_205),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_194),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_194),
.C(n_7),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_194),
.C(n_7),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_260),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_228),
.B1(n_233),
.B2(n_224),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_239),
.C(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_269),
.C(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_222),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_264),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_223),
.B1(n_221),
.B2(n_238),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_8),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_219),
.C(n_8),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_274),
.Y(n_284)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_280),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_6),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_279),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_6),
.C(n_8),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_260),
.B1(n_268),
.B2(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_9),
.C(n_10),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_9),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_9),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_9),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_261),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_287),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_286),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_263),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_262),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_276),
.B(n_277),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_298),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_279),
.C(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.C(n_299),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_10),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_10),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_10),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_302),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_294),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_297),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_304),
.C(n_11),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_11),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_12),
.B(n_297),
.Y(n_310)
);


endmodule