module fake_jpeg_13394_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_8),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_33),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_60),
.B(n_48),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_90),
.B(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_91),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_53),
.B1(n_68),
.B2(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_51),
.B1(n_61),
.B2(n_63),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_63),
.B1(n_71),
.B2(n_57),
.Y(n_111)
);

XOR2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_69),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_100),
.C(n_105),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_56),
.B(n_55),
.C(n_71),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2x1p5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_62),
.C(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_113),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_115),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_24),
.C(n_46),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_1),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_2),
.B(n_5),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_126),
.B(n_18),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_127),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_5),
.B(n_6),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_7),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_11),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_11),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_13),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_31),
.Y(n_148)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_16),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_140),
.C(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_19),
.C(n_20),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_22),
.C(n_25),
.Y(n_146)
);

NOR4xp25_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.D(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_117),
.C(n_129),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_117),
.B(n_136),
.C(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_34),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_156),
.C(n_145),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_137),
.B1(n_134),
.B2(n_39),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_143),
.B1(n_138),
.B2(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_162),
.B1(n_143),
.B2(n_138),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_141),
.B(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_157),
.C(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_144),
.C(n_159),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_134),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_37),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_38),
.Y(n_171)
);


endmodule