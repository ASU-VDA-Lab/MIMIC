module fake_jpeg_26763_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_17),
.Y(n_46)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_59),
.B1(n_65),
.B2(n_19),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_61),
.Y(n_66)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_63),
.Y(n_90)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_30),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_25),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_70),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_75),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_41),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_26),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

FAx1_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_38),
.CI(n_41),
.CON(n_76),
.SN(n_76)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_25),
.B(n_23),
.Y(n_117)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_42),
.B1(n_64),
.B2(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_92),
.B(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_46),
.B(n_26),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_22),
.C(n_31),
.Y(n_116)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_97),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_105),
.B(n_117),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_104),
.B1(n_108),
.B2(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_51),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_114),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_47),
.B1(n_40),
.B2(n_49),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_47),
.B1(n_40),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_113),
.B1(n_120),
.B2(n_84),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_91),
.B1(n_69),
.B2(n_71),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_82),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_75),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_29),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_118),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_42),
.B1(n_18),
.B2(n_31),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_71),
.B1(n_78),
.B2(n_88),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_125),
.B1(n_134),
.B2(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_90),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_78),
.B1(n_86),
.B2(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_136),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_78),
.B1(n_79),
.B2(n_85),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_105),
.C(n_116),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_89),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_60),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_60),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_143),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_84),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_73),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_163),
.C(n_173),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_108),
.B1(n_110),
.B2(n_101),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_159),
.B1(n_174),
.B2(n_125),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_167),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_119),
.B1(n_107),
.B2(n_115),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_176),
.B1(n_178),
.B2(n_131),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_107),
.C(n_114),
.Y(n_163)
);

OAI22x1_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_177),
.B1(n_21),
.B2(n_121),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

AND2x4_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_22),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_129),
.B(n_124),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_145),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_22),
.C(n_28),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_25),
.B1(n_27),
.B2(n_20),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_179),
.Y(n_190)
);

OAI22x1_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_21),
.B1(n_18),
.B2(n_4),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_194),
.B1(n_195),
.B2(n_207),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_127),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_168),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_130),
.C(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_192),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_127),
.B(n_136),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_193),
.B(n_196),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_128),
.C(n_122),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_203),
.C(n_204),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_140),
.B(n_139),
.C(n_126),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_172),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_123),
.C(n_141),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_141),
.C(n_21),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_141),
.B(n_2),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_1),
.Y(n_227)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_10),
.C(n_14),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_170),
.C(n_178),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_173),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_213),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_164),
.B1(n_153),
.B2(n_177),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_217),
.B1(n_220),
.B2(n_224),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_218),
.Y(n_254)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_219),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_164),
.B1(n_150),
.B2(n_167),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_155),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_157),
.CI(n_155),
.CON(n_219),
.SN(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_157),
.B1(n_161),
.B2(n_165),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_161),
.B1(n_10),
.B2(n_5),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_10),
.C(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_228),
.C(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_15),
.C(n_9),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_11),
.C(n_14),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_190),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_190),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_204),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_242),
.A2(n_244),
.B(n_1),
.Y(n_269)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_251),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_196),
.B(n_232),
.C(n_226),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_228),
.B(n_11),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_182),
.B1(n_195),
.B2(n_187),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_188),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_213),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_266),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_235),
.C(n_250),
.Y(n_271)
);

NAND2xp67_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_263),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_218),
.C(n_214),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_262),
.C(n_252),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_209),
.C(n_203),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_195),
.B(n_227),
.C(n_208),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_231),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_7),
.B(n_13),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_1),
.B(n_2),
.Y(n_272)
);

AOI31xp67_ASAP7_75t_SL g270 ( 
.A1(n_237),
.A2(n_236),
.A3(n_250),
.B(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_278),
.C(n_255),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_279),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_242),
.C(n_243),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_234),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_280),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_284),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_7),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_6),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_261),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_268),
.B1(n_263),
.B2(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_293),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_266),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_302),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_258),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_258),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_12),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_294),
.B(n_288),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_307),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_288),
.B(n_291),
.Y(n_309)
);

OAI21x1_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_301),
.B(n_311),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_302),
.B(n_12),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_310),
.C(n_306),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B1(n_313),
.B2(n_15),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_15),
.B(n_1),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_2),
.Y(n_321)
);


endmodule