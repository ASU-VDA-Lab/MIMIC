module fake_jpeg_5928_n_93 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_13),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_2),
.Y(n_59)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_3),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_55),
.B2(n_52),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_46),
.B1(n_51),
.B2(n_41),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_66),
.C(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_56),
.B1(n_49),
.B2(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_50),
.B1(n_40),
.B2(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_68),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_78),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_67),
.B1(n_47),
.B2(n_9),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_77),
.C(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_68),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_82),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_81),
.B1(n_80),
.B2(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_25),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_88),
.B(n_26),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_28),
.C(n_29),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_30),
.B(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_37),
.Y(n_93)
);


endmodule