module fake_jpeg_8307_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_7),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_27),
.B1(n_16),
.B2(n_17),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_39),
.A2(n_22),
.B1(n_25),
.B2(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_43),
.B1(n_52),
.B2(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_23),
.B1(n_27),
.B2(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_55),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_28),
.A2(n_27),
.B1(n_16),
.B2(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_22),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_59),
.B1(n_65),
.B2(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_69),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_28),
.B1(n_13),
.B2(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_33),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_15),
.B1(n_17),
.B2(n_13),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_13),
.B1(n_25),
.B2(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_75),
.B1(n_42),
.B2(n_43),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_87),
.B1(n_45),
.B2(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_49),
.B1(n_54),
.B2(n_38),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_95),
.B1(n_68),
.B2(n_44),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_60),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_52),
.B1(n_49),
.B2(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_100),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_56),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_18),
.C(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_110),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_115),
.B1(n_90),
.B2(n_19),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_60),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_20),
.B(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_57),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_114),
.B(n_89),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_26),
.B(n_19),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_116),
.B1(n_104),
.B2(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_44),
.B1(n_62),
.B2(n_67),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_45),
.B1(n_62),
.B2(n_34),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_96),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_127),
.C(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_115),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_96),
.A3(n_89),
.B1(n_29),
.B2(n_53),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_63),
.B(n_53),
.Y(n_123)
);

AOI22x1_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_26),
.B1(n_0),
.B2(n_3),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_80),
.B1(n_85),
.B2(n_20),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_128),
.B(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_138),
.B1(n_117),
.B2(n_90),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_92),
.B(n_64),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_132),
.B(n_128),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_112),
.B(n_99),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_80),
.B1(n_94),
.B2(n_63),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_139),
.B1(n_26),
.B2(n_1),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_97),
.Y(n_141)
);

AOI22x1_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_19),
.B1(n_26),
.B2(n_24),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_103),
.B1(n_114),
.B2(n_26),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_26),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_90),
.B1(n_26),
.B2(n_24),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_132),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_157),
.B(n_9),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_135),
.B1(n_129),
.B2(n_122),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_155),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_113),
.B(n_111),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_8),
.B(n_2),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_109),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_127),
.C(n_125),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

AOI22x1_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_136),
.B1(n_139),
.B2(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_7),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_7),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_124),
.B1(n_119),
.B2(n_3),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_181),
.B(n_158),
.Y(n_191)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_130),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_170),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_147),
.B1(n_156),
.B2(n_152),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_129),
.C(n_138),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_177),
.B(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_8),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_9),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_2),
.Y(n_184)
);

OA21x2_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_4),
.B(n_5),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_149),
.B(n_155),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_190),
.B1(n_169),
.B2(n_166),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_203),
.B1(n_177),
.B2(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_194),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_147),
.B(n_146),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_162),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_154),
.B(n_2),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_182),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_184),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_4),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_10),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_220),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_167),
.B1(n_163),
.B2(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_179),
.C(n_171),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_216),
.C(n_219),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_209),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_180),
.B1(n_165),
.B2(n_170),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_199),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_202),
.B1(n_187),
.B2(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_180),
.C(n_183),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_165),
.B1(n_174),
.B2(n_5),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_0),
.C(n_4),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_234),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_216),
.C(n_219),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_234),
.C(n_212),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_232),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_190),
.B1(n_194),
.B2(n_189),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_231),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_192),
.C(n_202),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_217),
.B(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_242),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_185),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_201),
.C(n_191),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_198),
.C(n_0),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_245),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_12),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_10),
.B(n_11),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_231),
.B(n_233),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_225),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_249),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_222),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_240),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_262),
.B1(n_253),
.B2(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_10),
.C(n_11),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_266),
.B(n_257),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

A2O1A1O1Ixp25_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_251),
.B(n_260),
.C(n_12),
.D(n_10),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_264),
.B(n_265),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_268),
.C(n_11),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_11),
.C(n_12),
.Y(n_273)
);


endmodule