module real_jpeg_4209_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g126 ( 
.A(n_0),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_1),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_2),
.A2(n_84),
.B1(n_137),
.B2(n_213),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_2),
.A2(n_84),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_2),
.A2(n_84),
.B1(n_248),
.B2(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_3),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_4),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_4),
.A2(n_74),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_5),
.A2(n_85),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_5),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_99),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_5),
.A2(n_99),
.B1(n_154),
.B2(n_203),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_5),
.A2(n_99),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_6),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_7),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g356 ( 
.A(n_7),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_8),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_8),
.A2(n_136),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_8),
.A2(n_136),
.B1(n_193),
.B2(n_295),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_8),
.A2(n_136),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_9),
.A2(n_42),
.B1(n_176),
.B2(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_165),
.C(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_9),
.B(n_122),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_9),
.B(n_65),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_9),
.B(n_181),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_9),
.B(n_213),
.Y(n_352)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_12),
.Y(n_208)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_12),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_13),
.A2(n_56),
.B1(n_61),
.B2(n_64),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_13),
.A2(n_64),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_14),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_14),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_14),
.A2(n_118),
.B1(n_179),
.B2(n_224),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_14),
.A2(n_76),
.B1(n_179),
.B2(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_15),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_15),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_16),
.A2(n_168),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_254),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_253),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_214),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_21),
.B(n_214),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_148),
.C(n_199),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_22),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_78),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_23),
.B(n_79),
.C(n_110),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_24),
.A2(n_46),
.B1(n_47),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.A3(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_28),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_29),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_29),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_29),
.Y(n_146)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_34),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_88)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_35),
.A2(n_102),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_41),
.A2(n_42),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_42),
.B(n_88),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_42),
.A2(n_48),
.B(n_297),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_42),
.A2(n_350),
.B(n_351),
.Y(n_349)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_54),
.B1(n_65),
.B2(n_68),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_48),
.A2(n_191),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_48),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_49),
.A2(n_69),
.B1(n_190),
.B2(n_195),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_49),
.A2(n_55),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_49),
.B(n_298),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_49),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_51),
.Y(n_269)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_53),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_59),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_63),
.Y(n_296)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_70),
.Y(n_291)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_77),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_109),
.B2(n_110),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_86),
.B(n_97),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_81),
.A2(n_88),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_87),
.B(n_98),
.Y(n_210)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_94),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_103),
.A2(n_206),
.B(n_209),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_103),
.Y(n_226)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_130),
.B(n_141),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g220 ( 
.A1(n_111),
.A2(n_122),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_111),
.B(n_221),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_111),
.A2(n_141),
.B(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_112),
.A2(n_131),
.B1(n_147),
.B2(n_212),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_113)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_114),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_117),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

AO22x2_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_122)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_125),
.Y(n_239)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_126),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_126),
.Y(n_308)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_135),
.Y(n_359)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_147),
.A2(n_212),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_148),
.A2(n_149),
.B1(n_199),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_189),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_150),
.B(n_189),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_175),
.B1(n_180),
.B2(n_182),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_151),
.A2(n_283),
.B(n_286),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_151),
.A2(n_180),
.B1(n_305),
.B2(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_151),
.A2(n_286),
.B(n_343),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_152),
.A2(n_181),
.B1(n_183),
.B2(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_164),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_159),
.B2(n_161),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_161),
.Y(n_289)
);

INVx5_ASAP7_75t_SL g346 ( 
.A(n_161),
.Y(n_346)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_175),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_164),
.A2(n_201),
.B(n_305),
.Y(n_304)
);

AOI22x1_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_170),
.B2(n_172),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_169),
.Y(n_301)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_178),
.Y(n_306)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_181),
.B(n_202),
.Y(n_286)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g360 ( 
.A(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.C(n_211),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_200),
.B(n_211),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_204),
.A2(n_205),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_233),
.B1(n_251),
.B2(n_252),
.Y(n_216)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_225),
.B1(n_231),
.B2(n_232),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_236),
.Y(n_344)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_241),
.Y(n_332)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_276),
.B(n_385),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_273),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_257),
.B(n_273),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.C(n_264),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_258),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_264),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.C(n_272),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_265),
.B(n_376),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_267),
.B(n_272),
.Y(n_376)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_379),
.B(n_384),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_368),
.B(n_378),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_337),
.B(n_367),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_311),
.B(n_336),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_292),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_292),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_282),
.A2(n_287),
.B1(n_288),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_284),
.B(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_303),
.C(n_310),
.Y(n_338)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_309),
.B2(n_310),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_328),
.B(n_335),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_318),
.B(n_327),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_326),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_323),
.B(n_325),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_333),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_339),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_353),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_347),
.B2(n_348),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_347),
.C(n_353),
.Y(n_369)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI32xp33_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_358),
.A3(n_360),
.B1(n_361),
.B2(n_365),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_357),
.Y(n_374)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_369),
.B(n_370),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_375),
.B2(n_377),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_374),
.C(n_377),
.Y(n_380)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);


endmodule