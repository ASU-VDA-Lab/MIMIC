module fake_jpeg_16973_n_394 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_394);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_394;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_48),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_34),
.B1(n_23),
.B2(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_69),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_77),
.A2(n_7),
.B(n_11),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_36),
.B1(n_31),
.B2(n_14),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_30),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_84),
.A2(n_118),
.B1(n_111),
.B2(n_105),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_88),
.B(n_94),
.Y(n_171)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_32),
.B1(n_28),
.B2(n_33),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_103),
.B1(n_40),
.B2(n_7),
.Y(n_166)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_38),
.B1(n_37),
.B2(n_29),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_49),
.B(n_18),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_39),
.B(n_26),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_120),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_67),
.A2(n_26),
.B1(n_17),
.B2(n_22),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_39),
.B(n_22),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_121),
.B(n_127),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_78),
.B(n_66),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_132),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_136),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_17),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_17),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_147),
.Y(n_192)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_114),
.B1(n_59),
.B2(n_105),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_165),
.B1(n_170),
.B2(n_72),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_70),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_46),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_159),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_17),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_22),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_157),
.Y(n_202)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_81),
.A2(n_22),
.B1(n_60),
.B2(n_58),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_154),
.A2(n_169),
.B(n_4),
.Y(n_210)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_98),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_46),
.C(n_44),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_106),
.C(n_5),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_44),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_98),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_167),
.Y(n_208)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_71),
.B(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_109),
.Y(n_189)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_107),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_104),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_72),
.B1(n_119),
.B2(n_81),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_175),
.A2(n_147),
.B1(n_130),
.B2(n_126),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_157),
.B1(n_161),
.B2(n_154),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_178),
.A2(n_213),
.B1(n_143),
.B2(n_167),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_13),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_183),
.A2(n_195),
.B(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_122),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_191),
.Y(n_237)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_107),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_216),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_207),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_138),
.A2(n_117),
.B(n_100),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_70),
.B1(n_91),
.B2(n_75),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_196),
.A2(n_199),
.B1(n_203),
.B2(n_215),
.Y(n_257)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_74),
.B1(n_75),
.B2(n_9),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_146),
.B(n_74),
.CI(n_113),
.CON(n_200),
.SN(n_200)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_127),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_0),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_135),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_210),
.A2(n_155),
.B1(n_134),
.B2(n_3),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_4),
.Y(n_211)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_143),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_4),
.B(n_10),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_183),
.B(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_11),
.C(n_3),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_171),
.C(n_129),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_0),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_165),
.A2(n_3),
.B(n_5),
.C(n_8),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_219),
.A2(n_258),
.B(n_191),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_221),
.B(n_229),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_131),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_137),
.B1(n_141),
.B2(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_230),
.B1(n_232),
.B2(n_238),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_247),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_121),
.C(n_145),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_242),
.C(n_246),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_123),
.C(n_155),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_228),
.B(n_233),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_126),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_176),
.A2(n_168),
.B1(n_145),
.B2(n_124),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_3),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_125),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_249),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_124),
.B1(n_160),
.B2(n_149),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_241),
.A2(n_252),
.B1(n_259),
.B2(n_240),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_133),
.C(n_125),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_144),
.B1(n_133),
.B2(n_8),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_253),
.B(n_206),
.Y(n_278)
);

OAI211xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_8),
.B(n_11),
.C(n_2),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_8),
.C(n_1),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_1),
.B1(n_2),
.B2(n_200),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_248),
.A2(n_212),
.B1(n_188),
.B2(n_209),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_180),
.B(n_1),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_202),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_201),
.B(n_190),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_179),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_206),
.B1(n_182),
.B2(n_185),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_211),
.A2(n_196),
.B(n_214),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_211),
.A2(n_175),
.B1(n_179),
.B2(n_174),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_272),
.B(n_283),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_242),
.C(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_270),
.C(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_184),
.C(n_174),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_227),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_172),
.B(n_177),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g273 ( 
.A1(n_221),
.A2(n_219),
.B1(n_259),
.B2(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_235),
.A2(n_213),
.B1(n_177),
.B2(n_172),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_278),
.B(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_284),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_248),
.B1(n_243),
.B2(n_238),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_231),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_185),
.B1(n_212),
.B2(n_209),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_286),
.A2(n_293),
.B1(n_280),
.B2(n_281),
.Y(n_318)
);

XOR2x1_ASAP7_75t_SL g288 ( 
.A(n_221),
.B(n_205),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_251),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_232),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_235),
.A2(n_188),
.B1(n_186),
.B2(n_197),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_204),
.B1(n_205),
.B2(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_294),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_296),
.A2(n_317),
.B1(n_320),
.B2(n_302),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_258),
.B(n_234),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_276),
.B1(n_264),
.B2(n_262),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_265),
.A2(n_226),
.B1(n_220),
.B2(n_241),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_302),
.B1(n_311),
.B2(n_313),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_234),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_226),
.C(n_247),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_287),
.B(n_223),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_310),
.B(n_321),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_246),
.B1(n_255),
.B2(n_233),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_252),
.B1(n_244),
.B2(n_249),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_263),
.B(n_239),
.C(n_204),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_316),
.C(n_293),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_244),
.C(n_283),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_273),
.A2(n_268),
.B1(n_286),
.B2(n_275),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_280),
.B1(n_290),
.B2(n_277),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_268),
.A2(n_273),
.B1(n_292),
.B2(n_274),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_276),
.C(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_295),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_323),
.A2(n_329),
.B1(n_342),
.B2(n_336),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_324),
.A2(n_336),
.B(n_344),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_333),
.C(n_334),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_314),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_343),
.B(n_300),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_285),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_264),
.C(n_291),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_313),
.B(n_277),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_320),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_304),
.B(n_317),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_318),
.B1(n_303),
.B2(n_316),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_338),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_307),
.C(n_315),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_311),
.C(n_309),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_312),
.B1(n_303),
.B2(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_341),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_312),
.A2(n_298),
.B1(n_299),
.B2(n_314),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_319),
.Y(n_343)
);

XOR2x2_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_297),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_300),
.C(n_299),
.Y(n_345)
);

NOR4xp25_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_340),
.C(n_342),
.D(n_356),
.Y(n_364)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_355),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_326),
.C(n_331),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_350),
.B(n_353),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_351),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_343),
.B(n_304),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_325),
.Y(n_354)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_334),
.C(n_328),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_333),
.C(n_338),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_361),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_360),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_344),
.C(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_337),
.Y(n_362)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_349),
.B1(n_359),
.B2(n_348),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_327),
.Y(n_365)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

AOI322xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_324),
.A3(n_330),
.B1(n_335),
.B2(n_341),
.C1(n_357),
.C2(n_358),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_371),
.B(n_373),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_361),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_369),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_372),
.A2(n_350),
.B1(n_348),
.B2(n_355),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_375),
.B(n_379),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g379 ( 
.A(n_365),
.B(n_362),
.CI(n_363),
.CON(n_379),
.SN(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_377),
.B(n_367),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_380),
.A2(n_370),
.B1(n_368),
.B2(n_378),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_379),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_367),
.B(n_373),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_383),
.A2(n_376),
.B(n_368),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_379),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_386),
.Y(n_388)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_387),
.A2(n_378),
.B(n_382),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_387),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_388),
.C(n_375),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_372),
.B(n_366),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_366),
.C(n_369),
.Y(n_394)
);


endmodule