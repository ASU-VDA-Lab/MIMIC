module fake_jpeg_14140_n_507 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_507);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_507;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_65),
.Y(n_123)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_63),
.B(n_69),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_18),
.B(n_11),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_72),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_67),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_68),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_18),
.B(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_71),
.B(n_80),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_22),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_73),
.Y(n_186)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_83),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_78),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_79),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_82),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_91),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_90),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_16),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_94),
.B(n_117),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_97),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_44),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_105),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_40),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_113),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_28),
.B(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_28),
.B(n_14),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_119),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_40),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_120),
.A2(n_117),
.B(n_93),
.Y(n_196)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_6),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_62),
.A2(n_50),
.B1(n_53),
.B2(n_43),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_128),
.A2(n_146),
.B1(n_150),
.B2(n_169),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_56),
.B1(n_55),
.B2(n_48),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_130),
.A2(n_133),
.B1(n_137),
.B2(n_142),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_105),
.B1(n_89),
.B2(n_75),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_27),
.B1(n_43),
.B2(n_42),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_64),
.A2(n_56),
.B1(n_55),
.B2(n_48),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_188),
.C(n_195),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_89),
.A2(n_20),
.B1(n_41),
.B2(n_37),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_79),
.B1(n_76),
.B2(n_67),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_74),
.A2(n_20),
.B(n_41),
.C(n_37),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_149),
.A2(n_153),
.B(n_161),
.C(n_198),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_38),
.B1(n_36),
.B2(n_31),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_78),
.A2(n_19),
.B1(n_33),
.B2(n_27),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_167),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_78),
.A2(n_33),
.B1(n_24),
.B2(n_19),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_60),
.A2(n_38),
.B1(n_36),
.B2(n_31),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_84),
.A2(n_109),
.B1(n_115),
.B2(n_101),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_82),
.A2(n_42),
.B1(n_24),
.B2(n_14),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_103),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_170),
.A2(n_171),
.B1(n_178),
.B2(n_195),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_113),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_57),
.A2(n_13),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_172),
.A2(n_192),
.B(n_196),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_118),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_85),
.A2(n_6),
.B1(n_97),
.B2(n_92),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_197),
.B1(n_199),
.B2(n_163),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_86),
.A2(n_119),
.B1(n_107),
.B2(n_100),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_140),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_100),
.A2(n_68),
.B1(n_93),
.B2(n_59),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_98),
.B(n_68),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_194),
.B(n_136),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_117),
.A2(n_88),
.B1(n_46),
.B2(n_40),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_98),
.A2(n_111),
.B1(n_112),
.B2(n_69),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_88),
.A2(n_46),
.B1(n_40),
.B2(n_105),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_163),
.B1(n_193),
.B2(n_147),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_61),
.A2(n_47),
.B1(n_67),
.B2(n_76),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_201),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_202),
.B(n_214),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_204),
.Y(n_302)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_206),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_208),
.Y(n_289)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_215),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_211),
.A2(n_178),
.B1(n_181),
.B2(n_238),
.Y(n_285)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g277 ( 
.A(n_212),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_135),
.B(n_123),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_213),
.B(n_221),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_143),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_140),
.A2(n_185),
.B1(n_164),
.B2(n_168),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_217),
.A2(n_232),
.B1(n_237),
.B2(n_230),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_218),
.Y(n_282)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_160),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_175),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_134),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_231),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_184),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_SL g313 ( 
.A(n_225),
.B(n_239),
.C(n_265),
.Y(n_313)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_139),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_155),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_262),
.C(n_256),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_200),
.B1(n_159),
.B2(n_188),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_144),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_122),
.Y(n_234)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_145),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_235),
.B(n_238),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_137),
.B(n_142),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_125),
.Y(n_241)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_154),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_173),
.B(n_126),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_243),
.B(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_126),
.B(n_190),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_258),
.B(n_267),
.Y(n_280)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_183),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_190),
.B(n_162),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_259),
.Y(n_294)
);

BUFx6f_ASAP7_75t_SL g251 ( 
.A(n_158),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_124),
.Y(n_252)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_167),
.Y(n_253)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_147),
.Y(n_254)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_158),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_124),
.Y(n_257)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_127),
.B(n_138),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_138),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_261),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_193),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_170),
.B(n_171),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_229),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_191),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_254),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_191),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_207),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_272),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_285),
.A2(n_305),
.B(n_306),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_202),
.B1(n_253),
.B2(n_211),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_286),
.A2(n_244),
.B1(n_234),
.B2(n_219),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_287),
.B(n_318),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_214),
.C(n_203),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_220),
.C(n_241),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_295),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_202),
.A2(n_242),
.B(n_256),
.Y(n_305)
);

INVx13_ASAP7_75t_L g307 ( 
.A(n_216),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_208),
.B(n_210),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_311),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_239),
.A2(n_246),
.B(n_262),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_314),
.A2(n_317),
.B(n_316),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_316),
.A2(n_247),
.B(n_251),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_240),
.A2(n_224),
.B(n_248),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_207),
.A2(n_237),
.B1(n_249),
.B2(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_225),
.B(n_236),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_320),
.A2(n_332),
.B(n_335),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_352),
.B1(n_356),
.B2(n_303),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_270),
.B(n_205),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_323),
.B(n_324),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_270),
.B(n_222),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_320),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_275),
.B(n_310),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_327),
.B(n_334),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_268),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_331),
.Y(n_359)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_287),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_209),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_336),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_271),
.B(n_206),
.Y(n_334)
);

A2O1A1O1Ixp25_ASAP7_75t_L g335 ( 
.A1(n_306),
.A2(n_257),
.B(n_259),
.C(n_260),
.D(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_294),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_355),
.Y(n_366)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_212),
.B1(n_226),
.B2(n_228),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_338),
.B(n_342),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_278),
.A2(n_298),
.B(n_285),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_278),
.B(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_345),
.Y(n_361)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_281),
.B(n_312),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_344),
.B(n_353),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_294),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_348),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_308),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_296),
.B(n_280),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_309),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_350),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_309),
.B(n_274),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_354),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_274),
.A2(n_296),
.B1(n_311),
.B2(n_289),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_282),
.B(n_302),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_274),
.A2(n_309),
.B(n_282),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_276),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_299),
.A2(n_277),
.B1(n_303),
.B2(n_284),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_293),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_380),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_292),
.C(n_308),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_346),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_370),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_371),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_343),
.A2(n_277),
.B1(n_291),
.B2(n_301),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_368),
.A2(n_374),
.B1(n_381),
.B2(n_358),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_353),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_343),
.A2(n_291),
.B1(n_301),
.B2(n_283),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_373),
.A2(n_378),
.B1(n_322),
.B2(n_352),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_315),
.B1(n_283),
.B2(n_290),
.Y(n_374)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_377),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_321),
.A2(n_340),
.B1(n_345),
.B2(n_332),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_290),
.A3(n_293),
.B1(n_273),
.B2(n_304),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_315),
.B1(n_304),
.B2(n_273),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_328),
.B(n_300),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_355),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_276),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_320),
.Y(n_396)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_362),
.Y(n_393)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_365),
.A2(n_332),
.B1(n_339),
.B2(n_350),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_394),
.A2(n_408),
.B1(n_412),
.B2(n_378),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_396),
.B(n_371),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_366),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_405),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g398 ( 
.A(n_363),
.B(n_324),
.C(n_347),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_398),
.B(n_404),
.Y(n_423)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_399),
.Y(n_416)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

INVx8_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_337),
.Y(n_402)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_402),
.Y(n_426)
);

OAI21xp33_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_349),
.B(n_329),
.Y(n_403)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_369),
.C(n_388),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_379),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_385),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_330),
.Y(n_406)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_372),
.A2(n_348),
.B1(n_326),
.B2(n_327),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_381),
.B1(n_376),
.B2(n_382),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_385),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_413),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_372),
.A2(n_323),
.B1(n_354),
.B2(n_329),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_364),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_325),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_325),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_417),
.A2(n_429),
.B(n_434),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_389),
.A2(n_382),
.B1(n_375),
.B2(n_373),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_422),
.A2(n_410),
.B1(n_404),
.B2(n_395),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_364),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_425),
.A2(n_395),
.B(n_361),
.Y(n_449)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_428),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_389),
.A2(n_376),
.B(n_375),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_367),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_431),
.C(n_433),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_360),
.C(n_387),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_435),
.B(n_414),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_361),
.C(n_388),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_407),
.C(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_397),
.Y(n_440)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_440),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_442),
.A2(n_426),
.B1(n_427),
.B2(n_424),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_405),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_443),
.B(n_439),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_444),
.B(n_450),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_445),
.A2(n_446),
.B1(n_415),
.B2(n_421),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

INVx13_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_448),
.A2(n_453),
.B(n_423),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_449),
.A2(n_425),
.B(n_434),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_408),
.C(n_396),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_413),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_454),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_419),
.A2(n_411),
.B1(n_401),
.B2(n_406),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_455),
.B1(n_424),
.B2(n_420),
.Y(n_465)
);

A2O1A1O1Ixp25_ASAP7_75t_L g453 ( 
.A1(n_420),
.A2(n_398),
.B(n_412),
.C(n_391),
.D(n_335),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_391),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_401),
.B1(n_399),
.B2(n_390),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_457),
.A2(n_459),
.B(n_460),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_461),
.A2(n_463),
.B1(n_442),
.B2(n_452),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_438),
.A2(n_417),
.B1(n_422),
.B2(n_429),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_438),
.A2(n_426),
.B1(n_427),
.B2(n_436),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_447),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_468),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_455),
.A2(n_399),
.B1(n_392),
.B2(n_393),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_450),
.C(n_441),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_471),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_440),
.B(n_453),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_478),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_458),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_444),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_476),
.C(n_441),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_474),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_457),
.B(n_334),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_447),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_488),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_477),
.A2(n_456),
.B(n_443),
.Y(n_482)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_482),
.Y(n_494)
);

MAJx2_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_463),
.C(n_430),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_475),
.B(n_451),
.CI(n_449),
.CON(n_485),
.SN(n_485)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_486),
.Y(n_490)
);

FAx1_ASAP7_75t_SL g486 ( 
.A(n_475),
.B(n_467),
.CI(n_453),
.CON(n_486),
.SN(n_486)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_477),
.A2(n_467),
.B(n_460),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_487),
.A2(n_445),
.B1(n_446),
.B2(n_472),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_493),
.Y(n_496)
);

MAJx2_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_480),
.C(n_486),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_445),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_481),
.A2(n_446),
.B(n_465),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_495),
.A2(n_490),
.B1(n_494),
.B2(n_481),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_498),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_490),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_499),
.A2(n_500),
.B(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_485),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_502),
.B(n_448),
.C(n_431),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_448),
.A3(n_384),
.B1(n_344),
.B2(n_338),
.C1(n_380),
.C2(n_335),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_503),
.B(n_338),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_505),
.C(n_501),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_338),
.Y(n_507)
);


endmodule