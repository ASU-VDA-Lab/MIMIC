module real_jpeg_14926_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_411, n_6, n_7, n_3, n_10, n_412, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_411;
input n_6;
input n_7;
input n_3;
input n_10;
input n_412;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_108),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_113),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_3),
.B(n_26),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_3),
.B(n_29),
.Y(n_326)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_50),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_5),
.B(n_26),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_5),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_38),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_6),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_38),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_6),
.B(n_108),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_6),
.B(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_6),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_8),
.B(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_8),
.B(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_8),
.B(n_29),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_8),
.B(n_38),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_8),
.B(n_43),
.Y(n_289)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_50),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_38),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_108),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_10),
.B(n_113),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_10),
.B(n_26),
.Y(n_247)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_11),
.B(n_32),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_11),
.B(n_29),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_11),
.B(n_50),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_11),
.B(n_38),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_13),
.B(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_29),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_13),
.B(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_13),
.B(n_32),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_13),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_50),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_38),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_13),
.B(n_43),
.Y(n_259)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_14),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_14),
.B(n_113),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_14),
.B(n_32),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_14),
.B(n_26),
.Y(n_308)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_15),
.Y(n_104)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_77),
.B(n_343),
.C(n_407),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_87),
.B(n_406),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_21),
.B(n_75),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_61),
.C(n_62),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_22),
.B(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_45),
.C(n_52),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_23),
.B(n_394),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_35),
.C(n_39),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_25),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_54),
.C(n_59),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_25),
.A2(n_60),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_25),
.B(n_232),
.C(n_233),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_25),
.A2(n_31),
.B1(n_60),
.B2(n_181),
.Y(n_384)
);

INVx5_ASAP7_75t_SL g122 ( 
.A(n_26),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_28),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_28),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_28),
.B(n_272),
.C(n_275),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_28),
.A2(n_276),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_30),
.B(n_36),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_31),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_31),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_31),
.B(n_177),
.C(n_179),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_31),
.A2(n_134),
.B1(n_135),
.B2(n_181),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_31),
.B(n_134),
.C(n_247),
.Y(n_387)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_32),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_36),
.B(n_107),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_41),
.B(n_156),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_41),
.B(n_226),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_42),
.B(n_155),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_42),
.B(n_109),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_42),
.B(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_45),
.A2(n_52),
.B1(n_53),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_45),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.C(n_49),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_46),
.B(n_49),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_47),
.A2(n_85),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

NOR3xp33_ASAP7_75t_L g407 ( 
.A(n_47),
.B(n_66),
.C(n_83),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_48),
.B(n_156),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_50),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_54),
.A2(n_55),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_55),
.B(n_115),
.C(n_232),
.Y(n_339)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_64),
.C(n_66),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_58),
.A2(n_59),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_59),
.B(n_245),
.C(n_247),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_61),
.B(n_62),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_70),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_72),
.C(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_64),
.A2(n_68),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_64),
.B(n_352),
.C(n_353),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_67),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_66),
.A2(n_67),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_67),
.B(n_286),
.C(n_288),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_86),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_83),
.A2(n_84),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_84),
.B(n_308),
.C(n_311),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_401),
.B(n_405),
.Y(n_87)
);

OAI321xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_369),
.A3(n_389),
.B1(n_399),
.B2(n_400),
.C(n_411),
.Y(n_88)
);

AOI321xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_297),
.A3(n_329),
.B1(n_363),
.B2(n_368),
.C(n_412),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_236),
.C(n_292),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_204),
.B(n_235),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_171),
.B(n_203),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_139),
.B(n_170),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_116),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_95),
.B(n_116),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_110),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_119),
.B1(n_120),
.B2(n_128),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_167),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.CI(n_99),
.CON(n_96),
.SN(n_96)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_100),
.A2(n_101),
.B1(n_110),
.B2(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_106),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_103),
.B(n_155),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_105),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_114),
.A2(n_115),
.B1(n_185),
.B2(n_186),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_114),
.A2(n_115),
.B1(n_231),
.B2(n_232),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_115),
.B(n_186),
.C(n_289),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_129),
.B2(n_138),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_128),
.C(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_124),
.C(n_127),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_132),
.C(n_133),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_134),
.A2(n_135),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_134),
.A2(n_135),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_134),
.B(n_343),
.C(n_345),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_136),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_135),
.B(n_324),
.C(n_326),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_136),
.A2(n_137),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_136),
.B(n_259),
.C(n_262),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_164),
.B(n_169),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_152),
.B(n_163),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_150),
.C(n_151),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_158),
.B(n_162),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_173),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_189),
.B2(n_190),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_191),
.C(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_183),
.C(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_187),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_201),
.B2(n_202),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_200),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_197),
.C(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_206),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_222),
.B2(n_234),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_221),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_209),
.B(n_221),
.C(n_234),
.Y(n_293)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_218),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_219),
.C(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_213),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.CI(n_216),
.CON(n_213),
.SN(n_213)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_222),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.CI(n_229),
.CON(n_222),
.SN(n_222)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_224),
.C(n_229),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_227),
.B(n_228),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_227),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_228),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g364 ( 
.A1(n_237),
.A2(n_365),
.B(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_268),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_238),
.B(n_268),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_256),
.C(n_267),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_239),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_255),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_248),
.C(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_246),
.A2(n_247),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_252),
.C(n_254),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_256),
.A2(n_257),
.B1(n_267),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_264),
.C(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_291),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_280),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_280),
.C(n_291),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_278),
.C(n_279),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_294),
.Y(n_365)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_298),
.A2(n_364),
.B(n_367),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_299),
.B(n_300),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_328),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_303),
.C(n_328),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_320),
.B2(n_321),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_304),
.B(n_322),
.C(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_314),
.C(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_331),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_362),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_347),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_347),
.C(n_362),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_338),
.C(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_345),
.Y(n_338)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_354),
.B2(n_355),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_356),
.C(n_361),
.Y(n_372)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_360),
.B2(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_361),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_370),
.B(n_371),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_390),
.Y(n_400)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.CI(n_388),
.CON(n_371),
.SN(n_371)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_381),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_378),
.C(n_381),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_379),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_386),
.C(n_387),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_398),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_396),
.B2(n_397),
.Y(n_391)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_392),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_397),
.C(n_398),
.Y(n_402)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_403),
.Y(n_405)
);


endmodule