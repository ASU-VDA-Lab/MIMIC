module fake_jpeg_30553_n_262 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_59),
.Y(n_80)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_66),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_19),
.B(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_75),
.B1(n_85),
.B2(n_87),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_29),
.B1(n_31),
.B2(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_1),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_41),
.B1(n_25),
.B2(n_38),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_29),
.B1(n_41),
.B2(n_38),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_93),
.B1(n_53),
.B2(n_55),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_106)
);

AOI22x1_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_2),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_37),
.B1(n_28),
.B2(n_39),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_45),
.A2(n_28),
.B1(n_39),
.B2(n_3),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_117),
.B1(n_106),
.B2(n_118),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_81),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_114),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_109),
.Y(n_134)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_54),
.B1(n_46),
.B2(n_44),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_107),
.A2(n_108),
.B1(n_71),
.B2(n_76),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_43),
.B1(n_57),
.B2(n_50),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_49),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_49),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_49),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_122),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_39),
.B1(n_3),
.B2(n_5),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_111),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_51),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_2),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_2),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_3),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_151),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_93),
.B1(n_91),
.B2(n_84),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_145),
.B1(n_152),
.B2(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_93),
.B1(n_91),
.B2(n_82),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_74),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_99),
.B1(n_70),
.B2(n_88),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_99),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_74),
.B1(n_70),
.B2(n_71),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_77),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_103),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_132),
.B(n_138),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_167),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_136),
.C(n_133),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_169),
.C(n_124),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_130),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_181),
.B(n_137),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_128),
.C(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_129),
.A3(n_115),
.B1(n_123),
.B2(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_172),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_5),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_5),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_6),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_116),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_157),
.B(n_141),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_146),
.B(n_7),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_187),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_146),
.B(n_145),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_161),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_149),
.B1(n_152),
.B2(n_154),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_194),
.B1(n_162),
.B2(n_163),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_135),
.B1(n_143),
.B2(n_137),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_185),
.B1(n_182),
.B2(n_194),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_156),
.B(n_139),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_193),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_156),
.B(n_139),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_148),
.B1(n_143),
.B2(n_137),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_166),
.C(n_169),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_208),
.C(n_215),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_216),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_158),
.C(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_211),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_180),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_210),
.B(n_213),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_160),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_217),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_174),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_215),
.C(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_191),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_227),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_199),
.B1(n_184),
.B2(n_196),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_203),
.B(n_204),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_218),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_218),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_189),
.B(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_206),
.C(n_203),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_237),
.C(n_223),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_192),
.B1(n_199),
.B2(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_184),
.B1(n_219),
.B2(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_206),
.C(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_239),
.B(n_240),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_159),
.B(n_187),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_243),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_236),
.B(n_228),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_245),
.B(n_231),
.CI(n_237),
.CON(n_247),
.SN(n_247)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_230),
.B(n_238),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_245),
.C(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_249),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_225),
.B(n_191),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_188),
.C(n_193),
.Y(n_258)
);

NAND4xp25_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_229),
.C(n_234),
.D(n_225),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_253),
.A2(n_250),
.B(n_165),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_257),
.A3(n_258),
.B1(n_254),
.B2(n_171),
.C1(n_181),
.C2(n_179),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_239),
.Y(n_257)
);

OAI311xp33_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_260),
.A3(n_7),
.B1(n_10),
.C1(n_12),
.Y(n_261)
);

AOI211xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_167),
.B(n_8),
.C(n_9),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_10),
.Y(n_262)
);


endmodule