module fake_jpeg_26165_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_11),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_23),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_18),
.B1(n_9),
.B2(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_13),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_9),
.B1(n_19),
.B2(n_14),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_42),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_20),
.B1(n_22),
.B2(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_44),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_24),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_43),
.B(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_10),
.B(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_29),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_26),
.CON(n_47),
.SN(n_47)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_50),
.B(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_27),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_46),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_40),
.B1(n_41),
.B2(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_59),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_40),
.Y(n_59)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_28),
.B1(n_33),
.B2(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_33),
.B1(n_25),
.B2(n_28),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_53),
.C(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_15),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_76),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_53),
.B(n_23),
.C(n_13),
.D(n_15),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_23),
.CON(n_78),
.SN(n_78)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_17),
.C(n_48),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_27),
.C(n_37),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_58),
.C(n_37),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_69),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_85),
.C(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_83),
.B1(n_71),
.B2(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_52),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_74),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_69),
.B(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_77),
.B(n_2),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_78),
.B1(n_33),
.B2(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_79),
.B1(n_77),
.B2(n_33),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_31),
.B1(n_35),
.B2(n_13),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_31),
.B1(n_13),
.B2(n_12),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_95),
.B1(n_93),
.B2(n_96),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_91),
.C(n_12),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_1),
.B(n_2),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_12),
.A3(n_15),
.B1(n_31),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.C(n_8),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_100),
.B(n_4),
.C(n_7),
.Y(n_105)
);

AOI321xp33_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.A3(n_1),
.B1(n_4),
.B2(n_8),
.C(n_24),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);


endmodule