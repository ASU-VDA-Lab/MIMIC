module fake_ibex_559_n_571 (n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_54, n_19, n_571);

input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_571;

wire n_151;
wire n_85;
wire n_507;
wire n_540;
wire n_395;
wire n_84;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_510;
wire n_193;
wire n_418;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_86;
wire n_255;
wire n_175;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_545;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_88;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_531;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_187;
wire n_105;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_89;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_523;
wire n_116;
wire n_370;
wire n_431;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_543;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_536;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_263;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_439;
wire n_433;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_365;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_283;
wire n_397;
wire n_366;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_238;
wire n_214;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_83;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_8),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_26),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_28),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_56),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_10),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_9),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_17),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_69),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_51),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_5),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_5),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_31),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_6),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_0),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_19),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_13),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_53),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_65),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_12),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_37),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_34),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_60),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_20),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_45),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_23),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_36),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_46),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_7),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_0),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_32),
.B(n_80),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_1),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_2),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_3),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_33),
.B(n_79),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_4),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

OAI22x1_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx11_ASAP7_75t_R g165 ( 
.A(n_115),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_86),
.B(n_41),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_85),
.A2(n_39),
.B(n_77),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_89),
.A2(n_38),
.B(n_72),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_98),
.A2(n_43),
.B(n_71),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_12),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_87),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

BUFx8_ASAP7_75t_SL g182 ( 
.A(n_117),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_14),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_15),
.B(n_16),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_21),
.B(n_24),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_107),
.B(n_29),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_82),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_108),
.B(n_30),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_67),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_113),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g205 ( 
.A1(n_149),
.A2(n_114),
.B(n_139),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_112),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_106),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_175),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_125),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_192),
.B(n_105),
.Y(n_230)
);

AO21x2_ASAP7_75t_L g231 ( 
.A1(n_149),
.A2(n_119),
.B(n_118),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_151),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_191),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

AO21x2_ASAP7_75t_L g241 ( 
.A1(n_152),
.A2(n_116),
.B(n_133),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_201),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

OR2x6_ASAP7_75t_L g252 ( 
.A(n_163),
.B(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_143),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_170),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_144),
.B(n_124),
.Y(n_259)
);

CKINVDCx6p67_ASAP7_75t_R g260 ( 
.A(n_180),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_198),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_198),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_162),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_144),
.Y(n_266)
);

BUFx6f_ASAP7_75t_SL g267 ( 
.A(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_220),
.B(n_199),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_209),
.A2(n_162),
.B1(n_196),
.B2(n_181),
.Y(n_270)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_183),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_220),
.B(n_197),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_184),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_240),
.B(n_195),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_184),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_236),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_218),
.B(n_157),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

BUFx8_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_179),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_206),
.B(n_179),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_177),
.Y(n_288)
);

OR2x6_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_163),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_232),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_206),
.B(n_194),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_213),
.B(n_145),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_205),
.A2(n_166),
.B1(n_160),
.B2(n_145),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_145),
.C(n_160),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_209),
.A2(n_202),
.B1(n_200),
.B2(n_154),
.Y(n_296)
);

BUFx6f_ASAP7_75t_SL g297 ( 
.A(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_213),
.B(n_160),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_227),
.B(n_190),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_227),
.B(n_190),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_231),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_210),
.B(n_189),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_241),
.B(n_189),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_203),
.B(n_165),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_209),
.B(n_177),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_241),
.B(n_189),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_211),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_L g311 ( 
.A(n_212),
.B(n_171),
.C(n_168),
.Y(n_311)
);

BUFx6f_ASAP7_75t_SL g312 ( 
.A(n_243),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_168),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_298),
.B(n_304),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_263),
.A2(n_224),
.B1(n_217),
.B2(n_226),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_221),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_225),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_237),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_226),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_225),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_238),
.B(n_233),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_208),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_223),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_270),
.B(n_219),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_216),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_264),
.A2(n_300),
.B(n_299),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_214),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_273),
.B(n_207),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_245),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_312),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

NOR2x1_ASAP7_75t_L g344 ( 
.A(n_265),
.B(n_246),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_229),
.B(n_255),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_303),
.B(n_311),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_289),
.A2(n_246),
.B1(n_242),
.B2(n_253),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_296),
.B(n_244),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_291),
.B(n_275),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_294),
.A2(n_288),
.B(n_278),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_306),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_248),
.Y(n_359)
);

BUFx4_ASAP7_75t_SL g360 ( 
.A(n_325),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_297),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_339),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_277),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

AOI21xp33_ASAP7_75t_L g365 ( 
.A1(n_328),
.A2(n_287),
.B(n_312),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_150),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_47),
.Y(n_369)
);

AND3x4_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_49),
.C(n_52),
.Y(n_370)
);

AO21x2_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_257),
.B(n_256),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

NAND2x1p5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_251),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_331),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_332),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

AND3x1_ASAP7_75t_SL g377 ( 
.A(n_358),
.B(n_326),
.C(n_342),
.Y(n_377)
);

OAI21x1_ASAP7_75t_SL g378 ( 
.A1(n_315),
.A2(n_349),
.B(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_336),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_345),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

OAI22x1_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_352),
.B1(n_356),
.B2(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

BUFx4f_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_325),
.Y(n_387)
);

AO21x1_ASAP7_75t_L g388 ( 
.A1(n_357),
.A2(n_307),
.B(n_301),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_314),
.A2(n_298),
.B(n_292),
.Y(n_389)
);

NAND2x1p5_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_323),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_272),
.Y(n_392)
);

INVx3_ASAP7_75t_SL g393 ( 
.A(n_342),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_314),
.A2(n_330),
.B(n_348),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_337),
.B(n_272),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_328),
.A2(n_209),
.B1(n_289),
.B2(n_234),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_319),
.A2(n_320),
.B1(n_316),
.B2(n_317),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_272),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_272),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

AO31x2_ASAP7_75t_L g401 ( 
.A1(n_346),
.A2(n_322),
.A3(n_314),
.B(n_309),
.Y(n_401)
);

AO21x2_ASAP7_75t_L g402 ( 
.A1(n_348),
.A2(n_346),
.B(n_357),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_272),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_314),
.A2(n_330),
.B(n_348),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_318),
.B(n_272),
.Y(n_405)
);

AO31x2_ASAP7_75t_L g406 ( 
.A1(n_346),
.A2(n_322),
.A3(n_314),
.B(n_309),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_272),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_337),
.B(n_272),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g411 ( 
.A1(n_346),
.A2(n_309),
.B(n_304),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_328),
.A2(n_209),
.B1(n_289),
.B2(n_234),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_325),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_337),
.B(n_272),
.Y(n_416)
);

INVx3_ASAP7_75t_SL g417 ( 
.A(n_387),
.Y(n_417)
);

NAND2x1p5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_364),
.Y(n_418)
);

NAND2x1p5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_364),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_360),
.Y(n_420)
);

OAI21x1_ASAP7_75t_SL g421 ( 
.A1(n_397),
.A2(n_378),
.B(n_374),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_410),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_409),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_416),
.Y(n_428)
);

AO21x2_ASAP7_75t_L g429 ( 
.A1(n_394),
.A2(n_388),
.B(n_411),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_362),
.A2(n_361),
.B1(n_375),
.B2(n_415),
.Y(n_430)
);

BUFx2_ASAP7_75t_SL g431 ( 
.A(n_414),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_412),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

INVx3_ASAP7_75t_SL g436 ( 
.A(n_407),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_393),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_389),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_396),
.A2(n_413),
.B1(n_385),
.B2(n_400),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

NOR2x1_ASAP7_75t_R g442 ( 
.A(n_376),
.B(n_380),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_373),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_363),
.Y(n_446)
);

OAI211xp5_ASAP7_75t_SL g447 ( 
.A1(n_396),
.A2(n_413),
.B(n_365),
.C(n_379),
.Y(n_447)
);

BUFx2_ASAP7_75t_R g448 ( 
.A(n_402),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_382),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g452 ( 
.A1(n_371),
.A2(n_402),
.B(n_366),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_401),
.A2(n_406),
.B(n_377),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_396),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_414),
.Y(n_458)
);

AO21x2_ASAP7_75t_L g459 ( 
.A1(n_394),
.A2(n_348),
.B(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

BUFx12f_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_432),
.Y(n_463)
);

OAI22xp33_ASAP7_75t_L g464 ( 
.A1(n_455),
.A2(n_440),
.B1(n_424),
.B2(n_422),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_421),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_455),
.A2(n_447),
.B1(n_430),
.B2(n_457),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_423),
.A2(n_462),
.B1(n_460),
.B2(n_428),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_433),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_459),
.Y(n_472)
);

INVx4_ASAP7_75t_SL g473 ( 
.A(n_441),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_461),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_447),
.A2(n_430),
.B1(n_454),
.B2(n_449),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_435),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_456),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_441),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_450),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_449),
.A2(n_431),
.B1(n_454),
.B2(n_420),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_437),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_483),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_483),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_485),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_445),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_464),
.A2(n_450),
.B1(n_446),
.B2(n_443),
.Y(n_492)
);

OAI221xp5_ASAP7_75t_SL g493 ( 
.A1(n_466),
.A2(n_438),
.B1(n_442),
.B2(n_448),
.C(n_458),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_429),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_452),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_467),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_465),
.B(n_475),
.Y(n_501)
);

INVx3_ASAP7_75t_SL g502 ( 
.A(n_473),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_469),
.A2(n_443),
.B1(n_437),
.B2(n_438),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_472),
.A2(n_450),
.B1(n_446),
.B2(n_461),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_488),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_496),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_481),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_489),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_478),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_501),
.A2(n_487),
.B1(n_484),
.B2(n_482),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_479),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_489),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_514),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_498),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_505),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_493),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_497),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_495),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_506),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_501),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_517),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_519),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_523),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_526),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_507),
.Y(n_532)
);

AOI21xp33_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_486),
.B(n_491),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_522),
.Y(n_534)
);

OAI32xp33_ASAP7_75t_L g535 ( 
.A1(n_520),
.A2(n_492),
.A3(n_506),
.B1(n_511),
.B2(n_508),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_534),
.A2(n_491),
.B1(n_522),
.B2(n_524),
.Y(n_536)
);

AOI21xp33_ASAP7_75t_L g537 ( 
.A1(n_535),
.A2(n_486),
.B(n_525),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_518),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_529),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_533),
.A2(n_535),
.B(n_527),
.C(n_528),
.Y(n_540)
);

AO22x1_ASAP7_75t_L g541 ( 
.A1(n_532),
.A2(n_524),
.B1(n_502),
.B2(n_521),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_474),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_524),
.B1(n_521),
.B2(n_501),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_540),
.A2(n_503),
.B(n_513),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_SL g546 ( 
.A(n_536),
.B(n_503),
.C(n_504),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_539),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_544),
.B(n_538),
.Y(n_548)
);

AOI221xp5_ASAP7_75t_L g549 ( 
.A1(n_545),
.A2(n_536),
.B1(n_529),
.B2(n_541),
.C(n_542),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_546),
.A2(n_543),
.B(n_465),
.Y(n_550)
);

NAND5xp2_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_474),
.C(n_418),
.D(n_419),
.E(n_481),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_547),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_552),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_552),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_550),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_553),
.A2(n_474),
.B1(n_417),
.B2(n_436),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_556),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_476),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_558),
.Y(n_559)
);

XOR2x1_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_417),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_560),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_559),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_562),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_562),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_484),
.Y(n_565)
);

AOI221xp5_ASAP7_75t_L g566 ( 
.A1(n_563),
.A2(n_478),
.B1(n_476),
.B2(n_484),
.C(n_426),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_564),
.C(n_565),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_568),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_569),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_502),
.B1(n_480),
.B2(n_482),
.Y(n_571)
);


endmodule