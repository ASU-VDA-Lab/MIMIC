module fake_aes_1468_n_1293 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1293);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1293;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVxp67_ASAP7_75t_L g284 ( .A(n_90), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_49), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_234), .Y(n_286) );
INVxp33_ASAP7_75t_SL g287 ( .A(n_71), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_249), .Y(n_288) );
INVxp33_ASAP7_75t_L g289 ( .A(n_23), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_146), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_279), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_62), .Y(n_294) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_63), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_217), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_208), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_83), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_170), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_99), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_87), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_267), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_102), .Y(n_305) );
CKINVDCx14_ASAP7_75t_R g306 ( .A(n_232), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_172), .B(n_9), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_228), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_127), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_199), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_6), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_255), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_86), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_24), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_25), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_0), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_84), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_152), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_49), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_88), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_183), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_103), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_220), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_105), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_171), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_200), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_0), .Y(n_327) );
NOR2xp67_ASAP7_75t_L g328 ( .A(n_75), .B(n_259), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_258), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_244), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_270), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_213), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_18), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_155), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_63), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_191), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_271), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_116), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_18), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_30), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_21), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_168), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_202), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_261), .B(n_39), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_166), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_65), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_37), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_242), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_69), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_134), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_44), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_273), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_100), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_128), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_32), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_178), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_32), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_264), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_198), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_29), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_28), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_201), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_173), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_182), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_238), .Y(n_365) );
INVxp33_ASAP7_75t_SL g366 ( .A(n_145), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_122), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_189), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_75), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_55), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_275), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_55), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_120), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_212), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_109), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_14), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_248), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_141), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_176), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_138), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_13), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_150), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_108), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_68), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_265), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_222), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_97), .B(n_34), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_121), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_268), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_38), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_133), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_94), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_177), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_5), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_257), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_154), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_80), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_184), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_231), .B(n_175), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_278), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_276), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_113), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_79), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_25), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_246), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_62), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_2), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_64), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_91), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_43), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_112), .Y(n_411) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_266), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_272), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_211), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_180), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_10), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_16), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_92), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_52), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_239), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_95), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_106), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_110), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_1), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_174), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_21), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_282), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_148), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_48), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_251), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_107), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_6), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_327), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_327), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_291), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_289), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_386), .B(n_1), .Y(n_437) );
AND3x2_ASAP7_75t_L g438 ( .A(n_354), .B(n_2), .C(n_3), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_288), .B(n_3), .Y(n_439) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_288), .A2(n_4), .B(n_5), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_291), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_291), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_341), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_341), .B(n_4), .Y(n_444) );
INVxp33_ASAP7_75t_SL g445 ( .A(n_300), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_286), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_291), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_289), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_322), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_322), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_348), .B(n_7), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_348), .B(n_352), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_290), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_296), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_285), .B(n_7), .Y(n_455) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_352), .A2(n_8), .B(n_9), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_322), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_297), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_299), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_300), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_322), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_306), .B(n_412), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_303), .Y(n_464) );
AOI22x1_ASAP7_75t_SL g465 ( .A1(n_349), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_355), .B(n_11), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_314), .B(n_12), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_451), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_441), .Y(n_471) );
BUFx8_ASAP7_75t_SL g472 ( .A(n_437), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_440), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_437), .A2(n_287), .B1(n_335), .B2(n_333), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_440), .Y(n_475) );
AND2x6_ASAP7_75t_L g476 ( .A(n_437), .B(n_326), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_436), .B(n_284), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_463), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_436), .B(n_306), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_448), .B(n_412), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_448), .B(n_329), .Y(n_487) );
BUFx10_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_435), .Y(n_489) );
BUFx10_ASAP7_75t_L g490 ( .A(n_437), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_463), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_445), .B(n_363), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_451), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_463), .B(n_349), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_440), .Y(n_495) );
INVx4_ASAP7_75t_L g496 ( .A(n_451), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_451), .B(n_315), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_435), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_451), .A2(n_316), .B1(n_346), .B2(n_319), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_460), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_442), .Y(n_501) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
INVx4_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_460), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_465), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_446), .B(n_410), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_435), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
OR2x6_ASAP7_75t_L g509 ( .A(n_444), .B(n_307), .Y(n_509) );
INVx4_ASAP7_75t_SL g510 ( .A(n_444), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_444), .A2(n_347), .B1(n_357), .B2(n_351), .Y(n_511) );
AND2x2_ASAP7_75t_SL g512 ( .A(n_456), .B(n_399), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_433), .Y(n_513) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_456), .B(n_305), .C(n_304), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_446), .B(n_385), .Y(n_515) );
INVx4_ASAP7_75t_SL g516 ( .A(n_452), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_452), .B(n_293), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_482), .B(n_453), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_482), .B(n_453), .Y(n_519) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_502), .B(n_456), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_506), .A2(n_469), .B(n_455), .C(n_458), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_484), .B(n_454), .Y(n_522) );
AND3x1_ASAP7_75t_L g523 ( .A(n_474), .B(n_467), .C(n_465), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_476), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_516), .Y(n_525) );
AO22x1_ASAP7_75t_L g526 ( .A1(n_487), .A2(n_287), .B1(n_366), .B2(n_390), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_484), .B(n_454), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_474), .A2(n_292), .B1(n_353), .B2(n_312), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_516), .Y(n_529) );
O2A1O1Ixp5_ASAP7_75t_L g530 ( .A1(n_502), .A2(n_439), .B(n_469), .C(n_455), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_502), .B(n_452), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_478), .B(n_458), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_515), .B(n_459), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_514), .A2(n_464), .B(n_459), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_510), .Y(n_535) );
NOR2x1p5_ASAP7_75t_L g536 ( .A(n_506), .B(n_390), .Y(n_536) );
AND2x2_ASAP7_75t_SL g537 ( .A(n_503), .B(n_456), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_487), .B(n_464), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_500), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_504), .A2(n_467), .B1(n_292), .B2(n_353), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_481), .B(n_491), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_476), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_510), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_510), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_472), .Y(n_545) );
NOR2x2_ASAP7_75t_L g546 ( .A(n_509), .B(n_312), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_504), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_481), .A2(n_392), .B1(n_420), .B2(n_380), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_510), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_488), .B(n_452), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_494), .B(n_408), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_510), .B(n_438), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_488), .B(n_309), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_509), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_496), .B(n_433), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_509), .B(n_438), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_503), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_513), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_509), .A2(n_392), .B1(n_420), .B2(n_380), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_488), .B(n_317), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_492), .B(n_408), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_503), .B(n_456), .Y(n_562) );
CKINVDCx16_ASAP7_75t_R g563 ( .A(n_505), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_497), .A2(n_366), .B1(n_432), .B2(n_295), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_496), .B(n_433), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_503), .B(n_360), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_497), .B(n_434), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_490), .B(n_339), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_497), .B(n_434), .Y(n_569) );
AOI22x1_ASAP7_75t_L g570 ( .A1(n_473), .A2(n_434), .B1(n_423), .B2(n_379), .Y(n_570) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_517), .B(n_443), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_511), .B(n_294), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_497), .B(n_476), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_473), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_476), .B(n_434), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_470), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_512), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_470), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_476), .B(n_434), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_470), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_470), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_499), .A2(n_417), .B1(n_340), .B2(n_424), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_493), .A2(n_443), .B(n_361), .C(n_370), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_490), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_475), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_476), .B(n_298), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_490), .B(n_320), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_493), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_493), .A2(n_372), .B1(n_376), .B2(n_369), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_493), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_512), .B(n_298), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_475), .B(n_414), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_483), .B(n_301), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_483), .B(n_321), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_485), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_485), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_486), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_514), .A2(n_325), .B(n_323), .Y(n_599) );
NOR2x2_ASAP7_75t_L g600 ( .A(n_471), .B(n_379), .Y(n_600) );
OAI22xp5_ASAP7_75t_SL g601 ( .A1(n_486), .A2(n_394), .B1(n_397), .B2(n_381), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_495), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_547), .B(n_495), .Y(n_603) );
INVx2_ASAP7_75t_SL g604 ( .A(n_539), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_554), .A2(n_508), .B1(n_404), .B2(n_406), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_521), .A2(n_593), .B(n_530), .C(n_534), .Y(n_606) );
BUFx3_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_575), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_595), .A2(n_508), .B(n_498), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_556), .B(n_403), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_564), .A2(n_419), .B1(n_426), .B2(n_416), .C(n_407), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_524), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_524), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_595), .A2(n_498), .B(n_388), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_556), .B(n_301), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_538), .A2(n_429), .B(n_331), .C(n_332), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_600), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_584), .A2(n_338), .B(n_342), .C(n_330), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_518), .B(n_308), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_536), .A2(n_308), .B1(n_364), .B2(n_310), .Y(n_621) );
NAND2xp33_ASAP7_75t_SL g622 ( .A(n_559), .B(n_310), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_519), .B(n_364), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_563), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_584), .A2(n_343), .B(n_350), .C(n_345), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_596), .A2(n_391), .B1(n_411), .B2(n_336), .Y(n_626) );
BUFx8_ASAP7_75t_SL g627 ( .A(n_552), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_522), .B(n_371), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_541), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_548), .B(n_371), .Y(n_630) );
O2A1O1Ixp5_ASAP7_75t_L g631 ( .A1(n_530), .A2(n_387), .B(n_344), .C(n_423), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_SL g632 ( .A1(n_599), .A2(n_358), .B(n_362), .C(n_356), .Y(n_632) );
AND2x2_ASAP7_75t_SL g633 ( .A(n_552), .B(n_311), .Y(n_633) );
INVx11_ASAP7_75t_L g634 ( .A(n_546), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_574), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_527), .B(n_378), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_597), .A2(n_328), .B1(n_367), .B2(n_365), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_532), .A2(n_374), .B(n_375), .C(n_368), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_571), .A2(n_384), .B1(n_311), .B2(n_382), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_573), .A2(n_389), .B(n_398), .C(n_377), .Y(n_641) );
HAxp5_ASAP7_75t_L g642 ( .A(n_523), .B(n_12), .CON(n_642), .SN(n_642) );
O2A1O1Ixp33_ASAP7_75t_SL g643 ( .A1(n_576), .A2(n_402), .B(n_405), .C(n_400), .Y(n_643) );
AOI21x1_ASAP7_75t_L g644 ( .A1(n_580), .A2(n_498), .B(n_477), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_557), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_598), .A2(n_413), .B(n_409), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_571), .A2(n_384), .B1(n_311), .B2(n_421), .Y(n_647) );
AOI21x1_ASAP7_75t_L g648 ( .A1(n_553), .A2(n_477), .B(n_471), .Y(n_648) );
OA22x2_ASAP7_75t_L g649 ( .A1(n_540), .A2(n_393), .B1(n_401), .B2(n_383), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_602), .A2(n_428), .B(n_425), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_568), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_566), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_531), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_589), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_577), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_564), .B(n_383), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_561), .B(n_401), .C(n_393), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_553), .A2(n_430), .B(n_480), .Y(n_658) );
NOR2xp67_ASAP7_75t_SL g659 ( .A(n_542), .B(n_415), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_542), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_579), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_581), .Y(n_662) );
NOR2xp33_ASAP7_75t_R g663 ( .A(n_592), .B(n_415), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_531), .A2(n_313), .B(n_395), .C(n_302), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_571), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_582), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_526), .B(n_318), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_558), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_533), .A2(n_326), .B(n_337), .C(n_334), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_551), .A2(n_334), .B(n_359), .C(n_337), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_566), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g673 ( .A(n_583), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_572), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_601), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_571), .A2(n_384), .B1(n_373), .B2(n_359), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_585), .B(n_324), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_590), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_578), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_560), .A2(n_501), .B(n_396), .Y(n_680) );
BUFx4f_ASAP7_75t_L g681 ( .A(n_578), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_567), .A2(n_396), .B(n_418), .C(n_373), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_528), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_578), .A2(n_384), .B1(n_418), .B2(n_447), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_560), .A2(n_449), .B(n_447), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_535), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_520), .B(n_422), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_569), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_544), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_555), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_550), .A2(n_594), .B1(n_520), .B2(n_537), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_587), .B(n_427), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_549), .B(n_431), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_550), .B(n_13), .Y(n_694) );
INVx3_ASAP7_75t_L g695 ( .A(n_529), .Y(n_695) );
NOR2xp33_ASAP7_75t_R g696 ( .A(n_525), .B(n_14), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_537), .A2(n_449), .B1(n_457), .B2(n_447), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_588), .A2(n_449), .B(n_447), .Y(n_698) );
BUFx4f_ASAP7_75t_L g699 ( .A(n_543), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_562), .B(n_449), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_528), .A2(n_468), .B1(n_466), .B2(n_462), .Y(n_701) );
AOI21x1_ASAP7_75t_L g702 ( .A1(n_588), .A2(n_462), .B(n_457), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_562), .B(n_457), .Y(n_703) );
INVx4_ASAP7_75t_L g704 ( .A(n_549), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_565), .B(n_457), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_570), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_554), .A2(n_462), .B1(n_468), .B2(n_466), .Y(n_707) );
INVx3_ASAP7_75t_L g708 ( .A(n_529), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_575), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_595), .A2(n_462), .B(n_479), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_SL g711 ( .A1(n_599), .A2(n_468), .B(n_489), .C(n_479), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_539), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_554), .A2(n_435), .B1(n_450), .B2(n_461), .Y(n_713) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_524), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_539), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_554), .B(n_435), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_554), .B(n_435), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_554), .B(n_435), .Y(n_718) );
CKINVDCx6p67_ASAP7_75t_R g719 ( .A(n_539), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_539), .B(n_15), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_595), .A2(n_489), .B(n_479), .Y(n_721) );
BUFx3_ASAP7_75t_L g722 ( .A(n_539), .Y(n_722) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_524), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_547), .B(n_15), .Y(n_724) );
O2A1O1Ixp33_ASAP7_75t_L g725 ( .A1(n_538), .A2(n_16), .B(n_17), .C(n_19), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_547), .B(n_17), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_595), .A2(n_489), .B(n_479), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_638), .A2(n_461), .B(n_450), .C(n_507), .Y(n_728) );
BUFx10_ASAP7_75t_L g729 ( .A(n_604), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_609), .A2(n_507), .B(n_489), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_608), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_619), .A2(n_461), .B(n_450), .C(n_507), .Y(n_732) );
AO21x1_ASAP7_75t_L g733 ( .A1(n_697), .A2(n_461), .B(n_450), .Y(n_733) );
INVx6_ASAP7_75t_L g734 ( .A(n_722), .Y(n_734) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_612), .A2(n_641), .B(n_617), .C(n_625), .Y(n_735) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_665), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_606), .A2(n_19), .B(n_20), .C(n_22), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_632), .A2(n_461), .B(n_450), .Y(n_738) );
O2A1O1Ixp33_ASAP7_75t_SL g739 ( .A1(n_711), .A2(n_158), .B(n_283), .C(n_281), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_719), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_629), .B(n_20), .Y(n_741) );
NOR2xp33_ASAP7_75t_R g742 ( .A(n_624), .B(n_22), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_671), .A2(n_461), .B(n_507), .C(n_26), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g744 ( .A(n_618), .B(n_23), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_706), .A2(n_507), .B(n_461), .Y(n_745) );
BUFx3_ASAP7_75t_L g746 ( .A(n_715), .Y(n_746) );
O2A1O1Ixp5_ASAP7_75t_L g747 ( .A1(n_631), .A2(n_461), .B(n_159), .C(n_160), .Y(n_747) );
INVx5_ASAP7_75t_L g748 ( .A(n_627), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_669), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_678), .B(n_24), .Y(n_750) );
INVx1_ASAP7_75t_SL g751 ( .A(n_712), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_618), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_683), .B(n_27), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_633), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_721), .A2(n_89), .B(n_85), .Y(n_755) );
BUFx12f_ASAP7_75t_SL g756 ( .A(n_610), .Y(n_756) );
AO31x2_ASAP7_75t_L g757 ( .A1(n_697), .A2(n_27), .A3(n_28), .B(n_29), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_651), .B(n_30), .Y(n_758) );
O2A1O1Ixp33_ASAP7_75t_SL g759 ( .A1(n_652), .A2(n_162), .B(n_277), .C(n_269), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_622), .A2(n_31), .B1(n_33), .B2(n_34), .Y(n_760) );
AND2x6_ASAP7_75t_L g761 ( .A(n_652), .B(n_31), .Y(n_761) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_672), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_649), .A2(n_33), .B1(n_35), .B2(n_36), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_649), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_700), .A2(n_96), .B(n_93), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_637), .A2(n_39), .B(n_40), .C(n_41), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_656), .B(n_40), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_630), .B(n_41), .Y(n_768) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_672), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_607), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_611), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_700), .A2(n_101), .B(n_98), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_703), .A2(n_111), .B(n_104), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_703), .A2(n_115), .B(n_114), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_656), .B(n_42), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_616), .B(n_42), .Y(n_776) );
NAND2x1p5_ASAP7_75t_L g777 ( .A(n_681), .B(n_44), .Y(n_777) );
BUFx3_ASAP7_75t_L g778 ( .A(n_610), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_653), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_640), .Y(n_780) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_665), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_694), .Y(n_782) );
AO31x2_ASAP7_75t_L g783 ( .A1(n_637), .A2(n_45), .A3(n_46), .B(n_47), .Y(n_783) );
AND3x2_ASAP7_75t_L g784 ( .A(n_634), .B(n_720), .C(n_667), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_709), .A2(n_118), .B(n_117), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_688), .Y(n_786) );
OAI22xp5_ASAP7_75t_SL g787 ( .A1(n_675), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_787) );
CKINVDCx8_ASAP7_75t_R g788 ( .A(n_673), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_674), .A2(n_48), .B1(n_50), .B2(n_51), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_645), .Y(n_790) );
AO31x2_ASAP7_75t_L g791 ( .A1(n_684), .A2(n_50), .A3(n_51), .B(n_52), .Y(n_791) );
INVx1_ASAP7_75t_SL g792 ( .A(n_696), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_635), .A2(n_53), .B1(n_54), .B2(n_56), .Y(n_793) );
NOR2xp33_ASAP7_75t_SL g794 ( .A(n_681), .B(n_53), .Y(n_794) );
O2A1O1Ixp33_ASAP7_75t_SL g795 ( .A1(n_605), .A2(n_670), .B(n_717), .C(n_716), .Y(n_795) );
NOR2x1_ASAP7_75t_SL g796 ( .A(n_704), .B(n_54), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_603), .A2(n_56), .B(n_57), .C(n_58), .Y(n_797) );
OR2x6_ASAP7_75t_L g798 ( .A(n_725), .B(n_57), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_SL g799 ( .A1(n_718), .A2(n_187), .B(n_263), .C(n_262), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_654), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_727), .A2(n_185), .B(n_256), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_642), .B(n_58), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_620), .B(n_59), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_623), .B(n_59), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_705), .A2(n_186), .B(n_254), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_655), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_628), .B(n_60), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_661), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_635), .A2(n_60), .B1(n_61), .B2(n_64), .Y(n_809) );
INVx8_ASAP7_75t_L g810 ( .A(n_613), .Y(n_810) );
AO32x2_ASAP7_75t_L g811 ( .A1(n_684), .A2(n_61), .A3(n_65), .B1(n_66), .B2(n_67), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_705), .A2(n_188), .B(n_253), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_662), .Y(n_813) );
NAND3xp33_ASAP7_75t_SL g814 ( .A(n_664), .B(n_66), .C(n_67), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_621), .B(n_68), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_701), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_666), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_665), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_690), .A2(n_190), .B(n_252), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_657), .B(n_69), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_SL g821 ( .A1(n_693), .A2(n_181), .B(n_247), .C(n_245), .Y(n_821) );
AO31x2_ASAP7_75t_L g822 ( .A1(n_713), .A2(n_70), .A3(n_71), .B(n_72), .Y(n_822) );
AO31x2_ASAP7_75t_L g823 ( .A1(n_713), .A2(n_70), .A3(n_72), .B(n_73), .Y(n_823) );
O2A1O1Ixp33_ASAP7_75t_L g824 ( .A1(n_626), .A2(n_73), .B(n_74), .C(n_76), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_668), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_644), .A2(n_192), .B(n_243), .Y(n_826) );
O2A1O1Ixp33_ASAP7_75t_L g827 ( .A1(n_626), .A2(n_74), .B(n_76), .C(n_77), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_636), .A2(n_77), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_724), .A2(n_78), .B1(n_81), .B2(n_82), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_615), .A2(n_687), .B(n_692), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_643), .A2(n_82), .B(n_83), .C(n_119), .Y(n_831) );
AND2x4_ASAP7_75t_L g832 ( .A(n_704), .B(n_123), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_691), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_833) );
A2O1A1Ixp33_ASAP7_75t_L g834 ( .A1(n_646), .A2(n_129), .B(n_130), .C(n_131), .Y(n_834) );
O2A1O1Ixp33_ASAP7_75t_SL g835 ( .A1(n_682), .A2(n_132), .B(n_135), .C(n_136), .Y(n_835) );
AO32x2_ASAP7_75t_L g836 ( .A1(n_707), .A2(n_137), .A3(n_139), .B1(n_140), .B2(n_142), .Y(n_836) );
AO32x2_ASAP7_75t_L g837 ( .A1(n_707), .A2(n_143), .A3(n_144), .B1(n_147), .B2(n_149), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_726), .A2(n_151), .B1(n_153), .B2(n_156), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_663), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_686), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_650), .A2(n_157), .B1(n_161), .B2(n_163), .C(n_164), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_687), .A2(n_165), .B1(n_167), .B2(n_169), .Y(n_842) );
AO31x2_ASAP7_75t_L g843 ( .A1(n_710), .A2(n_179), .A3(n_193), .B(n_194), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_677), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_L g845 ( .A1(n_658), .A2(n_195), .B(n_196), .C(n_197), .Y(n_845) );
INVx2_ASAP7_75t_SL g846 ( .A(n_699), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_679), .Y(n_847) );
O2A1O1Ixp5_ASAP7_75t_L g848 ( .A1(n_659), .A2(n_203), .B(n_204), .C(n_205), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_689), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g850 ( .A1(n_680), .A2(n_206), .B(n_207), .Y(n_850) );
OAI21x1_ASAP7_75t_SL g851 ( .A1(n_648), .A2(n_209), .B(n_210), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_679), .A2(n_214), .B1(n_215), .B2(n_216), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_695), .A2(n_218), .B(n_219), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g854 ( .A1(n_702), .A2(n_221), .B(n_223), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_676), .A2(n_225), .B1(n_226), .B2(n_227), .C(n_229), .Y(n_855) );
INVx6_ASAP7_75t_L g856 ( .A(n_613), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_639), .A2(n_230), .B1(n_233), .B2(n_235), .C(n_236), .Y(n_857) );
AOI221x1_ASAP7_75t_L g858 ( .A1(n_685), .A2(n_237), .B1(n_240), .B2(n_241), .C(n_280), .Y(n_858) );
OAI21xp5_ASAP7_75t_L g859 ( .A1(n_698), .A2(n_695), .B(n_708), .Y(n_859) );
OAI21xp5_ASAP7_75t_L g860 ( .A1(n_708), .A2(n_647), .B(n_699), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_614), .Y(n_861) );
OAI21x1_ASAP7_75t_L g862 ( .A1(n_614), .A2(n_660), .B(n_714), .Y(n_862) );
NAND2xp5_ASAP7_75t_SL g863 ( .A(n_723), .B(n_547), .Y(n_863) );
AOI221x1_ASAP7_75t_L g864 ( .A1(n_723), .A2(n_697), .B1(n_606), .B2(n_637), .C(n_706), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_733), .A2(n_738), .B(n_851), .Y(n_865) );
OAI21xp5_ASAP7_75t_L g866 ( .A1(n_747), .A2(n_864), .B(n_743), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_746), .Y(n_867) );
INVx3_ASAP7_75t_L g868 ( .A(n_810), .Y(n_868) );
AOI21x1_ASAP7_75t_L g869 ( .A1(n_745), .A2(n_826), .B(n_858), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_740), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_786), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_782), .B(n_749), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_859), .A2(n_739), .B(n_835), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_808), .Y(n_874) );
OA21x2_ASAP7_75t_L g875 ( .A1(n_854), .A2(n_819), .B(n_848), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_816), .A2(n_832), .B1(n_754), .B2(n_798), .Y(n_876) );
AO31x2_ASAP7_75t_L g877 ( .A1(n_732), .A2(n_728), .A3(n_833), .B(n_845), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_731), .Y(n_878) );
A2O1A1Ixp33_ASAP7_75t_L g879 ( .A1(n_735), .A2(n_737), .B(n_775), .C(n_820), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_768), .B(n_753), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_803), .B(n_779), .Y(n_881) );
AND2x4_ASAP7_75t_SL g882 ( .A(n_729), .B(n_762), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_825), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_751), .B(n_750), .Y(n_884) );
OR2x2_ASAP7_75t_L g885 ( .A(n_752), .B(n_778), .Y(n_885) );
OA21x2_ASAP7_75t_L g886 ( .A1(n_850), .A2(n_801), .B(n_755), .Y(n_886) );
CKINVDCx11_ASAP7_75t_R g887 ( .A(n_729), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_802), .B(n_734), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_815), .A2(n_758), .B1(n_776), .B2(n_756), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_767), .B(n_769), .Y(n_890) );
OAI211xp5_ASAP7_75t_SL g891 ( .A1(n_763), .A2(n_764), .B(n_788), .C(n_824), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_807), .B(n_741), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_804), .B(n_806), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_748), .Y(n_894) );
CKINVDCx6p67_ASAP7_75t_R g895 ( .A(n_748), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_813), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_817), .B(n_771), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_805), .A2(n_812), .B(n_773), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_765), .A2(n_772), .B(n_774), .Y(n_899) );
OA21x2_ASAP7_75t_L g900 ( .A1(n_834), .A2(n_785), .B(n_853), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_780), .B(n_800), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_798), .A2(n_814), .B1(n_787), .B2(n_792), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_849), .B(n_790), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_832), .A2(n_777), .B1(n_760), .B2(n_829), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_844), .B(n_784), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_734), .B(n_744), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_761), .A2(n_770), .B1(n_828), .B2(n_839), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_796), .Y(n_908) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_761), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_846), .B(n_827), .Y(n_910) );
BUFx8_ASAP7_75t_L g911 ( .A(n_761), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_759), .A2(n_831), .B(n_860), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_761), .Y(n_913) );
BUFx4f_ASAP7_75t_L g914 ( .A(n_810), .Y(n_914) );
NAND2xp5_ASAP7_75t_SL g915 ( .A(n_794), .B(n_742), .Y(n_915) );
BUFx12f_ASAP7_75t_L g916 ( .A(n_748), .Y(n_916) );
OR2x2_ASAP7_75t_L g917 ( .A(n_840), .B(n_863), .Y(n_917) );
BUFx10_ASAP7_75t_L g918 ( .A(n_856), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_766), .B(n_789), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_757), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_856), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_797), .B(n_809), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_793), .B(n_861), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_818), .A2(n_852), .B(n_842), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_847), .B(n_838), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_811), .B(n_783), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_736), .Y(n_927) );
AOI21xp5_ASAP7_75t_L g928 ( .A1(n_799), .A2(n_821), .B(n_841), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_736), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_757), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_855), .A2(n_857), .B1(n_781), .B2(n_736), .C(n_783), .Y(n_931) );
INVx3_ASAP7_75t_SL g932 ( .A(n_781), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_822), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_811), .B(n_783), .Y(n_934) );
INVxp67_ASAP7_75t_L g935 ( .A(n_781), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_811), .A2(n_791), .B1(n_822), .B2(n_823), .Y(n_936) );
NOR2x1_ASAP7_75t_SL g937 ( .A(n_836), .B(n_837), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g938 ( .A1(n_836), .A2(n_539), .B1(n_651), .B2(n_474), .C(n_683), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_843), .A2(n_795), .B(n_730), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_843), .A2(n_795), .B(n_730), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_837), .A2(n_795), .B(n_730), .Y(n_941) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_795), .A2(n_730), .B(n_706), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_751), .B(n_539), .Y(n_943) );
A2O1A1Ixp33_ASAP7_75t_L g944 ( .A1(n_735), .A2(n_737), .B(n_775), .C(n_671), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_749), .Y(n_945) );
AO31x2_ASAP7_75t_L g946 ( .A1(n_733), .A2(n_864), .A3(n_858), .B(n_697), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_751), .B(n_539), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_795), .A2(n_730), .B(n_706), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_751), .B(n_539), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_749), .Y(n_950) );
AND2x4_ASAP7_75t_L g951 ( .A(n_786), .B(n_652), .Y(n_951) );
AO21x2_ASAP7_75t_L g952 ( .A1(n_733), .A2(n_738), .B(n_851), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_751), .B(n_539), .Y(n_953) );
OAI21xp5_ASAP7_75t_L g954 ( .A1(n_830), .A2(n_606), .B(n_632), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_749), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_786), .B(n_683), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_795), .A2(n_730), .B(n_706), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_795), .A2(n_730), .B(n_706), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_786), .B(n_683), .Y(n_959) );
OAI21x1_ASAP7_75t_L g960 ( .A1(n_730), .A2(n_745), .B(n_862), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_749), .Y(n_961) );
NOR2x1_ASAP7_75t_R g962 ( .A(n_748), .B(n_740), .Y(n_962) );
INVx3_ASAP7_75t_L g963 ( .A(n_810), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_786), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_786), .B(n_683), .Y(n_965) );
AO21x2_ASAP7_75t_L g966 ( .A1(n_733), .A2(n_738), .B(n_851), .Y(n_966) );
OAI21xp5_ASAP7_75t_L g967 ( .A1(n_830), .A2(n_606), .B(n_632), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_749), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_749), .Y(n_969) );
AOI21xp5_ASAP7_75t_L g970 ( .A1(n_795), .A2(n_730), .B(n_706), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_786), .Y(n_971) );
AO31x2_ASAP7_75t_L g972 ( .A1(n_733), .A2(n_864), .A3(n_858), .B(n_697), .Y(n_972) );
A2O1A1Ixp33_ASAP7_75t_L g973 ( .A1(n_735), .A2(n_737), .B(n_775), .C(n_671), .Y(n_973) );
OAI211xp5_ASAP7_75t_SL g974 ( .A1(n_750), .A2(n_618), .B(n_474), .C(n_612), .Y(n_974) );
A2O1A1Ixp33_ASAP7_75t_L g975 ( .A1(n_735), .A2(n_737), .B(n_775), .C(n_671), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_735), .A2(n_523), .B1(n_528), .B2(n_612), .C(n_683), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_749), .Y(n_977) );
A2O1A1Ixp33_ASAP7_75t_L g978 ( .A1(n_735), .A2(n_737), .B(n_775), .C(n_671), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_795), .A2(n_730), .B(n_706), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_786), .Y(n_980) );
A2O1A1Ixp33_ASAP7_75t_L g981 ( .A1(n_735), .A2(n_737), .B(n_775), .C(n_671), .Y(n_981) );
BUFx6f_ASAP7_75t_L g982 ( .A(n_736), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_786), .B(n_683), .Y(n_983) );
AO31x2_ASAP7_75t_L g984 ( .A1(n_733), .A2(n_864), .A3(n_858), .B(n_697), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_816), .A2(n_683), .B1(n_539), .B2(n_622), .Y(n_985) );
AO21x2_ASAP7_75t_L g986 ( .A1(n_939), .A2(n_940), .B(n_941), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_876), .B(n_956), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_976), .B(n_959), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_901), .Y(n_989) );
AO21x2_ASAP7_75t_L g990 ( .A1(n_942), .A2(n_957), .B(n_948), .Y(n_990) );
INVx3_ASAP7_75t_L g991 ( .A(n_982), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_871), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_878), .B(n_897), .Y(n_993) );
AO21x2_ASAP7_75t_L g994 ( .A1(n_958), .A2(n_979), .B(n_970), .Y(n_994) );
OAI221xp5_ASAP7_75t_L g995 ( .A1(n_889), .A2(n_985), .B1(n_974), .B2(n_902), .C(n_880), .Y(n_995) );
NOR2xp33_ASAP7_75t_R g996 ( .A(n_870), .B(n_887), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_876), .A2(n_911), .B1(n_904), .B2(n_938), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_965), .B(n_983), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_897), .B(n_896), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_907), .A2(n_904), .B1(n_913), .B2(n_919), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_901), .B(n_903), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_943), .B(n_949), .Y(n_1002) );
OR2x6_ASAP7_75t_L g1003 ( .A(n_909), .B(n_908), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_903), .B(n_951), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_951), .B(n_964), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_971), .B(n_980), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_953), .B(n_945), .Y(n_1007) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_914), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_950), .B(n_955), .Y(n_1009) );
INVx4_ASAP7_75t_L g1010 ( .A(n_914), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_890), .B(n_947), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_891), .A2(n_884), .B1(n_910), .B2(n_911), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_920), .B(n_930), .Y(n_1013) );
AND2x4_ASAP7_75t_L g1014 ( .A(n_927), .B(n_982), .Y(n_1014) );
OA21x2_ASAP7_75t_L g1015 ( .A1(n_873), .A2(n_866), .B(n_936), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1016 ( .A(n_867), .Y(n_1016) );
OAI21xp5_ASAP7_75t_L g1017 ( .A1(n_879), .A2(n_978), .B(n_975), .Y(n_1017) );
OA21x2_ASAP7_75t_L g1018 ( .A1(n_866), .A2(n_954), .B(n_967), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_882), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_961), .B(n_968), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_874), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_872), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_872), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1024 ( .A(n_905), .B(n_915), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_883), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_969), .Y(n_1026) );
AND2x4_ASAP7_75t_L g1027 ( .A(n_929), .B(n_977), .Y(n_1027) );
AOI211xp5_ASAP7_75t_SL g1028 ( .A1(n_944), .A2(n_981), .B(n_973), .C(n_925), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_926), .Y(n_1029) );
AO21x2_ASAP7_75t_L g1030 ( .A1(n_954), .A2(n_967), .B(n_912), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_934), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_960), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_937), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_881), .B(n_893), .Y(n_1034) );
BUFx3_ASAP7_75t_L g1035 ( .A(n_932), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_881), .B(n_888), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_885), .B(n_892), .Y(n_1037) );
AO21x2_ASAP7_75t_L g1038 ( .A1(n_869), .A2(n_865), .B(n_966), .Y(n_1038) );
INVx3_ASAP7_75t_L g1039 ( .A(n_868), .Y(n_1039) );
AO21x2_ASAP7_75t_L g1040 ( .A1(n_952), .A2(n_966), .B(n_898), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_917), .B(n_922), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_906), .A2(n_916), .B1(n_894), .B2(n_963), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_946), .Y(n_1043) );
AO21x2_ASAP7_75t_L g1044 ( .A1(n_952), .A2(n_899), .B(n_928), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_935), .B(n_984), .Y(n_1045) );
INVx4_ASAP7_75t_SL g1046 ( .A(n_984), .Y(n_1046) );
AND2x4_ASAP7_75t_L g1047 ( .A(n_921), .B(n_868), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_984), .B(n_972), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_963), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_923), .B(n_931), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_886), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_918), .B(n_877), .Y(n_1052) );
INVx2_ASAP7_75t_SL g1053 ( .A(n_918), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_877), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_895), .Y(n_1055) );
AND2x4_ASAP7_75t_L g1056 ( .A(n_924), .B(n_877), .Y(n_1056) );
OAI222xp33_ASAP7_75t_L g1057 ( .A1(n_962), .A2(n_876), .B1(n_904), .B2(n_938), .C1(n_618), .C2(n_559), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_875), .B(n_900), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_878), .B(n_897), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_974), .A2(n_523), .B1(n_976), .B2(n_528), .C(n_683), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_891), .A2(n_683), .B1(n_876), .B2(n_974), .Y(n_1061) );
AOI33xp33_ASAP7_75t_L g1062 ( .A1(n_985), .A2(n_528), .A3(n_564), .B1(n_474), .B2(n_976), .B3(n_618), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_933), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g1064 ( .A(n_887), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_933), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_933), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_901), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_908), .B(n_927), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_947), .Y(n_1069) );
AO21x2_ASAP7_75t_L g1070 ( .A1(n_939), .A2(n_940), .B(n_941), .Y(n_1070) );
INVxp67_ASAP7_75t_L g1071 ( .A(n_987), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_989), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1029), .B(n_1031), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1001), .B(n_1004), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1001), .B(n_1004), .Y(n_1075) );
INVx3_ASAP7_75t_L g1076 ( .A(n_1033), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1022), .B(n_1023), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_1067), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1048), .B(n_1018), .Y(n_1079) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_1003), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_997), .A2(n_995), .B1(n_1061), .B2(n_1060), .Y(n_1081) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_1045), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_993), .B(n_1059), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1048), .B(n_1018), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_1045), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1018), .B(n_1054), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_987), .B(n_1011), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_1017), .A2(n_1028), .B1(n_988), .B2(n_1012), .C(n_1000), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_1011), .B(n_1013), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1018), .B(n_1054), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1037), .B(n_1036), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1022), .B(n_1023), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_1050), .A2(n_1041), .B1(n_1034), .B2(n_1069), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1033), .B(n_1063), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_1050), .A2(n_1041), .B1(n_1034), .B2(n_1024), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1065), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1066), .B(n_1030), .Y(n_1097) );
INVxp67_ASAP7_75t_L g1098 ( .A(n_1052), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1030), .B(n_1043), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1100 ( .A(n_1052), .B(n_1056), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1051), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_999), .B(n_1006), .Y(n_1102) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_1003), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_999), .B(n_1006), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1009), .B(n_1020), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1009), .B(n_1020), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_998), .B(n_1002), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_1056), .B(n_1046), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1021), .B(n_1025), .Y(n_1109) );
AOI21xp5_ASAP7_75t_L g1110 ( .A1(n_1038), .A2(n_994), .B(n_990), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1021), .B(n_1025), .Y(n_1111) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_1003), .Y(n_1112) );
AOI222xp33_ASAP7_75t_L g1113 ( .A1(n_1057), .A2(n_1026), .B1(n_1007), .B2(n_1062), .C1(n_1016), .C2(n_1010), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1005), .B(n_992), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_1046), .B(n_1003), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1005), .B(n_1015), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1117 ( .A(n_1100), .B(n_1046), .Y(n_1117) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1076), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1105), .B(n_1106), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1105), .B(n_1027), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1121 ( .A(n_1076), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1079), .B(n_1058), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1106), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1101), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1102), .B(n_1027), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1089), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1102), .B(n_1027), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1079), .B(n_1058), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1084), .B(n_1040), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1087), .B(n_1040), .Y(n_1130) );
NAND2xp5_ASAP7_75t_SL g1131 ( .A(n_1113), .B(n_1068), .Y(n_1131) );
OAI31xp33_ASAP7_75t_L g1132 ( .A1(n_1088), .A2(n_1008), .A3(n_1049), .B(n_1035), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1072), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1084), .B(n_1040), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1087), .B(n_1038), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1072), .Y(n_1136) );
INVx2_ASAP7_75t_SL g1137 ( .A(n_1076), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1089), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_1115), .B(n_1032), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1104), .B(n_1024), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1109), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1084), .B(n_1038), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_1078), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1116), .B(n_1044), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1104), .B(n_1074), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1074), .B(n_1024), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1116), .B(n_1044), .Y(n_1147) );
AND2x4_ASAP7_75t_SL g1148 ( .A(n_1115), .B(n_1014), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1109), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1075), .B(n_1024), .Y(n_1150) );
NAND2x1_ASAP7_75t_L g1151 ( .A(n_1076), .B(n_991), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1111), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1071), .B(n_1044), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1096), .Y(n_1154) );
AND2x4_ASAP7_75t_SL g1155 ( .A(n_1114), .B(n_1014), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1073), .B(n_1094), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_1088), .A2(n_1068), .B1(n_1042), .B2(n_1010), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1094), .B(n_986), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1097), .B(n_1083), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1071), .B(n_986), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1097), .B(n_1070), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1122), .B(n_1097), .Y(n_1162) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1124), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_1119), .B(n_1055), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1122), .B(n_1086), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1128), .B(n_1086), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1167 ( .A(n_1123), .B(n_1055), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1159), .B(n_1082), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1156), .B(n_1075), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1170 ( .A(n_1133), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1159), .B(n_1082), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1128), .B(n_1086), .Y(n_1172) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1136), .Y(n_1173) );
BUFx3_ASAP7_75t_L g1174 ( .A(n_1151), .Y(n_1174) );
INVx1_ASAP7_75t_SL g1175 ( .A(n_1155), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1156), .B(n_1083), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1126), .B(n_1114), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1142), .B(n_1090), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1142), .B(n_1090), .Y(n_1179) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1154), .Y(n_1180) );
AND2x4_ASAP7_75t_L g1181 ( .A(n_1139), .B(n_1108), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1141), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1129), .B(n_1099), .Y(n_1183) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_1131), .A2(n_1113), .B1(n_1081), .B2(n_1095), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1149), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1135), .B(n_1085), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1161), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1129), .B(n_1090), .Y(n_1188) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1138), .B(n_1035), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1157), .A2(n_1093), .B1(n_1098), .B2(n_1091), .Y(n_1190) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_1143), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1152), .Y(n_1192) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1161), .Y(n_1193) );
INVx2_ASAP7_75t_SL g1194 ( .A(n_1173), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1162), .B(n_1134), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1183), .B(n_1130), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1170), .Y(n_1197) );
INVx1_ASAP7_75t_SL g1198 ( .A(n_1175), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1180), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1162), .B(n_1134), .Y(n_1200) );
INVxp67_ASAP7_75t_L g1201 ( .A(n_1173), .Y(n_1201) );
NOR2xp67_ASAP7_75t_SL g1202 ( .A(n_1174), .B(n_1064), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1163), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1168), .Y(n_1204) );
OAI21xp5_ASAP7_75t_L g1205 ( .A1(n_1184), .A2(n_1132), .B(n_1107), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1188), .B(n_1145), .Y(n_1206) );
A2O1A1Ixp33_ASAP7_75t_L g1207 ( .A1(n_1184), .A2(n_1155), .B(n_1148), .C(n_1080), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1208 ( .A(n_1191), .Y(n_1208) );
INVxp67_ASAP7_75t_SL g1209 ( .A(n_1191), .Y(n_1209) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_1190), .A2(n_1112), .B1(n_1103), .B2(n_1080), .Y(n_1210) );
INVx1_ASAP7_75t_SL g1211 ( .A(n_1175), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1168), .Y(n_1212) );
BUFx3_ASAP7_75t_L g1213 ( .A(n_1174), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1188), .B(n_1144), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1178), .B(n_1144), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1178), .B(n_1147), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1183), .B(n_1130), .Y(n_1217) );
OAI21xp5_ASAP7_75t_L g1218 ( .A1(n_1190), .A2(n_1107), .B(n_1053), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1171), .Y(n_1219) );
INVx1_ASAP7_75t_SL g1220 ( .A(n_1171), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1204), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1212), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1219), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1197), .Y(n_1224) );
AOI21xp33_ASAP7_75t_SL g1225 ( .A1(n_1207), .A2(n_1064), .B(n_1164), .Y(n_1225) );
AOI22xp5_ASAP7_75t_L g1226 ( .A1(n_1205), .A2(n_1189), .B1(n_1167), .B2(n_1193), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1220), .B(n_1179), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1196), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1196), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_1218), .A2(n_1140), .B1(n_1150), .B2(n_1146), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1201), .B(n_1176), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1217), .B(n_1179), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1217), .Y(n_1233) );
INVxp33_ASAP7_75t_L g1234 ( .A(n_1202), .Y(n_1234) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_1194), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1214), .B(n_1169), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1209), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1194), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1208), .B(n_1165), .Y(n_1239) );
INVxp67_ASAP7_75t_L g1240 ( .A(n_1198), .Y(n_1240) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1203), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1208), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1228), .Y(n_1243) );
AOI21xp33_ASAP7_75t_L g1244 ( .A1(n_1234), .A2(n_1202), .B(n_1210), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_1225), .A2(n_1207), .B1(n_1211), .B2(n_1206), .Y(n_1245) );
AOI21xp5_ASAP7_75t_L g1246 ( .A1(n_1234), .A2(n_1213), .B(n_1151), .Y(n_1246) );
O2A1O1Ixp33_ASAP7_75t_L g1247 ( .A1(n_1240), .A2(n_1053), .B(n_1213), .C(n_1019), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_1224), .Y(n_1248) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_1226), .A2(n_1019), .B1(n_1091), .B2(n_1118), .C(n_1121), .Y(n_1249) );
AOI21xp5_ASAP7_75t_L g1250 ( .A1(n_1235), .A2(n_1181), .B(n_1127), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1229), .Y(n_1251) );
OAI322xp33_ASAP7_75t_L g1252 ( .A1(n_1231), .A2(n_1186), .A3(n_1216), .B1(n_1215), .B2(n_1195), .C1(n_1200), .C2(n_1177), .Y(n_1252) );
NAND3xp33_ASAP7_75t_SL g1253 ( .A(n_1237), .B(n_996), .C(n_1103), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1233), .B(n_1182), .Y(n_1254) );
XOR2x2_ASAP7_75t_L g1255 ( .A(n_1231), .B(n_1010), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_1235), .A2(n_1166), .B1(n_1165), .B2(n_1172), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_1230), .A2(n_1187), .B1(n_1193), .B2(n_1185), .Y(n_1257) );
OAI21xp5_ASAP7_75t_SL g1258 ( .A1(n_1245), .A2(n_1230), .B(n_1148), .Y(n_1258) );
AOI22x1_ASAP7_75t_SL g1259 ( .A1(n_1255), .A2(n_1242), .B1(n_1238), .B2(n_1223), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1260 ( .A1(n_1252), .A2(n_1222), .B1(n_1221), .B2(n_1239), .C(n_1227), .Y(n_1260) );
OAI21xp5_ASAP7_75t_L g1261 ( .A1(n_1247), .A2(n_1239), .B(n_1232), .Y(n_1261) );
NAND5xp2_ASAP7_75t_L g1262 ( .A(n_1244), .B(n_1112), .C(n_1098), .D(n_1110), .E(n_1158), .Y(n_1262) );
AOI22xp5_ASAP7_75t_L g1263 ( .A1(n_1253), .A2(n_1182), .B1(n_1185), .B2(n_1192), .Y(n_1263) );
NAND3xp33_ASAP7_75t_L g1264 ( .A(n_1246), .B(n_1110), .C(n_1241), .Y(n_1264) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_1250), .A2(n_1241), .B(n_1174), .Y(n_1265) );
AOI211xp5_ASAP7_75t_L g1266 ( .A1(n_1249), .A2(n_1160), .B(n_1186), .C(n_1153), .Y(n_1266) );
AOI211xp5_ASAP7_75t_L g1267 ( .A1(n_1249), .A2(n_1160), .B(n_1153), .C(n_1135), .Y(n_1267) );
O2A1O1Ixp33_ASAP7_75t_L g1268 ( .A1(n_1258), .A2(n_1248), .B(n_1256), .C(n_1243), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1269 ( .A1(n_1260), .A2(n_1257), .B1(n_1251), .B2(n_1254), .C(n_1236), .Y(n_1269) );
NOR2x1_ASAP7_75t_L g1270 ( .A(n_1264), .B(n_1068), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1263), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1272 ( .A(n_1259), .B(n_1192), .C(n_1199), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1261), .Y(n_1273) );
NOR3xp33_ASAP7_75t_L g1274 ( .A(n_1262), .B(n_1008), .C(n_1039), .Y(n_1274) );
NAND3xp33_ASAP7_75t_L g1275 ( .A(n_1273), .B(n_1266), .C(n_1267), .Y(n_1275) );
INVxp67_ASAP7_75t_SL g1276 ( .A(n_1270), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1271), .Y(n_1277) );
OAI221xp5_ASAP7_75t_L g1278 ( .A1(n_1268), .A2(n_1265), .B1(n_1080), .B2(n_1121), .C(n_1137), .Y(n_1278) );
OR2x2_ASAP7_75t_SL g1279 ( .A(n_1272), .B(n_1187), .Y(n_1279) );
AND2x2_ASAP7_75t_SL g1280 ( .A(n_1277), .B(n_1274), .Y(n_1280) );
AOI22xp5_ASAP7_75t_L g1281 ( .A1(n_1276), .A2(n_1269), .B1(n_1147), .B2(n_1181), .Y(n_1281) );
NOR3xp33_ASAP7_75t_SL g1282 ( .A(n_1275), .B(n_1120), .C(n_1125), .Y(n_1282) );
INVx3_ASAP7_75t_L g1283 ( .A(n_1278), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1283), .Y(n_1284) );
INVx2_ASAP7_75t_L g1285 ( .A(n_1280), .Y(n_1285) );
INVx2_ASAP7_75t_SL g1286 ( .A(n_1281), .Y(n_1286) );
OA22x2_ASAP7_75t_L g1287 ( .A1(n_1284), .A2(n_1282), .B1(n_1279), .B2(n_1047), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_1285), .B(n_1181), .Y(n_1288) );
AOI21xp5_ASAP7_75t_L g1289 ( .A1(n_1288), .A2(n_1286), .B(n_1047), .Y(n_1289) );
NOR2xp67_ASAP7_75t_SL g1290 ( .A(n_1287), .B(n_1039), .Y(n_1290) );
OAI21xp5_ASAP7_75t_L g1291 ( .A1(n_1289), .A2(n_1092), .B(n_1077), .Y(n_1291) );
AO21x2_ASAP7_75t_L g1292 ( .A1(n_1291), .A2(n_1290), .B(n_1092), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_1292), .A2(n_1187), .B1(n_1193), .B2(n_1117), .Y(n_1293) );
endmodule