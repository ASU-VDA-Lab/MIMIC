module fake_jpeg_3624_n_432 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_49),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_46),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_48),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_51),
.B(n_57),
.Y(n_132)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_67),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx2_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_78),
.Y(n_112)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_70),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_71),
.B(n_75),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_38),
.B1(n_32),
.B2(n_28),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_74),
.B(n_77),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_1),
.Y(n_83)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_17),
.B(n_1),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_31),
.C(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_92),
.B(n_4),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_39),
.B1(n_16),
.B2(n_44),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_93),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_39),
.B1(n_24),
.B2(n_42),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_115),
.B1(n_118),
.B2(n_76),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_16),
.B1(n_18),
.B2(n_33),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_74),
.A2(n_16),
.B1(n_33),
.B2(n_40),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_45),
.A2(n_31),
.B1(n_40),
.B2(n_26),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_42),
.B1(n_38),
.B2(n_24),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_49),
.A2(n_32),
.B1(n_28),
.B2(n_26),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_119),
.A2(n_121),
.B1(n_104),
.B2(n_143),
.Y(n_180)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_55),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_4),
.B(n_5),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_72),
.B(n_71),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_4),
.C(n_5),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_4),
.Y(n_164)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_48),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_149),
.A2(n_151),
.B(n_165),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_150),
.B(n_157),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_62),
.B(n_50),
.C(n_64),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_68),
.B1(n_66),
.B2(n_61),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_153),
.A2(n_183),
.B1(n_186),
.B2(n_177),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_84),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_85),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_161),
.B(n_168),
.Y(n_215)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_46),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_167),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_175),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_82),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_93),
.A2(n_52),
.B(n_64),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_166),
.A2(n_193),
.B(n_170),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_111),
.B(n_80),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_47),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

OR2x4_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_73),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_176),
.A2(n_179),
.B(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_185),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_169),
.B1(n_177),
.B2(n_159),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_98),
.A2(n_54),
.B1(n_73),
.B2(n_65),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_197),
.B1(n_126),
.B2(n_140),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_128),
.A2(n_65),
.B1(n_79),
.B2(n_8),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_189),
.B1(n_196),
.B2(n_131),
.Y(n_212)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_195),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

NAND2x1_ASAP7_75t_SL g204 ( 
.A(n_188),
.B(n_107),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_7),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_102),
.B(n_8),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_155),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_96),
.B(n_9),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_107),
.C(n_100),
.Y(n_203)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_146),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_119),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_121),
.B1(n_140),
.B2(n_109),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_206),
.B1(n_213),
.B2(n_217),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_138),
.B1(n_103),
.B2(n_106),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_201),
.B1(n_209),
.B2(n_222),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_190),
.B1(n_192),
.B2(n_197),
.Y(n_201)
);

AOI221xp5_ASAP7_75t_L g260 ( 
.A1(n_203),
.A2(n_225),
.B1(n_205),
.B2(n_224),
.C(n_214),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_204),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_127),
.B1(n_113),
.B2(n_108),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_152),
.A2(n_126),
.B1(n_131),
.B2(n_165),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_168),
.B1(n_193),
.B2(n_194),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_151),
.A2(n_148),
.B1(n_156),
.B2(n_160),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_157),
.A2(n_185),
.B1(n_164),
.B2(n_150),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_225),
.B1(n_237),
.B2(n_232),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_174),
.B1(n_158),
.B2(n_194),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_226),
.A2(n_227),
.B(n_233),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_221),
.C(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_187),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_178),
.B1(n_184),
.B2(n_173),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_159),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_239),
.A2(n_173),
.B1(n_172),
.B2(n_162),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_242),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_172),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_244),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_188),
.B(n_226),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_273),
.B(n_262),
.Y(n_298)
);

NOR2x1p5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_249),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_188),
.B1(n_199),
.B2(n_213),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_247),
.A2(n_253),
.B(n_267),
.Y(n_295)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_236),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_251),
.A2(n_259),
.B1(n_265),
.B2(n_275),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_201),
.B(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_215),
.B1(n_221),
.B2(n_200),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_251),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_263),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_204),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_268),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_203),
.B1(n_206),
.B2(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_218),
.C(n_229),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_269),
.C(n_264),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_220),
.A2(n_216),
.B(n_208),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_229),
.B(n_211),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_204),
.C(n_220),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_220),
.A2(n_212),
.B1(n_211),
.B2(n_232),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_198),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_219),
.A2(n_234),
.B1(n_198),
.B2(n_207),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_234),
.B(n_273),
.C(n_245),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_257),
.B(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_297),
.C(n_303),
.Y(n_311)
);

O2A1O1Ixp33_ASAP7_75t_SL g285 ( 
.A1(n_273),
.A2(n_246),
.B(n_267),
.C(n_271),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_285),
.A2(n_298),
.B(n_302),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_261),
.B(n_244),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_259),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_287),
.B(n_290),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_255),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_287),
.C(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_242),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_256),
.A2(n_246),
.B(n_269),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_301),
.A2(n_295),
.B(n_298),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_243),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_243),
.B1(n_246),
.B2(n_240),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_262),
.B1(n_270),
.B2(n_241),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_272),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_306),
.Y(n_324)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_314),
.B1(n_313),
.B2(n_328),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_248),
.B1(n_274),
.B2(n_275),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_303),
.B1(n_305),
.B2(n_297),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_315),
.A2(n_316),
.B1(n_323),
.B2(n_311),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_282),
.A2(n_301),
.B1(n_291),
.B2(n_284),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_311),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_318),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_278),
.B(n_307),
.Y(n_320)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_284),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_325),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_304),
.A2(n_290),
.B1(n_292),
.B2(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_304),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_326),
.A2(n_330),
.B(n_310),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_280),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_329),
.C(n_331),
.Y(n_341)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_328),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_279),
.B(n_288),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_300),
.C(n_299),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_277),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_334),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_277),
.C(n_302),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_327),
.Y(n_348)
);

NAND2xp67_ASAP7_75t_SL g334 ( 
.A(n_283),
.B(n_298),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_315),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_345),
.B1(n_350),
.B2(n_353),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_349),
.B(n_352),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_344),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_321),
.B(n_317),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_348),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_340),
.C(n_341),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_326),
.A2(n_310),
.B1(n_322),
.B2(n_324),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_351),
.B1(n_344),
.B2(n_356),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_316),
.B(n_319),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_320),
.A2(n_329),
.B1(n_309),
.B2(n_334),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_333),
.A2(n_331),
.B(n_308),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_309),
.A2(n_314),
.B1(n_313),
.B2(n_312),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_354),
.B(n_357),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_317),
.Y(n_355)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_321),
.B(n_230),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_362),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_339),
.Y(n_363)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_339),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_365),
.B(n_373),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_341),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_372),
.Y(n_385)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_371),
.Y(n_383)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_353),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_369),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_355),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_377),
.C(n_367),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_351),
.C(n_346),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_345),
.B1(n_346),
.B2(n_343),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_378),
.A2(n_391),
.B1(n_364),
.B2(n_368),
.Y(n_397)
);

NOR2x1_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_349),
.Y(n_379)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_384),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_360),
.B(n_336),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

BUFx12_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_388),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_359),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_368),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_381),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_369),
.B1(n_363),
.B2(n_376),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_371),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_382),
.A2(n_392),
.B1(n_381),
.B2(n_393),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_397),
.B1(n_383),
.B2(n_386),
.Y(n_410)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_372),
.C(n_375),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_398),
.B(n_405),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_360),
.Y(n_403)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_379),
.A2(n_391),
.B(n_382),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_385),
.C(n_390),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_407),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_385),
.C(n_384),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_410),
.A2(n_408),
.B1(n_400),
.B2(n_395),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_402),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_404),
.B(n_405),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_396),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_412),
.A2(n_401),
.B1(n_400),
.B2(n_394),
.Y(n_415)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_415),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g421 ( 
.A1(n_416),
.A2(n_409),
.B(n_410),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_420),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_403),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_414),
.C(n_411),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_421),
.Y(n_425)
);

BUFx24_ASAP7_75t_SL g426 ( 
.A(n_424),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_425),
.A2(n_419),
.B(n_423),
.Y(n_427)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_427),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_415),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_429),
.Y(n_430)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_428),
.C(n_422),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_418),
.Y(n_432)
);


endmodule