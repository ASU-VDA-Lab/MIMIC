module fake_jpeg_12531_n_646 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_646);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_646;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_4),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_62),
.B(n_67),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_64),
.Y(n_183)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_68),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_41),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_71),
.B(n_85),
.Y(n_132)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_79),
.Y(n_191)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_80),
.Y(n_150)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_81),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_82),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_83),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_2),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_87),
.Y(n_206)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_88),
.Y(n_210)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_108),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_2),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_102),
.B(n_106),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_2),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_25),
.B(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_116),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_25),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_115),
.B(n_126),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_34),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_22),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_29),
.B(n_4),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_22),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_22),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_133),
.B(n_172),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_135),
.B(n_157),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_143),
.B(n_197),
.Y(n_240)
);

BUFx16f_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_69),
.A2(n_23),
.B1(n_56),
.B2(n_26),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_149),
.A2(n_27),
.B1(n_59),
.B2(n_55),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_60),
.A2(n_128),
.B1(n_105),
.B2(n_88),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_151),
.A2(n_189),
.B1(n_201),
.B2(n_37),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_56),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_152),
.A2(n_59),
.B(n_55),
.Y(n_250)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx11_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_72),
.B(n_40),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_160),
.B(n_168),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_73),
.B(n_44),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_86),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_171),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_92),
.B(n_49),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_75),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_181),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_99),
.B(n_44),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_176),
.B(n_178),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_29),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_77),
.B(n_56),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_207),
.C(n_27),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_79),
.B(n_51),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx16f_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_63),
.A2(n_45),
.B1(n_23),
.B2(n_52),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_64),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_196),
.B(n_36),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_66),
.B(n_49),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_74),
.A2(n_45),
.B1(n_52),
.B2(n_40),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_76),
.B(n_31),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_55),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_78),
.B(n_23),
.C(n_47),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_220),
.Y(n_335)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_222),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g223 ( 
.A(n_139),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_223),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_129),
.B1(n_112),
.B2(n_103),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_225),
.A2(n_233),
.B1(n_243),
.B2(n_255),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_226),
.Y(n_347)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_134),
.B(n_45),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_230),
.B(n_37),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_231),
.B(n_250),
.Y(n_309)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_232),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_132),
.B(n_51),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_235),
.A2(n_244),
.B(n_286),
.Y(n_346)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_236),
.Y(n_339)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_100),
.B1(n_87),
.B2(n_84),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_31),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_245),
.B(n_263),
.Y(n_298)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_247),
.Y(n_345)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

INVx8_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_254),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_179),
.A2(n_59),
.B1(n_36),
.B2(n_30),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_256),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_167),
.Y(n_259)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_261),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_148),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_262),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_138),
.B(n_36),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_265),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_272),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_268),
.B(n_269),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_30),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g270 ( 
.A(n_133),
.B(n_30),
.C(n_27),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_285),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_170),
.A2(n_37),
.B1(n_5),
.B2(n_6),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_271),
.A2(n_185),
.B1(n_204),
.B2(n_147),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_131),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_159),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_277),
.Y(n_320)
);

CKINVDCx12_ASAP7_75t_R g275 ( 
.A(n_161),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_275),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_164),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_278),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_216),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_136),
.B(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_281),
.Y(n_330)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_155),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_166),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_282),
.B(n_284),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_181),
.A2(n_37),
.B1(n_6),
.B2(n_8),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_244),
.B1(n_235),
.B2(n_267),
.Y(n_332)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_175),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_141),
.B(n_4),
.Y(n_286)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_193),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_291),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_290),
.Y(n_306)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_188),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_193),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_154),
.B(n_158),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_204),
.Y(n_314)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_208),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_294),
.Y(n_340)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_137),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_187),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_297),
.B(n_319),
.C(n_194),
.Y(n_393)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_243),
.A2(n_151),
.B(n_171),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_299),
.A2(n_322),
.B1(n_333),
.B2(n_253),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_225),
.A2(n_191),
.B1(n_150),
.B2(n_146),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_301),
.A2(n_307),
.B1(n_277),
.B2(n_287),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_159),
.B(n_185),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_303),
.A2(n_316),
.B(n_334),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_258),
.A2(n_191),
.B1(n_150),
.B2(n_146),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_308),
.A2(n_249),
.B1(n_206),
.B2(n_228),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_343),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_242),
.B(n_240),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_162),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_325),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_242),
.A2(n_218),
.B1(n_216),
.B2(n_162),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_147),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_210),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_326),
.B(n_344),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_271),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_218),
.B1(n_211),
.B2(n_198),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_294),
.A2(n_195),
.B1(n_210),
.B2(n_202),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_233),
.A2(n_142),
.B(n_153),
.C(n_165),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_224),
.B(n_199),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_297),
.B(n_229),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_357),
.B(n_358),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_259),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_359),
.A2(n_392),
.B1(n_398),
.B2(n_299),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_366),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_325),
.B(n_284),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_361),
.B(n_364),
.Y(n_433)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_247),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_365),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_329),
.B(n_255),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_234),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_332),
.B(n_226),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_285),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_368),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_276),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_313),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_383),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_326),
.A2(n_252),
.B(n_221),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_371),
.A2(n_376),
.B(n_390),
.Y(n_430)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_252),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_377),
.Y(n_409)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_302),
.A2(n_246),
.B(n_238),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_330),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_291),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_379),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_274),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_380),
.Y(n_406)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_303),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_273),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_386),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_309),
.B(n_199),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_387),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_319),
.B(n_241),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_273),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_314),
.B(n_260),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_302),
.B(n_142),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_391),
.A2(n_396),
.B1(n_301),
.B2(n_312),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_394),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_306),
.B(n_194),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_299),
.A2(n_211),
.B1(n_198),
.B2(n_206),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_265),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_399),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_349),
.A2(n_186),
.B1(n_219),
.B2(n_9),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_300),
.B(n_6),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_346),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_401),
.B(n_403),
.C(n_405),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_378),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_426),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_310),
.C(n_348),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_341),
.C(n_342),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_410),
.A2(n_396),
.B1(n_365),
.B2(n_366),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_414),
.A2(n_424),
.B1(n_418),
.B2(n_427),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_383),
.A2(n_312),
.B1(n_307),
.B2(n_299),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_418),
.A2(n_424),
.B1(n_397),
.B2(n_398),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_328),
.C(n_311),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_431),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_391),
.A2(n_299),
.B1(n_300),
.B2(n_343),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_381),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g426 ( 
.A(n_377),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_295),
.C(n_352),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_295),
.C(n_352),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_336),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_354),
.A2(n_334),
.B1(n_340),
.B2(n_306),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_434),
.A2(n_374),
.B1(n_365),
.B2(n_385),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_354),
.A2(n_340),
.B(n_320),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_437),
.A2(n_365),
.B(n_360),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_381),
.A2(n_371),
.B(n_364),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_438),
.A2(n_392),
.B(n_359),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_439),
.A2(n_447),
.B1(n_404),
.B2(n_405),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_407),
.B(n_370),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_441),
.B(n_453),
.Y(n_477)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

INVx13_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_443),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_374),
.Y(n_444)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_445),
.A2(n_456),
.B1(n_461),
.B2(n_465),
.Y(n_503)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_446),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_415),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_460),
.Y(n_483)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_450),
.Y(n_507)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_458),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_358),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_376),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_455),
.B(n_336),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_457),
.A2(n_473),
.B(n_404),
.Y(n_492)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_407),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_462),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_425),
.B(n_379),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_434),
.A2(n_382),
.B1(n_373),
.B2(n_390),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_399),
.Y(n_462)
);

AO22x1_ASAP7_75t_L g463 ( 
.A1(n_437),
.A2(n_420),
.B1(n_373),
.B2(n_430),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_464),
.Y(n_485)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_429),
.A2(n_394),
.B1(n_395),
.B2(n_388),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_367),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_468),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_368),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_469),
.Y(n_487)
);

OAI32xp33_ASAP7_75t_L g468 ( 
.A1(n_409),
.A2(n_361),
.A3(n_390),
.B1(n_389),
.B2(n_360),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_384),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_412),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_335),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_435),
.B(n_369),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_417),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_408),
.C(n_401),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_475),
.B(n_481),
.C(n_482),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_408),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_478),
.B(n_470),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_445),
.A2(n_409),
.B1(n_430),
.B2(n_400),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_479),
.A2(n_488),
.B1(n_463),
.B2(n_444),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_416),
.C(n_431),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_438),
.B1(n_414),
.B2(n_416),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_489),
.A2(n_496),
.B1(n_505),
.B2(n_501),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_492),
.A2(n_498),
.B(n_501),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g522 ( 
.A(n_493),
.Y(n_522)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_335),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_495),
.B(n_504),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_450),
.A2(n_413),
.B1(n_411),
.B2(n_375),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_417),
.C(n_423),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_497),
.B(n_449),
.C(n_451),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_455),
.A2(n_411),
.B(n_362),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_459),
.B(n_380),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_457),
.A2(n_372),
.B(n_337),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_502),
.A2(n_446),
.B(n_442),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_339),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_439),
.A2(n_447),
.B1(n_455),
.B2(n_448),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_304),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_506),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_475),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_509),
.B(n_524),
.Y(n_550)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_488),
.A2(n_463),
.B1(n_468),
.B2(n_444),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_513),
.A2(n_505),
.B1(n_489),
.B2(n_507),
.Y(n_543)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_474),
.Y(n_514)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_514),
.Y(n_541)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_516),
.A2(n_525),
.B1(n_491),
.B2(n_477),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_480),
.Y(n_518)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_518),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_466),
.Y(n_520)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_520),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_521),
.A2(n_490),
.B1(n_486),
.B2(n_480),
.Y(n_559)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_484),
.Y(n_523)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_481),
.B(n_454),
.Y(n_524)
);

AOI22x1_ASAP7_75t_L g525 ( 
.A1(n_491),
.A2(n_462),
.B1(n_441),
.B2(n_456),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_472),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_527),
.B(n_532),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_528),
.A2(n_537),
.B(n_506),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_530),
.C(n_535),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_493),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_499),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_476),
.B(n_458),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_533),
.Y(n_556)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_476),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_536),
.Y(n_560)
);

MAJx2_ASAP7_75t_L g535 ( 
.A(n_497),
.B(n_356),
.C(n_443),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_500),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_443),
.B(n_317),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_538),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_482),
.C(n_485),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_542),
.B(n_547),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_552),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_519),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_562),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_522),
.A2(n_503),
.B1(n_479),
.B2(n_507),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_545),
.A2(n_558),
.B1(n_559),
.B2(n_508),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_485),
.C(n_502),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_518),
.B(n_490),
.Y(n_548)
);

AOI221xp5_ASAP7_75t_L g563 ( 
.A1(n_548),
.A2(n_514),
.B1(n_515),
.B2(n_511),
.C(n_486),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_502),
.C(n_498),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_553),
.B(n_561),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_554),
.B(n_517),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_SL g558 ( 
.A(n_520),
.B(n_508),
.C(n_506),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_510),
.B(n_516),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_533),
.Y(n_562)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_563),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_539),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_564),
.B(n_580),
.Y(n_593)
);

XOR2x2_ASAP7_75t_L g588 ( 
.A(n_565),
.B(n_571),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_SL g567 ( 
.A(n_553),
.B(n_526),
.C(n_509),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_567),
.B(n_578),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_529),
.C(n_535),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_570),
.C(n_576),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_550),
.B(n_537),
.C(n_517),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_SL g572 ( 
.A(n_540),
.B(n_525),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_573),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_513),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_547),
.A2(n_525),
.B(n_528),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_575),
.A2(n_570),
.B(n_579),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_542),
.B(n_490),
.C(n_500),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_315),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_543),
.B(n_337),
.C(n_317),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_581),
.C(n_548),
.Y(n_587)
);

FAx1_ASAP7_75t_SL g580 ( 
.A(n_538),
.B(n_356),
.CI(n_315),
.CON(n_580),
.SN(n_580)
);

XNOR2x1_ASAP7_75t_SL g581 ( 
.A(n_545),
.B(n_347),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_539),
.B(n_350),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_583),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_556),
.Y(n_586)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_586),
.Y(n_603)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_566),
.A2(n_559),
.B1(n_541),
.B2(n_549),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_589),
.A2(n_597),
.B1(n_599),
.B2(n_339),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_576),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_592),
.B(n_594),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_582),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_554),
.C(n_541),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_595),
.B(n_596),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_549),
.C(n_546),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_577),
.A2(n_555),
.B1(n_560),
.B2(n_557),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_577),
.A2(n_555),
.B1(n_558),
.B2(n_557),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_600),
.B(n_353),
.C(n_327),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_580),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_350),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_598),
.B(n_574),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_607),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_585),
.B(n_573),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_584),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_574),
.C(n_568),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_580),
.C(n_581),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_608),
.B(n_610),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_591),
.B(n_546),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_345),
.C(n_353),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_611),
.B(n_586),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_589),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_613),
.B(n_602),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_614),
.A2(n_593),
.B(n_599),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_595),
.B(n_327),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_615),
.B(n_596),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_616),
.Y(n_627)
);

OAI21x1_ASAP7_75t_SL g630 ( 
.A1(n_618),
.A2(n_588),
.B(n_608),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_619),
.B(n_620),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_606),
.A2(n_593),
.B1(n_587),
.B2(n_590),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_621),
.A2(n_626),
.B(n_605),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_623),
.B(n_10),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_584),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_624),
.B(n_625),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_603),
.B(n_588),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_628),
.A2(n_630),
.B(n_633),
.Y(n_636)
);

AOI322xp5_ASAP7_75t_L g631 ( 
.A1(n_622),
.A2(n_614),
.A3(n_345),
.B1(n_219),
.B2(n_347),
.C1(n_12),
.C2(n_13),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_631),
.B(n_634),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_617),
.A2(n_8),
.B(n_9),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_629),
.A2(n_618),
.B(n_623),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_637),
.A2(n_627),
.B(n_11),
.C(n_14),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_624),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_638),
.A2(n_639),
.B(n_10),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_627),
.A2(n_10),
.B(n_11),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_640),
.A2(n_641),
.B(n_636),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_635),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_10),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_15),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_15),
.B(n_621),
.Y(n_646)
);


endmodule