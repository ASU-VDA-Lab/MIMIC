module fake_jpeg_5730_n_113 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_10),
.B(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_13),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_22),
.C(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_22),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_22),
.C(n_12),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_22),
.B(n_19),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_12),
.C(n_16),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_25),
.B1(n_24),
.B2(n_14),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_41),
.B1(n_40),
.B2(n_17),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_11),
.B2(n_14),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_35),
.B1(n_11),
.B2(n_37),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_15),
.B1(n_28),
.B2(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_50),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_47),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_51),
.B1(n_46),
.B2(n_47),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.C(n_61),
.Y(n_63)
);

NOR2xp67_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_62),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_29),
.C(n_21),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_71),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_67),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_51),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_17),
.B(n_16),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_15),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_60),
.B1(n_58),
.B2(n_28),
.Y(n_76)
);

XOR2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_61),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_21),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_19),
.C(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_2),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_19),
.B(n_15),
.C(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_74),
.B1(n_78),
.B2(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_63),
.B(n_72),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_87),
.B1(n_81),
.B2(n_6),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_75),
.C(n_83),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_3),
.CI(n_5),
.CON(n_88),
.SN(n_88)
);

AOI21x1_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_90),
.B(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_97),
.C(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_6),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_3),
.C(n_6),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_97),
.C(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_91),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_102),
.B(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_8),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_7),
.B(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_8),
.C(n_109),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_111),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_110),
.Y(n_113)
);


endmodule