module fake_jpeg_25923_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_44),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_35),
.B1(n_18),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_64),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_35),
.B1(n_18),
.B2(n_19),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_56),
.Y(n_86)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_25),
.B(n_22),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_33),
.B(n_1),
.Y(n_91)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_22),
.B(n_21),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_67),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_28),
.Y(n_73)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_76),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_92),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_16),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_14),
.Y(n_118)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_40),
.B1(n_41),
.B2(n_38),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_87),
.B(n_33),
.C(n_93),
.Y(n_107)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_82),
.B(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_26),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_37),
.B1(n_26),
.B2(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_33),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_104),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx10_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_53),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_113),
.B(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_100),
.B(n_114),
.C(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_65),
.C(n_67),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_51),
.C(n_54),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_52),
.B1(n_56),
.B2(n_66),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_75),
.B1(n_76),
.B2(n_72),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_57),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_118),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_79),
.B(n_24),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_83),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_129),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_74),
.B(n_92),
.C(n_93),
.D(n_25),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_130),
.B(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_75),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_132),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_50),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_138),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_50),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_141),
.C(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_115),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_113),
.B(n_107),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_157),
.B(n_159),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_155),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_160),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_96),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_163),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_143),
.B(n_126),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_34),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_107),
.B1(n_105),
.B2(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_83),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_139),
.B1(n_141),
.B2(n_134),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_51),
.C(n_54),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_71),
.B1(n_90),
.B2(n_89),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_SL g171 ( 
.A(n_152),
.B(n_127),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_186),
.B1(n_170),
.B2(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_127),
.B1(n_71),
.B2(n_89),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_181),
.B1(n_185),
.B2(n_190),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_20),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_177),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_51),
.B1(n_97),
.B2(n_50),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_34),
.B1(n_32),
.B2(n_25),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_158),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_16),
.C(n_15),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_162),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_167),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_166),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_163),
.C(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_179),
.C(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_202),
.B(n_210),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_164),
.B1(n_146),
.B2(n_147),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_175),
.B1(n_185),
.B2(n_182),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_178),
.B(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_211),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_168),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_207),
.C(n_173),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_169),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_220),
.B(n_208),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_222),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_173),
.C(n_157),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_226),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_147),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_224),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_0),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_208),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_202),
.B1(n_195),
.B2(n_194),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_198),
.Y(n_239)
);

OAI221xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_240),
.B1(n_189),
.B2(n_5),
.C(n_6),
.Y(n_247)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_229),
.B1(n_228),
.B2(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_218),
.C(n_214),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_216),
.B(n_224),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_247),
.B(n_3),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_207),
.B1(n_196),
.B2(n_30),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_254),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_235),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_256),
.B(n_242),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_232),
.C(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_255),
.C(n_5),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_232),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_254),
.B(n_8),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_248),
.B(n_6),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_7),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_248),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_7),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_266),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.C1(n_261),
.C2(n_74),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_10),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_267),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_12),
.Y(n_271)
);


endmodule