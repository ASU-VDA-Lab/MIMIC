module fake_jpeg_27266_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx10_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_4),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_3),
.B(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_1),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_13),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_6),
.B1(n_13),
.B2(n_11),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_10),
.B1(n_14),
.B2(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_12),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_24),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_14),
.C(n_10),
.Y(n_24)
);

OAI322xp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_7),
.A3(n_9),
.B1(n_16),
.B2(n_18),
.C1(n_21),
.C2(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_21),
.B1(n_10),
.B2(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_32),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_29),
.B(n_28),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_7),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_7),
.B(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule