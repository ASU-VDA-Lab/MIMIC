module fake_jpeg_25999_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_20),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_29),
.Y(n_50)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AO22x1_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_54),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_31),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_25),
.B1(n_22),
.B2(n_27),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_33),
.B1(n_39),
.B2(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_16),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_63),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_23),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_70),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_33),
.B1(n_41),
.B2(n_20),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_62),
.B1(n_61),
.B2(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_41),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_38),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_83),
.B(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_90),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_92),
.B1(n_99),
.B2(n_100),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_61),
.B1(n_24),
.B2(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_96),
.Y(n_118)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_103),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_40),
.B(n_56),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_37),
.B1(n_57),
.B2(n_24),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_40),
.A3(n_18),
.B1(n_60),
.B2(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_40),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_56),
.C(n_70),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_80),
.B(n_76),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_116),
.B(n_120),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_75),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_65),
.B1(n_72),
.B2(n_66),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_117),
.B1(n_100),
.B2(n_68),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_91),
.B(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_65),
.B1(n_72),
.B2(n_66),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_80),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_60),
.B(n_49),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_89),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_95),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_125),
.C(n_127),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_103),
.C(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_88),
.C(n_102),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_131),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_88),
.C(n_99),
.Y(n_131)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_140),
.B1(n_114),
.B2(n_138),
.C(n_120),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_85),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_113),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_74),
.C(n_56),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_137),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_74),
.C(n_56),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_148),
.B(n_150),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_111),
.C(n_112),
.Y(n_146)
);

OA21x2_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_10),
.B(n_9),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_121),
.B1(n_123),
.B2(n_109),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_94),
.B1(n_57),
.B2(n_18),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

OAI31xp33_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_120),
.A3(n_123),
.B(n_113),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_57),
.B(n_60),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_0),
.B(n_1),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_124),
.C(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_160),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_110),
.B1(n_135),
.B2(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_151),
.B(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_15),
.C(n_12),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_12),
.C(n_11),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_152),
.B(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_163),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_161),
.B1(n_159),
.B2(n_173),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_142),
.B1(n_165),
.B2(n_145),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.C(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_158),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_166),
.B(n_180),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_177),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_180),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_179),
.B(n_1),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_160),
.C(n_3),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_183),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_176),
.B(n_6),
.C(n_7),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_189),
.C(n_188),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_5),
.C(n_7),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_185),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_193),
.C(n_5),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_190),
.Y(n_193)
);


endmodule