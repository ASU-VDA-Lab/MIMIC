module fake_jpeg_11816_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_7),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_58),
.B(n_13),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_64),
.Y(n_112)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_29),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_78),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_97),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_96),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_38),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_104),
.B(n_128),
.Y(n_169)
);

INVx6_ASAP7_75t_SL g127 ( 
.A(n_64),
.Y(n_127)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_58),
.B(n_25),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_155),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_35),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_139),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_59),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_142),
.B(n_150),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_36),
.B1(n_47),
.B2(n_46),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_47),
.B1(n_36),
.B2(n_56),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_35),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_24),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_86),
.B(n_42),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_156),
.B(n_158),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_71),
.B(n_35),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_103),
.A2(n_46),
.B1(n_41),
.B2(n_25),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_83),
.B1(n_81),
.B2(n_79),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_52),
.B(n_33),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_26),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_164),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_152),
.Y(n_165)
);

BUFx2_ASAP7_75t_SL g224 ( 
.A(n_165),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_99),
.B1(n_97),
.B2(n_88),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_174),
.B1(n_208),
.B2(n_218),
.Y(n_233)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_77),
.B1(n_76),
.B2(n_75),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_176),
.A2(n_44),
.B1(n_23),
.B2(n_22),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_178),
.A2(n_187),
.B1(n_189),
.B2(n_193),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

CKINVDCx12_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_32),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_198),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_36),
.B1(n_46),
.B2(n_41),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_119),
.A2(n_36),
.B1(n_46),
.B2(n_32),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_143),
.A2(n_42),
.B1(n_25),
.B2(n_32),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_119),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_200),
.Y(n_231)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_195),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g271 ( 
.A(n_196),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_131),
.Y(n_198)
);

NAND2x1_ASAP7_75t_SL g199 ( 
.A(n_109),
.B(n_22),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_199),
.B(n_112),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_126),
.B(n_28),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_124),
.B(n_28),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_201),
.B(n_209),
.Y(n_253)
);

OR2x2_ASAP7_75t_SL g202 ( 
.A(n_152),
.B(n_11),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g257 ( 
.A(n_202),
.B(n_22),
.C(n_44),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_141),
.B(n_61),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_207),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

BUFx24_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_145),
.A2(n_60),
.B1(n_54),
.B2(n_53),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_135),
.B(n_30),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_117),
.B(n_30),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_105),
.B(n_33),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_105),
.B(n_23),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_123),
.A2(n_48),
.B1(n_34),
.B2(n_24),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g221 ( 
.A(n_137),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_116),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_107),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_229),
.B(n_267),
.Y(n_284)
);

AO22x2_ASAP7_75t_L g232 ( 
.A1(n_178),
.A2(n_115),
.B1(n_148),
.B2(n_116),
.Y(n_232)
);

AO22x1_ASAP7_75t_SL g292 ( 
.A1(n_232),
.A2(n_167),
.B1(n_165),
.B2(n_179),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_171),
.A2(n_157),
.B1(n_154),
.B2(n_140),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_245),
.B1(n_138),
.B2(n_195),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_220),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_113),
.C(n_112),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_264),
.C(n_207),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_115),
.B1(n_132),
.B2(n_154),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_140),
.B1(n_107),
.B2(n_148),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_249),
.B(n_44),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_254),
.B(n_31),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_207),
.B(n_48),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_177),
.B(n_147),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_261),
.B(n_266),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_204),
.B(n_121),
.C(n_132),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_147),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_202),
.B(n_222),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_269),
.A2(n_193),
.B1(n_189),
.B2(n_187),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_274),
.B(n_31),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_275),
.A2(n_283),
.B1(n_297),
.B2(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_276),
.B(n_281),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_277),
.A2(n_288),
.B1(n_302),
.B2(n_315),
.Y(n_324)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_278),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_SL g330 ( 
.A(n_279),
.B(n_290),
.Y(n_330)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_223),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_280),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_224),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_234),
.B(n_169),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_286),
.B(n_291),
.Y(n_336)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_233),
.A2(n_185),
.B1(n_184),
.B2(n_173),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_231),
.B(n_34),
.Y(n_291)
);

OA22x2_ASAP7_75t_L g348 ( 
.A1(n_292),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_203),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_293),
.B(n_298),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_138),
.B1(n_168),
.B2(n_205),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_167),
.A3(n_175),
.B1(n_180),
.B2(n_181),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_299),
.B(n_303),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_229),
.B(n_210),
.C(n_206),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_305),
.C(n_249),
.Y(n_326)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_242),
.A2(n_196),
.B1(n_188),
.B2(n_182),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_226),
.B(n_166),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_164),
.C(n_137),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_306),
.B(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_225),
.B(n_10),
.Y(n_308)
);

INVx13_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_309),
.A2(n_310),
.B1(n_312),
.B2(n_318),
.Y(n_327)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_311),
.A2(n_302),
.B(n_310),
.Y(n_355)
);

INVx13_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_239),
.A2(n_246),
.B1(n_232),
.B2(n_242),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_245),
.A2(n_23),
.B1(n_57),
.B2(n_137),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_0),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_317),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_244),
.B(n_240),
.Y(n_333)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_320),
.Y(n_345)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_232),
.B1(n_249),
.B2(n_257),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_325),
.A2(n_334),
.B1(n_339),
.B2(n_340),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_326),
.B(n_354),
.C(n_312),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_232),
.B(n_249),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_331),
.A2(n_332),
.B(n_355),
.Y(n_397)
);

AO22x1_ASAP7_75t_L g332 ( 
.A1(n_311),
.A2(n_244),
.B1(n_256),
.B2(n_263),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_284),
.A2(n_270),
.B1(n_248),
.B2(n_250),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_337),
.B(n_282),
.Y(n_390)
);

AO22x1_ASAP7_75t_SL g338 ( 
.A1(n_313),
.A2(n_270),
.B1(n_260),
.B2(n_258),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_347),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_279),
.A2(n_230),
.B1(n_260),
.B2(n_258),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_275),
.A2(n_252),
.B1(n_251),
.B2(n_262),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_284),
.A2(n_262),
.B1(n_251),
.B2(n_259),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_361),
.B1(n_320),
.B2(n_294),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_259),
.B1(n_241),
.B2(n_240),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_346),
.A2(n_351),
.B1(n_356),
.B2(n_306),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_241),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_1),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_274),
.A2(n_285),
.B1(n_305),
.B2(n_316),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_292),
.A2(n_9),
.B1(n_15),
.B2(n_13),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_296),
.A2(n_1),
.B(n_3),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_358),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_292),
.A2(n_1),
.B(n_3),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_277),
.A2(n_15),
.B1(n_12),
.B2(n_10),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_328),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_364),
.Y(n_399)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_291),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_368),
.B(n_384),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_314),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_375),
.C(n_381),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_356),
.Y(n_406)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_344),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_373),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_352),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_319),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_345),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_377),
.B(n_390),
.Y(n_414)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_307),
.Y(n_379)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_330),
.B(n_290),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_382),
.A2(n_396),
.B1(n_324),
.B2(n_355),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_289),
.Y(n_383)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_301),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_358),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_386),
.B(n_391),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_304),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_389),
.C(n_395),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_299),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_329),
.B(n_280),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_335),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_343),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_321),
.A2(n_287),
.B1(n_318),
.B2(n_295),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_397),
.A2(n_331),
.B(n_360),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_400),
.A2(n_379),
.B(n_348),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_321),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_413),
.C(n_424),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_383),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_405),
.B(n_367),
.Y(n_445)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_332),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_387),
.B1(n_364),
.B2(n_370),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_417),
.B(n_404),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_333),
.B(n_327),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_381),
.B(n_348),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_422),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_394),
.A2(n_355),
.B(n_332),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_396),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_340),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_338),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_428),
.C(n_365),
.Y(n_432)
);

OA22x2_ASAP7_75t_L g426 ( 
.A1(n_397),
.A2(n_346),
.B1(n_348),
.B2(n_338),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_349),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_342),
.C(n_362),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_402),
.A2(n_376),
.B1(n_382),
.B2(n_365),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_429),
.A2(n_437),
.B1(n_400),
.B2(n_426),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_446),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_427),
.B(n_357),
.Y(n_433)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_439),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_401),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_448),
.Y(n_455)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_441),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_414),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_445),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_392),
.C(n_385),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_454),
.C(n_424),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_412),
.B(n_374),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_278),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_425),
.Y(n_459)
);

NAND2xp67_ASAP7_75t_SL g449 ( 
.A(n_423),
.B(n_380),
.Y(n_449)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

A2O1A1O1Ixp25_ASAP7_75t_L g450 ( 
.A1(n_411),
.A2(n_342),
.B(n_362),
.C(n_349),
.D(n_309),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g458 ( 
.A(n_450),
.B(n_419),
.CI(n_428),
.CON(n_458),
.SN(n_458)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_399),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_453),
.A2(n_408),
.B1(n_323),
.B2(n_409),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_323),
.C(n_371),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_470),
.C(n_472),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_435),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_457),
.B(n_460),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_469),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_465),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_413),
.C(n_416),
.Y(n_460)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_429),
.A2(n_426),
.B1(n_422),
.B2(n_406),
.Y(n_466)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_466),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_443),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_422),
.C(n_426),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_420),
.C(n_418),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_473),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_432),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_484),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_447),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_464),
.A2(n_452),
.B1(n_437),
.B2(n_430),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_485),
.A2(n_489),
.B1(n_468),
.B2(n_476),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_431),
.C(n_446),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_490),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_439),
.B1(n_430),
.B2(n_438),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_407),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_455),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_492),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_442),
.C(n_438),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_442),
.B(n_449),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_493),
.A2(n_468),
.B1(n_482),
.B2(n_480),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_497),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_471),
.C(n_470),
.Y(n_497)
);

XNOR2x1_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_465),
.Y(n_498)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_498),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_471),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_503),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_505),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_464),
.C(n_467),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_502),
.B(n_504),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_479),
.B(n_466),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_476),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_485),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_481),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_508),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_487),
.B(n_458),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_495),
.Y(n_523)
);

AOI21xp33_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_483),
.B(n_486),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_513),
.A2(n_517),
.B(n_450),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_506),
.A2(n_463),
.B(n_458),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_514),
.A2(n_516),
.B(n_441),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_497),
.A2(n_408),
.B(n_475),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_453),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g520 ( 
.A(n_519),
.B(n_505),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_520),
.A2(n_521),
.B(n_522),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_499),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_524),
.C(n_511),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_503),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_526),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_498),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_529),
.B(n_436),
.Y(n_531)
);

AOI322xp5_ASAP7_75t_L g529 ( 
.A1(n_522),
.A2(n_513),
.A3(n_510),
.B1(n_409),
.B2(n_436),
.C1(n_407),
.C2(n_378),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_532),
.A3(n_530),
.B1(n_31),
.B2(n_9),
.C1(n_6),
.C2(n_3),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_12),
.B(n_10),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_4),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_8),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_536),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_6),
.B1(n_8),
.B2(n_531),
.Y(n_538)
);


endmodule