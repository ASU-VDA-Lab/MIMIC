module fake_netlist_1_1431_n_650 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_650);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_650;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_58), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_36), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_78), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_14), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_75), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_16), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_62), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_69), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_31), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_61), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_66), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_15), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_37), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_25), .Y(n_97) );
BUFx2_ASAP7_75t_SL g98 ( .A(n_42), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_32), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_52), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_53), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_50), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_2), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_34), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_22), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_64), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_10), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_70), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_60), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_21), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_54), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_39), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_27), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_16), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_5), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_4), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
NOR2xp67_ASAP7_75t_L g121 ( .A(n_5), .B(n_74), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_35), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_55), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_4), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_6), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_3), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_94), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_83), .B(n_0), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_111), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_111), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_114), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_117), .B(n_110), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_107), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_89), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_106), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_109), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_79), .Y(n_139) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_108), .B(n_76), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_123), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_114), .B(n_0), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_82), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_86), .B(n_1), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_86), .B(n_1), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_80), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
NAND2xp33_ASAP7_75t_R g153 ( .A(n_88), .B(n_29), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_98), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_93), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_98), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_114), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_95), .B(n_2), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_87), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_115), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_95), .B(n_3), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_119), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_92), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_119), .B(n_6), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_135), .B(n_126), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_135), .B(n_126), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVx8_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_132), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_128), .B(n_101), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_146), .B(n_124), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_132), .A2(n_124), .B1(n_125), .B2(n_104), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_165), .B(n_122), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_128), .A2(n_116), .B1(n_90), .B2(n_120), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_163), .B(n_122), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_132), .B(n_80), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_129), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_146), .B(n_102), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_137), .B(n_139), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_130), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
AND2x6_ASAP7_75t_L g201 ( .A(n_166), .B(n_102), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_131), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_158), .B(n_103), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_137), .B(n_96), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_160), .B(n_103), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_139), .B(n_96), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_167), .B(n_90), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_134), .B(n_91), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_167), .B(n_91), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_166), .B(n_112), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_141), .B(n_99), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_168), .B(n_112), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_149), .B(n_99), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_169), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_151), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_140), .A2(n_105), .B1(n_120), .B2(n_118), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_149), .B(n_118), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_136), .B(n_113), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_152), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_217), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_175), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_195), .B(n_162), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_206), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_201), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_195), .B(n_169), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_209), .Y(n_239) );
NAND3xp33_ASAP7_75t_SL g240 ( .A(n_189), .B(n_138), .C(n_159), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g241 ( .A1(n_224), .A2(n_133), .B1(n_150), .B2(n_147), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_204), .Y(n_243) );
NAND3xp33_ASAP7_75t_SL g244 ( .A(n_176), .B(n_127), .C(n_147), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_197), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_195), .B(n_162), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_205), .B(n_212), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_205), .B(n_157), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_213), .B(n_150), .C(n_153), .Y(n_251) );
INVx3_ASAP7_75t_SL g252 ( .A(n_175), .Y(n_252) );
BUFx8_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_209), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_205), .B(n_140), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_212), .B(n_157), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_171), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_171), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_178), .Y(n_261) );
NOR3xp33_ASAP7_75t_SL g262 ( .A(n_228), .B(n_144), .C(n_156), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_212), .B(n_152), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_214), .B(n_156), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_172), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_172), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_174), .A2(n_151), .B(n_101), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_214), .B(n_140), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_174), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_215), .B(n_169), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_186), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_192), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_184), .Y(n_274) );
INVx4_ASAP7_75t_L g275 ( .A(n_178), .Y(n_275) );
OR2x6_ASAP7_75t_L g276 ( .A(n_186), .B(n_151), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_192), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_170), .B(n_113), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_170), .B(n_100), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_178), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_193), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_184), .Y(n_284) );
NOR3xp33_ASAP7_75t_SL g285 ( .A(n_182), .B(n_100), .C(n_121), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_186), .A2(n_161), .B1(n_131), .B2(n_9), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_215), .B(n_161), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_193), .Y(n_288) );
INVx11_ASAP7_75t_L g289 ( .A(n_201), .Y(n_289) );
NOR3xp33_ASAP7_75t_SL g290 ( .A(n_220), .B(n_7), .C(n_8), .Y(n_290) );
NOR2xp33_ASAP7_75t_R g291 ( .A(n_194), .B(n_38), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_178), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_226), .B(n_161), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_252), .B(n_194), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_259), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_259), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_238), .B(n_201), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_252), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_221), .B(n_219), .Y(n_300) );
BUFx4_ASAP7_75t_SL g301 ( .A(n_243), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_252), .B(n_255), .Y(n_302) );
AOI21x1_ASAP7_75t_L g303 ( .A1(n_260), .A2(n_229), .B(n_219), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_233), .B(n_222), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_234), .A2(n_177), .B(n_190), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_265), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_253), .Y(n_309) );
CKINVDCx8_ASAP7_75t_R g310 ( .A(n_243), .Y(n_310) );
INVx5_ASAP7_75t_L g311 ( .A(n_232), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
INVx5_ASAP7_75t_L g313 ( .A(n_232), .Y(n_313) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_275), .B(n_226), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_233), .B(n_203), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_187), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_255), .A2(n_201), .B1(n_178), .B2(n_184), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_230), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_266), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_238), .B(n_179), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_232), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_230), .Y(n_323) );
AND2x2_ASAP7_75t_SL g324 ( .A(n_275), .B(n_226), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g325 ( .A1(n_253), .A2(n_173), .B1(n_178), .B2(n_179), .Y(n_325) );
AO32x2_ASAP7_75t_L g326 ( .A1(n_286), .A2(n_216), .A3(n_183), .B1(n_223), .B2(n_188), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_241), .A2(n_173), .B1(n_180), .B2(n_199), .C(n_210), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_240), .B(n_216), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_232), .B(n_229), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_238), .B(n_198), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_269), .A2(n_248), .B1(n_250), .B2(n_257), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_247), .A2(n_207), .B(n_211), .C(n_223), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_264), .B(n_223), .Y(n_334) );
NAND2xp33_ASAP7_75t_L g335 ( .A(n_261), .B(n_272), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_273), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_230), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_249), .A2(n_256), .B(n_263), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_273), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_276), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_276), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_271), .B(n_7), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_236), .A2(n_227), .B1(n_181), .B2(n_218), .Y(n_343) );
OAI22xp33_ASAP7_75t_SL g344 ( .A1(n_310), .A2(n_276), .B1(n_244), .B2(n_278), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_299), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_305), .A2(n_268), .B1(n_236), .B2(n_257), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_342), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_334), .Y(n_348) );
OAI222xp33_ASAP7_75t_L g349 ( .A1(n_310), .A2(n_276), .B1(n_272), .B2(n_279), .C1(n_268), .C2(n_292), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_312), .A2(n_233), .B1(n_232), .B2(n_242), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_297), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_299), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_334), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_297), .A2(n_239), .B(n_292), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_330), .B(n_262), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_304), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_302), .B(n_275), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_295), .B(n_261), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_302), .A2(n_242), .B1(n_274), .B2(n_284), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_330), .B(n_251), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_307), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_304), .A2(n_315), .B1(n_327), .B2(n_324), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_315), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_315), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_315), .B(n_292), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_311), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_314), .B(n_280), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_301), .Y(n_371) );
NAND2xp33_ASAP7_75t_R g372 ( .A(n_328), .B(n_291), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_340), .B(n_242), .Y(n_373) );
INVx8_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_316), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_365), .A2(n_328), .B1(n_325), .B2(n_321), .C(n_285), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_360), .A2(n_314), .B1(n_324), .B2(n_341), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_352), .B(n_314), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_363), .A2(n_324), .B1(n_309), .B2(n_298), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_357), .A2(n_309), .B1(n_319), .B2(n_316), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_344), .A2(n_339), .B1(n_336), .B2(n_307), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_347), .A2(n_332), .B(n_338), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_375), .Y(n_383) );
BUFx12f_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_351), .A2(n_333), .B1(n_339), .B2(n_336), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_348), .A2(n_290), .B(n_317), .C(n_331), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_295), .Y(n_387) );
INVx8_ASAP7_75t_L g388 ( .A(n_374), .Y(n_388) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_354), .A2(n_303), .B(n_296), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_360), .A2(n_294), .B1(n_306), .B2(n_300), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_361), .A2(n_303), .B(n_296), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_372), .A2(n_300), .B1(n_320), .B2(n_287), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_360), .A2(n_289), .B1(n_320), .B2(n_300), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_355), .B(n_311), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_371), .A2(n_313), .B1(n_322), .B2(n_311), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_349), .A2(n_329), .B(n_239), .C(n_318), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_368), .B(n_300), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_368), .B(n_308), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_360), .A2(n_323), .B1(n_337), .B2(n_318), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_392), .Y(n_402) );
OR2x6_ASAP7_75t_L g403 ( .A(n_388), .B(n_374), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_385), .A2(n_345), .B1(n_368), .B2(n_373), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_381), .B(n_131), .C(n_350), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_392), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_397), .B(n_345), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_384), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_383), .B(n_358), .Y(n_409) );
NAND2xp33_ASAP7_75t_SL g410 ( .A(n_377), .B(n_353), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_399), .B(n_369), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_394), .B(n_131), .C(n_353), .Y(n_412) );
NAND4xp75_ASAP7_75t_L g413 ( .A(n_394), .B(n_359), .C(n_367), .D(n_366), .Y(n_413) );
AO21x1_ASAP7_75t_L g414 ( .A1(n_398), .A2(n_361), .B(n_356), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_380), .B(n_370), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_391), .B(n_369), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_384), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_391), .Y(n_418) );
OAI211xp5_ASAP7_75t_SL g419 ( .A1(n_376), .A2(n_346), .B(n_362), .C(n_293), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_379), .A2(n_373), .B1(n_343), .B2(n_370), .C(n_369), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_378), .B(n_353), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_353), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_400), .B(n_308), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_400), .B(n_308), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_389), .A2(n_266), .B(n_283), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_400), .B(n_326), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_427), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_421), .B(n_382), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_425), .B(n_400), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_421), .B(n_382), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
AOI21xp5_ASAP7_75t_SL g439 ( .A1(n_404), .A2(n_395), .B(n_389), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_430), .B(n_393), .Y(n_442) );
OAI221xp5_ASAP7_75t_SL g443 ( .A1(n_415), .A2(n_386), .B1(n_390), .B2(n_401), .C(n_396), .Y(n_443) );
INVx5_ASAP7_75t_L g444 ( .A(n_403), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_427), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_431), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_407), .B(n_313), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_431), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_430), .B(n_393), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_426), .B(n_388), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_417), .B(n_8), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_422), .B(n_9), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_422), .B(n_10), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_423), .B(n_11), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_409), .Y(n_455) );
INVx5_ASAP7_75t_L g456 ( .A(n_403), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_416), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_420), .A2(n_337), .B1(n_308), .B2(n_318), .C(n_323), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_429), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_403), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_416), .Y(n_462) );
NOR2x1p5_ASAP7_75t_L g463 ( .A(n_408), .B(n_337), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_419), .B(n_11), .C(n_12), .D(n_13), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_424), .B(n_12), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_411), .B(n_13), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_411), .B(n_337), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_411), .B(n_17), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_403), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_424), .B(n_17), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_405), .B(n_322), .C(n_313), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_410), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_451), .B(n_428), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_465), .B(n_412), .C(n_410), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_455), .B(n_413), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_444), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_432), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_442), .B(n_413), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_476), .A2(n_322), .B(n_313), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_467), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_449), .B(n_414), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_434), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_440), .Y(n_490) );
NAND2xp33_ASAP7_75t_L g491 ( .A(n_444), .B(n_261), .Y(n_491) );
AOI32xp33_ASAP7_75t_L g492 ( .A1(n_467), .A2(n_18), .A3(n_19), .B1(n_335), .B2(n_274), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_449), .B(n_18), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_435), .B(n_19), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_457), .B(n_322), .Y(n_495) );
AND2x4_ASAP7_75t_SL g496 ( .A(n_461), .B(n_258), .Y(n_496) );
INVx5_ASAP7_75t_L g497 ( .A(n_444), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_444), .B(n_322), .Y(n_498) );
NAND2xp33_ASAP7_75t_SL g499 ( .A(n_461), .B(n_261), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_464), .B(n_227), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_469), .Y(n_502) );
NAND4xp25_ASAP7_75t_SL g503 ( .A(n_472), .B(n_322), .C(n_313), .D(n_326), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_452), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_435), .B(n_20), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_464), .B(n_23), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_458), .B(n_24), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_432), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_458), .B(n_26), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_462), .B(n_28), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_448), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_462), .B(n_452), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_453), .B(n_270), .Y(n_513) );
NOR4xp25_ASAP7_75t_SL g514 ( .A(n_443), .B(n_326), .C(n_33), .D(n_40), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_444), .B(n_261), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_448), .Y(n_516) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_463), .B(n_231), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_453), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_473), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_438), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_437), .B(n_30), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_445), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_437), .B(n_218), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_447), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_471), .B(n_41), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g526 ( .A(n_456), .B(n_242), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_456), .B(n_242), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_445), .B(n_44), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_446), .B(n_181), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_504), .A2(n_456), .B1(n_447), .B2(n_450), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_486), .A2(n_473), .B1(n_466), .B2(n_454), .C(n_439), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_479), .A2(n_447), .B(n_456), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_518), .B(n_441), .Y(n_533) );
NAND3xp33_ASAP7_75t_L g534 ( .A(n_492), .B(n_454), .C(n_441), .Y(n_534) );
AOI31xp33_ASAP7_75t_SL g535 ( .A1(n_481), .A2(n_456), .A3(n_436), .B(n_439), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_501), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_520), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_525), .A2(n_459), .B(n_477), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_502), .B(n_474), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_480), .Y(n_540) );
NOR2xp67_ASAP7_75t_L g541 ( .A(n_497), .B(n_446), .Y(n_541) );
AOI322xp5_ASAP7_75t_L g542 ( .A1(n_494), .A2(n_477), .A3(n_468), .B1(n_474), .B2(n_475), .C1(n_470), .C2(n_460), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_488), .Y(n_543) );
AOI21xp33_ASAP7_75t_SL g544 ( .A1(n_498), .A2(n_468), .B(n_46), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_519), .B(n_45), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_497), .A2(n_326), .B1(n_284), .B2(n_274), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_478), .A2(n_254), .B1(n_246), .B2(n_283), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_493), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_494), .B(n_208), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_489), .Y(n_550) );
AOI222xp33_ASAP7_75t_L g551 ( .A1(n_487), .A2(n_254), .B1(n_246), .B2(n_326), .C1(n_208), .C2(n_191), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_490), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_522), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_491), .A2(n_270), .B(n_277), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_522), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_512), .B(n_47), .Y(n_556) );
OAI22xp33_ASAP7_75t_SL g557 ( .A1(n_482), .A2(n_48), .B1(n_49), .B2(n_51), .Y(n_557) );
NAND3xp33_ASAP7_75t_SL g558 ( .A(n_514), .B(n_277), .C(n_282), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_497), .B(n_56), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_484), .A2(n_185), .B(n_191), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_523), .B(n_185), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_483), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_508), .Y(n_565) );
OAI22xp33_ASAP7_75t_SL g566 ( .A1(n_497), .A2(n_57), .B1(n_59), .B2(n_63), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_511), .B(n_68), .Y(n_567) );
NOR3xp33_ASAP7_75t_SL g568 ( .A(n_503), .B(n_326), .C(n_202), .Y(n_568) );
O2A1O1Ixp5_ASAP7_75t_L g569 ( .A1(n_498), .A2(n_282), .B(n_284), .C(n_237), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_516), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_505), .B(n_200), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_505), .A2(n_200), .B(n_202), .Y(n_574) );
OAI211xp5_ASAP7_75t_SL g575 ( .A1(n_513), .A2(n_237), .B(n_202), .C(n_225), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
NOR2xp33_ASAP7_75t_R g577 ( .A(n_561), .B(n_497), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_564), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_537), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_533), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_540), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_543), .B(n_550), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_541), .B(n_499), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_552), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_553), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g586 ( .A1(n_548), .A2(n_521), .A3(n_517), .B1(n_506), .B2(n_507), .C1(n_509), .C2(n_527), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_555), .B(n_521), .Y(n_587) );
XNOR2xp5_ASAP7_75t_L g588 ( .A(n_539), .B(n_531), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_563), .B(n_529), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_557), .A2(n_500), .B(n_510), .Y(n_590) );
INVx3_ASAP7_75t_SL g591 ( .A(n_559), .Y(n_591) );
INVx3_ASAP7_75t_SL g592 ( .A(n_559), .Y(n_592) );
NOR4xp25_ASAP7_75t_SL g593 ( .A(n_544), .B(n_515), .C(n_491), .D(n_524), .Y(n_593) );
NAND4xp25_ASAP7_75t_SL g594 ( .A(n_542), .B(n_485), .C(n_506), .D(n_509), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_568), .B(n_526), .Y(n_595) );
NOR4xp25_ASAP7_75t_SL g596 ( .A(n_538), .B(n_524), .C(n_496), .D(n_526), .Y(n_596) );
NOR3xp33_ASAP7_75t_SL g597 ( .A(n_532), .B(n_534), .C(n_530), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_573), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_565), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_562), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_570), .B(n_571), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_530), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_532), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_574), .B(n_496), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_578), .Y(n_607) );
OAI22xp33_ASAP7_75t_SL g608 ( .A1(n_591), .A2(n_545), .B1(n_549), .B2(n_572), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_594), .A2(n_538), .B1(n_560), .B2(n_507), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_597), .A2(n_574), .B(n_575), .C(n_528), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_602), .B(n_551), .Y(n_611) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_588), .B(n_547), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_597), .A2(n_566), .B(n_554), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g614 ( .A1(n_590), .A2(n_535), .B(n_546), .C(n_558), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_591), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_582), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_603), .B(n_567), .C(n_528), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_592), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_580), .B(n_500), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_594), .A2(n_200), .B1(n_202), .B2(n_225), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_598), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_590), .A2(n_245), .B(n_258), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_611), .A2(n_592), .B1(n_605), .B2(n_600), .Y(n_623) );
OAI31xp33_ASAP7_75t_L g624 ( .A1(n_615), .A2(n_583), .A3(n_604), .B(n_605), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_609), .A2(n_596), .B(n_593), .C(n_586), .Y(n_625) );
AOI21xp33_ASAP7_75t_SL g626 ( .A1(n_618), .A2(n_606), .B(n_576), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_612), .B(n_579), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_616), .B(n_584), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_613), .A2(n_595), .B(n_581), .C(n_585), .Y(n_629) );
CKINVDCx6p67_ASAP7_75t_R g630 ( .A(n_607), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_608), .A2(n_577), .B(n_587), .C(n_589), .Y(n_631) );
AND4x1_ASAP7_75t_L g632 ( .A(n_614), .B(n_599), .C(n_601), .D(n_245), .Y(n_632) );
AOI221xp5_ASAP7_75t_SL g633 ( .A1(n_609), .A2(n_245), .B1(n_258), .B2(n_621), .C(n_622), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_610), .A2(n_245), .B1(n_617), .B2(n_619), .Y(n_634) );
NOR3xp33_ASAP7_75t_SL g635 ( .A(n_618), .B(n_613), .C(n_594), .Y(n_635) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_609), .A2(n_597), .B(n_620), .Y(n_636) );
XOR2xp5_ASAP7_75t_L g637 ( .A(n_618), .B(n_612), .Y(n_637) );
BUFx2_ASAP7_75t_L g638 ( .A(n_630), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_628), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_628), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_636), .B(n_635), .Y(n_641) );
BUFx4f_ASAP7_75t_SL g642 ( .A(n_637), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_641), .A2(n_625), .B1(n_634), .B2(n_627), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_638), .B(n_629), .C(n_633), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_639), .A2(n_624), .B1(n_632), .B2(n_631), .C(n_623), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_644), .B(n_642), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_643), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_646), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_647), .B(n_645), .C(n_642), .Y(n_649) );
AO21x2_ASAP7_75t_L g650 ( .A1(n_649), .A2(n_640), .B(n_626), .Y(n_650) );
endmodule