module fake_netlist_1_6313_n_699 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_699);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_699;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g77 ( .A(n_69), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_30), .Y(n_78) );
BUFx3_ASAP7_75t_L g79 ( .A(n_33), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_53), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_22), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_23), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_39), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_0), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_76), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_73), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_58), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_8), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_44), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_61), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_38), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_25), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_34), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_0), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_19), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_40), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_42), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_6), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_18), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_37), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_59), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
OR2x2_ASAP7_75t_L g112 ( .A(n_67), .B(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_60), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_4), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_15), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_21), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_17), .Y(n_118) );
NOR2xp67_ASAP7_75t_L g119 ( .A(n_74), .B(n_49), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_45), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_72), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_63), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_82), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_85), .B(n_1), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_99), .Y(n_130) );
NOR2xp33_ASAP7_75t_R g131 ( .A(n_78), .B(n_28), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g132 ( .A(n_83), .B(n_29), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_109), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_91), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_96), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_106), .B(n_2), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_98), .B(n_2), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_102), .B(n_3), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_109), .Y(n_145) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_123), .B(n_32), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_79), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_104), .B(n_3), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_92), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_93), .A2(n_35), .B(n_70), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_107), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_110), .B(n_4), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_99), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_81), .B(n_71), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_85), .B(n_5), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_118), .A2(n_5), .B1(n_7), .B2(n_9), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_81), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_88), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_108), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_88), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_99), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_94), .B(n_7), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_101), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_99), .Y(n_167) );
OAI22xp33_ASAP7_75t_L g168 ( .A1(n_135), .A2(n_89), .B1(n_112), .B2(n_109), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_160), .B(n_124), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_133), .B(n_103), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_159), .Y(n_176) );
NAND3x1_ASAP7_75t_L g177 ( .A(n_158), .B(n_89), .C(n_121), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_125), .B(n_124), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_129), .B(n_108), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_163), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_125), .B(n_120), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_127), .B(n_90), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_127), .B(n_77), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_128), .B(n_137), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_126), .A2(n_77), .B1(n_90), .B2(n_100), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_150), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_129), .B(n_121), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_128), .B(n_100), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_137), .B(n_111), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_145), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_136), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_141), .B(n_147), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_158), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_157), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_141), .B(n_122), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_143), .B(n_95), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_148), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_152), .Y(n_209) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_132), .B(n_112), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_152), .B(n_114), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_153), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_145), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_130), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_130), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
BUFx4f_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_139), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_161), .B(n_105), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_165), .B(n_113), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_140), .B(n_117), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_142), .B(n_117), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_130), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_149), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_201), .Y(n_231) );
INVx6_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_230), .B(n_146), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_212), .B(n_154), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_166), .B1(n_156), .B2(n_86), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_218), .B(n_79), .Y(n_238) );
OAI22xp33_ASAP7_75t_L g239 ( .A1(n_202), .A2(n_109), .B1(n_166), .B2(n_151), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_189), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_185), .B(n_80), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_170), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_201), .B(n_80), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_220), .B(n_119), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_227), .B(n_109), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_203), .B(n_195), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_221), .B(n_151), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_178), .A2(n_151), .B(n_155), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_181), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_190), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_178), .A2(n_167), .B(n_164), .C(n_155), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_186), .A2(n_167), .B(n_164), .C(n_155), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_227), .B(n_151), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_227), .B(n_155), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_180), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_187), .B(n_10), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_181), .Y(n_263) );
NOR2x2_ASAP7_75t_L g264 ( .A(n_176), .B(n_13), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_179), .B(n_155), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_184), .B(n_144), .Y(n_266) );
OAI22xp5_ASAP7_75t_SL g267 ( .A1(n_202), .A2(n_200), .B1(n_182), .B2(n_188), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_220), .A2(n_167), .B(n_164), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_190), .B(n_167), .Y(n_269) );
BUFx12f_ASAP7_75t_L g270 ( .A(n_188), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_180), .A2(n_144), .B1(n_130), .B2(n_164), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_190), .B(n_13), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_180), .Y(n_273) );
NOR2xp33_ASAP7_75t_SL g274 ( .A(n_210), .B(n_144), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g275 ( .A(n_210), .B(n_144), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_183), .B(n_144), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_217), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_226), .B(n_167), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_173), .B(n_14), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_180), .A2(n_167), .B1(n_15), .B2(n_16), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_228), .B(n_14), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_205), .B(n_16), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_207), .B(n_50), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_209), .B(n_17), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_199), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_223), .B(n_18), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_199), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_194), .B(n_180), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_180), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_SL g293 ( .A1(n_225), .A2(n_52), .B(n_66), .C(n_26), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_197), .B(n_19), .Y(n_294) );
NAND2x1_ASAP7_75t_L g295 ( .A(n_208), .B(n_55), .Y(n_295) );
AND2x6_ASAP7_75t_SL g296 ( .A(n_200), .B(n_20), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_272), .A2(n_177), .B1(n_197), .B2(n_206), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_261), .B(n_208), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_233), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_261), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_236), .B(n_174), .Y(n_306) );
AND3x1_ASAP7_75t_SL g307 ( .A(n_264), .B(n_177), .C(n_168), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_250), .B(n_211), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_272), .A2(n_204), .B1(n_192), .B2(n_198), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_272), .A2(n_192), .B1(n_198), .B2(n_213), .Y(n_310) );
AOI21x1_ASAP7_75t_L g311 ( .A1(n_253), .A2(n_229), .B(n_224), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_231), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_239), .A2(n_169), .B(n_213), .C(n_193), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_231), .Y(n_314) );
AOI21xp33_ASAP7_75t_L g315 ( .A1(n_274), .A2(n_169), .B(n_193), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_231), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_261), .B(n_172), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_280), .A2(n_172), .B1(n_175), .B2(n_191), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_255), .A2(n_191), .B1(n_175), .B2(n_229), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_292), .B(n_250), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_231), .B(n_20), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_234), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_249), .Y(n_323) );
O2A1O1Ixp5_ASAP7_75t_SL g324 ( .A1(n_247), .A2(n_222), .B(n_219), .C(n_224), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_290), .B(n_27), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_260), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_235), .B(n_36), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_239), .A2(n_216), .B(n_214), .C(n_51), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_248), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_258), .A2(n_216), .B(n_214), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_232), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_234), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_240), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_294), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_269), .A2(n_219), .B(n_222), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_240), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_273), .B(n_222), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_252), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_267), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_269), .A2(n_219), .B(n_222), .Y(n_341) );
CKINVDCx6p67_ASAP7_75t_R g342 ( .A(n_270), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_232), .Y(n_343) );
BUFx2_ASAP7_75t_SL g344 ( .A(n_273), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_290), .B(n_41), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_259), .B(n_43), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_237), .B(n_56), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_330), .A2(n_251), .B(n_265), .Y(n_351) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_313), .A2(n_278), .B(n_282), .C(n_283), .Y(n_352) );
OR2x6_ASAP7_75t_L g353 ( .A(n_344), .B(n_270), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_306), .A2(n_286), .B(n_288), .C(n_242), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_306), .B(n_262), .Y(n_355) );
OAI22xp5_ASAP7_75t_SL g356 ( .A1(n_340), .A2(n_264), .B1(n_294), .B2(n_280), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_342), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_297), .A2(n_275), .B1(n_246), .B2(n_238), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_329), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_335), .A2(n_259), .B1(n_275), .B2(n_232), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_339), .A2(n_287), .B1(n_289), .B2(n_284), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_305), .B(n_284), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_328), .B(n_281), .C(n_247), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_308), .A2(n_279), .B1(n_276), .B2(n_266), .C(n_285), .Y(n_364) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_342), .B(n_340), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_311), .A2(n_295), .B(n_268), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_311), .A2(n_285), .B(n_263), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_339), .A2(n_243), .B1(n_263), .B2(n_254), .Y(n_369) );
AO31x2_ASAP7_75t_L g370 ( .A1(n_298), .A2(n_257), .A3(n_256), .B(n_254), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_324), .A2(n_241), .B(n_243), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_324), .A2(n_241), .B(n_271), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_301), .Y(n_373) );
OA21x2_ASAP7_75t_L g374 ( .A1(n_336), .A2(n_257), .B(n_256), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_308), .B(n_296), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_310), .A2(n_293), .B1(n_219), .B2(n_222), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_298), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_318), .B(n_271), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_309), .B(n_293), .Y(n_379) );
AOI33xp33_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_307), .A3(n_326), .B1(n_325), .B2(n_323), .B3(n_337), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_356), .A2(n_325), .B1(n_347), .B2(n_344), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_352), .A2(n_303), .B(n_341), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_375), .A2(n_325), .B1(n_345), .B2(n_321), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_377), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_303), .B(n_327), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_355), .A2(n_333), .B1(n_337), .B2(n_334), .C(n_322), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_368), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_375), .A2(n_314), .B(n_312), .Y(n_389) );
OA21x2_ASAP7_75t_L g390 ( .A1(n_371), .A2(n_346), .B(n_315), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_353), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_373), .B(n_334), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_354), .A2(n_333), .B1(n_322), .B2(n_312), .C(n_316), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_358), .A2(n_332), .B1(n_312), .B2(n_343), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_361), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_348), .B(n_316), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_358), .A2(n_319), .B1(n_343), .B2(n_299), .C(n_338), .Y(n_399) );
AO31x2_ASAP7_75t_L g400 ( .A1(n_379), .A2(n_343), .A3(n_299), .B(n_302), .Y(n_400) );
INVx4_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_365), .A2(n_302), .B1(n_304), .B2(n_331), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_353), .B(n_304), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_357), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_361), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_317), .B(n_302), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_384), .B(n_370), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_400), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_387), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_384), .B(n_370), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_404), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_400), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_400), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_384), .B(n_370), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_388), .B(n_367), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_388), .B(n_370), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_400), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_388), .B(n_351), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_394), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_391), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_391), .B(n_374), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_397), .B(n_369), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_397), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_398), .B(n_360), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_405), .B(n_374), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_405), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_389), .B(n_369), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_381), .B(n_374), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_390), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_390), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_390), .Y(n_440) );
NAND2x1_ASAP7_75t_L g441 ( .A(n_401), .B(n_302), .Y(n_441) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_407), .A2(n_372), .B(n_366), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_425), .Y(n_446) );
AOI322xp5_ASAP7_75t_L g447 ( .A1(n_422), .A2(n_381), .A3(n_392), .B1(n_383), .B2(n_386), .C1(n_376), .C2(n_396), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_409), .B(n_401), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_425), .B(n_406), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_425), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_437), .B(n_406), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_437), .B(n_406), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_414), .B(n_389), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_434), .B(n_401), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_441), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_408), .B(n_406), .Y(n_456) );
BUFx8_ASAP7_75t_L g457 ( .A(n_427), .Y(n_457) );
OAI321xp33_ASAP7_75t_L g458 ( .A1(n_434), .A2(n_392), .A3(n_395), .B1(n_403), .B2(n_399), .C(n_402), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_392), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_430), .B(n_401), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_435), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_436), .A2(n_395), .B1(n_399), .B2(n_386), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_433), .A2(n_403), .B1(n_387), .B2(n_363), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_408), .B(n_387), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_433), .A2(n_382), .B1(n_364), .B2(n_385), .C(n_387), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_429), .B(n_382), .Y(n_468) );
OAI33xp33_ASAP7_75t_L g469 ( .A1(n_431), .A2(n_378), .A3(n_385), .B1(n_65), .B2(n_68), .B3(n_62), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_429), .B(n_390), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_411), .B(n_390), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_411), .B(n_407), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_429), .B(n_299), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_416), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_419), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_419), .B(n_302), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_428), .A2(n_57), .B1(n_219), .B2(n_331), .C(n_423), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_432), .B(n_331), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_410), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_413), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_413), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_415), .B(n_331), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_427), .B(n_331), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_432), .B(n_423), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_415), .B(n_423), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_415), .B(n_420), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_418), .B(n_420), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_410), .B(n_418), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_428), .B(n_421), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_471), .B(n_418), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_471), .B(n_420), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_443), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_475), .B(n_421), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_488), .B(n_439), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_473), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_488), .B(n_439), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_459), .B(n_417), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_472), .B(n_439), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_472), .B(n_438), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_460), .B(n_438), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_444), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_475), .B(n_421), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_489), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_460), .B(n_438), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_477), .B(n_440), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_474), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_455), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_444), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_454), .B(n_469), .C(n_453), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_459), .B(n_417), .Y(n_516) );
NOR2xp67_ASAP7_75t_SL g517 ( .A(n_458), .B(n_410), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_489), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_485), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_474), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_477), .B(n_417), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_450), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_478), .B(n_440), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_450), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_480), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_478), .B(n_440), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_484), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_451), .B(n_417), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_451), .B(n_421), .Y(n_531) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_446), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_490), .B(n_410), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_452), .B(n_442), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_457), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_463), .A2(n_441), .B1(n_410), .B2(n_442), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_493), .B(n_442), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_452), .B(n_442), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_491), .B(n_410), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_446), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_490), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_470), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_456), .B(n_466), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_456), .B(n_466), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_470), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_461), .B(n_468), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_468), .B(n_449), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_449), .Y(n_550) );
INVx4_ASAP7_75t_L g551 ( .A(n_448), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_461), .B(n_465), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_509), .B(n_463), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_509), .B(n_479), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_518), .B(n_462), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_515), .A2(n_445), .B1(n_467), .B2(n_464), .C(n_462), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_496), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_518), .B(n_447), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_539), .B(n_448), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_515), .A2(n_457), .B1(n_448), .B2(n_445), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_494), .B(n_482), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_539), .B(n_457), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_494), .B(n_482), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_543), .B(n_479), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_528), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_543), .B(n_455), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_538), .B(n_492), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_536), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_494), .B(n_483), .Y(n_573) );
OAI211xp5_ASAP7_75t_L g574 ( .A1(n_536), .A2(n_481), .B(n_483), .C(n_476), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_528), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_495), .B(n_483), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_495), .B(n_486), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_552), .A2(n_486), .B1(n_476), .B2(n_487), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_498), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_538), .B(n_486), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_544), .B(n_486), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_552), .A2(n_487), .B1(n_522), .B2(n_516), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_551), .B(n_521), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
AOI31xp33_ASAP7_75t_L g585 ( .A1(n_513), .A2(n_537), .A3(n_550), .B(n_546), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_500), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_544), .B(n_547), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_495), .B(n_546), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_507), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_507), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_551), .B(n_519), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_514), .Y(n_592) );
NOR2x1_ASAP7_75t_R g593 ( .A(n_551), .B(n_513), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_522), .A2(n_516), .B1(n_503), .B2(n_531), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_499), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_537), .B(n_551), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_548), .B(n_550), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_514), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_522), .A2(n_503), .B1(n_516), .B2(n_531), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_547), .B(n_546), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_511), .B(n_525), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_523), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_545), .B(n_505), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_545), .B(n_505), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_553), .Y(n_605) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_593), .B(n_522), .Y(n_606) );
NOR4xp25_ASAP7_75t_L g607 ( .A(n_556), .B(n_497), .C(n_508), .D(n_523), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_560), .B(n_517), .C(n_519), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_597), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_565), .A2(n_517), .B(n_503), .C(n_516), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_587), .B(n_511), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_553), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_567), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_583), .B(n_503), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_558), .A2(n_548), .B1(n_497), .B2(n_508), .C(n_521), .Y(n_615) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_565), .B(n_526), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_597), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_600), .B(n_511), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_571), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_572), .B(n_526), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_595), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_562), .A2(n_540), .B1(n_535), .B2(n_504), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_598), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_588), .B(n_549), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_585), .A2(n_541), .B1(n_532), .B2(n_533), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_557), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_570), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_582), .A2(n_540), .B1(n_535), .B2(n_549), .C(n_505), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_588), .B(n_549), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_603), .B(n_504), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_594), .A2(n_599), .B1(n_580), .B2(n_573), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_578), .A2(n_504), .B1(n_530), .B2(n_525), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_574), .A2(n_530), .B1(n_499), .B2(n_501), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_579), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_589), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_566), .B(n_575), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_559), .A2(n_501), .B1(n_506), .B2(n_510), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_590), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_626), .B(n_603), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_607), .A2(n_596), .B1(n_604), .B2(n_568), .C(n_555), .Y(n_642) );
XNOR2x1_ASAP7_75t_L g643 ( .A(n_616), .B(n_591), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_609), .B(n_604), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_615), .A2(n_596), .B1(n_580), .B2(n_573), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_616), .A2(n_584), .B(n_554), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_606), .A2(n_601), .B1(n_554), .B2(n_577), .Y(n_648) );
AOI321xp33_ASAP7_75t_L g649 ( .A1(n_633), .A2(n_581), .A3(n_564), .B1(n_576), .B2(n_577), .C(n_561), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_617), .B(n_563), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_630), .B(n_563), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_605), .B(n_569), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_627), .A2(n_569), .B(n_532), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_635), .A2(n_634), .B1(n_623), .B2(n_612), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_619), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_621), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_613), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_631), .B(n_576), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_632), .B(n_561), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_610), .A2(n_575), .B(n_566), .Y(n_660) );
XNOR2xp5_ASAP7_75t_L g661 ( .A(n_639), .B(n_506), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_624), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_611), .B(n_592), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_643), .A2(n_608), .B(n_620), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_643), .A2(n_614), .B(n_611), .Y(n_665) );
OAI21xp33_ASAP7_75t_SL g666 ( .A1(n_646), .A2(n_618), .B(n_638), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_654), .A2(n_614), .B1(n_637), .B2(n_640), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_645), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_657), .A2(n_638), .B(n_618), .Y(n_669) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_653), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_648), .B(n_636), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_642), .B(n_629), .C(n_628), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_651), .A2(n_625), .A3(n_602), .B1(n_541), .B2(n_586), .C1(n_533), .C2(n_527), .Y(n_673) );
NOR2xp67_ASAP7_75t_SL g674 ( .A(n_660), .B(n_542), .Y(n_674) );
OAI32xp33_ASAP7_75t_L g675 ( .A1(n_646), .A2(n_527), .A3(n_586), .B1(n_506), .B2(n_510), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_652), .B(n_510), .Y(n_676) );
OAI31xp33_ASAP7_75t_L g677 ( .A1(n_661), .A2(n_500), .A3(n_502), .B(n_512), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_666), .A2(n_649), .B1(n_647), .B2(n_652), .C(n_663), .Y(n_678) );
AOI211x1_ASAP7_75t_SL g679 ( .A1(n_664), .A2(n_644), .B(n_650), .C(n_659), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_667), .A2(n_662), .B1(n_656), .B2(n_655), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_670), .B(n_641), .C(n_658), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_665), .A2(n_641), .B(n_658), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_668), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_671), .A2(n_500), .B1(n_502), .B2(n_512), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_672), .A2(n_502), .B1(n_512), .B2(n_520), .Y(n_685) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_678), .B(n_673), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g687 ( .A1(n_679), .A2(n_677), .B(n_669), .C(n_676), .Y(n_687) );
NOR3xp33_ASAP7_75t_SL g688 ( .A(n_682), .B(n_675), .C(n_677), .Y(n_688) );
NOR4xp75_ASAP7_75t_L g689 ( .A(n_681), .B(n_674), .C(n_524), .D(n_529), .Y(n_689) );
AO22x1_ASAP7_75t_L g690 ( .A1(n_686), .A2(n_683), .B1(n_685), .B2(n_684), .Y(n_690) );
NOR3xp33_ASAP7_75t_SL g691 ( .A(n_687), .B(n_680), .C(n_524), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g692 ( .A1(n_688), .A2(n_689), .B(n_524), .C(n_529), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_690), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_692), .Y(n_694) );
OAI22xp5_ASAP7_75t_SL g695 ( .A1(n_693), .A2(n_691), .B1(n_529), .B2(n_534), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_695), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_696), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_693), .B1(n_694), .B2(n_520), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_698), .A2(n_520), .B1(n_534), .B2(n_686), .Y(n_699) );
endmodule