module fake_ariane_365_n_2361 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2361);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2361;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_279;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_967;
wire n_437;
wire n_274;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_307;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_363;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_308;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_118),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_69),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_25),
.Y(n_245)
);

CKINVDCx6p67_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_42),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_65),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx11_ASAP7_75t_R g251 ( 
.A(n_36),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_26),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_123),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_84),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_77),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_120),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_33),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_5),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_33),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_42),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_180),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_128),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_223),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_119),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_75),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_52),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_186),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_39),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_126),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_63),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_132),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_75),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_124),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_88),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_164),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_181),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_159),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_185),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_13),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_101),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_20),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_220),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_93),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_153),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_63),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_210),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_146),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_211),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_69),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_87),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_234),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_152),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_138),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_121),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_122),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_61),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_222),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_214),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_32),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_78),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_105),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_8),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_154),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_189),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_56),
.Y(n_320)
);

INVxp33_ASAP7_75t_R g321 ( 
.A(n_213),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_16),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_94),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_19),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_83),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_65),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_208),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_133),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_102),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_106),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_2),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_98),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_162),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_96),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_66),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_60),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_17),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_92),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_204),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_18),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_225),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_24),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_115),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_90),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_34),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_169),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_86),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_178),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_127),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_175),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_27),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_191),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_196),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_198),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_129),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_17),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_167),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_71),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_174),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_59),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_30),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_44),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_78),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_43),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_149),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_171),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_131),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_37),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_104),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_8),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_163),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_111),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_61),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_91),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_89),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_184),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_103),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_160),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_55),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_4),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_76),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_116),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_4),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_201),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_141),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_91),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_3),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_143),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_142),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_203),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_73),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_72),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_46),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_66),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_32),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_147),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_232),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_45),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_70),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_93),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_205),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_49),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_54),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_5),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_89),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_113),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_71),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_218),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_41),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_130),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_45),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_72),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_48),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_158),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_84),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_94),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_125),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_39),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_83),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_85),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_176),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_29),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_38),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_145),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_187),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_9),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_37),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_44),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_55),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_16),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_156),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_1),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_41),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_170),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_150),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_92),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_60),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_24),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_20),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_179),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_227),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_107),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_36),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_23),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_99),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_57),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_19),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_100),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_193),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_6),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_200),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_108),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_48),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_215),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_109),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_14),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_237),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_237),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_251),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_364),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_242),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_242),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_260),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g465 ( 
.A(n_314),
.B(n_0),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_262),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_296),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_262),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_309),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_265),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_265),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_331),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_266),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_282),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_282),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_266),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_334),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_273),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_273),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_358),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_418),
.B(n_344),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_276),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_276),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_389),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_283),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_409),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_241),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_282),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_414),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_283),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_290),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_290),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_259),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_291),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_246),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_314),
.B(n_0),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_359),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_238),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_406),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_410),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_291),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_372),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_259),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_1),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_300),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_300),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_243),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_439),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_305),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_305),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_318),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_318),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_329),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_329),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_347),
.B(n_6),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_245),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_249),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_330),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_330),
.B(n_7),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_430),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_253),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_342),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_256),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_440),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_342),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_261),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_254),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_349),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_268),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_277),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_328),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_280),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_372),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_349),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_284),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_356),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_427),
.B(n_247),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_356),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_282),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_372),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_259),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_360),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_360),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_282),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_247),
.B(n_7),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_286),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_366),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_366),
.B(n_10),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_303),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_373),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_252),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_397),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_298),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_373),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_377),
.B(n_10),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_377),
.B(n_11),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_378),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_378),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_302),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_379),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_236),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_379),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_397),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_432),
.B(n_11),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_247),
.B(n_12),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_397),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_303),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_236),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_310),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_435),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_365),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_244),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_311),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_315),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_552),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_540),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_502),
.B(n_458),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_442),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_558),
.B(n_294),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_575),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_540),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_540),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_458),
.B(n_303),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_459),
.B(n_449),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_459),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_474),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_552),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_487),
.A2(n_412),
.B1(n_263),
.B2(n_269),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_463),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_466),
.B(n_449),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_475),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_475),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_521),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_466),
.B(n_326),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_468),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_468),
.B(n_453),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_470),
.B(n_326),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_488),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_470),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_509),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_471),
.B(n_473),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_473),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_488),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_476),
.B(n_478),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_545),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_476),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_489),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_545),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_479),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_326),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_482),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_482),
.B(n_348),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_483),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_483),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_485),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_460),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_490),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_490),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_491),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_491),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_492),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_494),
.B(n_348),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_494),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_501),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_501),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_481),
.B(n_453),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_505),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_505),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_507),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_542),
.B(n_348),
.Y(n_646)
);

NOR2x1_ASAP7_75t_L g647 ( 
.A(n_507),
.B(n_319),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_510),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_506),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_550),
.B(n_294),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_510),
.B(n_294),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_498),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_511),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_511),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_512),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_512),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_467),
.A2(n_412),
.B1(n_323),
.B2(n_327),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_513),
.B(n_264),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_513),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_514),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_514),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_515),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_569),
.B(n_563),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_508),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_515),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_503),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_519),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_516),
.B(n_321),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_519),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_523),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_526),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_529),
.B(n_322),
.Y(n_674)
);

OAI22x1_ASAP7_75t_SL g675 ( 
.A1(n_497),
.A2(n_457),
.B1(n_332),
.B2(n_333),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_643),
.B(n_517),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_643),
.B(n_518),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_584),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_586),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_612),
.B(n_264),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_626),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_612),
.B(n_462),
.Y(n_684)
);

BUFx6f_ASAP7_75t_SL g685 ( 
.A(n_668),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_626),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_642),
.A2(n_549),
.B1(n_556),
.B2(n_520),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_626),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_626),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_666),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_584),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_663),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_640),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_643),
.B(n_522),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_627),
.B(n_529),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_663),
.B(n_495),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_641),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_641),
.Y(n_700)
);

AND3x2_ASAP7_75t_L g701 ( 
.A(n_630),
.B(n_586),
.C(n_652),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_593),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_641),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_593),
.Y(n_704)
);

AOI22x1_ASAP7_75t_L g705 ( 
.A1(n_627),
.A2(n_361),
.B1(n_374),
.B2(n_322),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_612),
.B(n_524),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_641),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_641),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_627),
.B(n_535),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_627),
.B(n_535),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_593),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_599),
.Y(n_712)
);

XNOR2x2_ASAP7_75t_L g713 ( 
.A(n_657),
.B(n_321),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_643),
.B(n_527),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_641),
.Y(n_716)
);

BUFx4f_ASAP7_75t_L g717 ( 
.A(n_658),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_645),
.Y(n_718)
);

INVxp33_ASAP7_75t_L g719 ( 
.A(n_618),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_599),
.Y(n_720)
);

INVx5_ASAP7_75t_L g721 ( 
.A(n_658),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_599),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_645),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_612),
.B(n_530),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_637),
.B(n_656),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_635),
.B(n_531),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_666),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_623),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_645),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_623),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_650),
.B(n_537),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_666),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_650),
.B(n_537),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_637),
.B(n_656),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_600),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_600),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_664),
.B(n_244),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_600),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_609),
.B(n_469),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_585),
.A2(n_557),
.B1(n_566),
.B2(n_546),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_645),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_645),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_637),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_607),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_645),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_595),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_640),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_637),
.B(n_539),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_635),
.B(n_533),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_595),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_609),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_607),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_640),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_595),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_647),
.A2(n_567),
.B1(n_541),
.B2(n_553),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_595),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_640),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_651),
.B(n_539),
.Y(n_760)
);

INVxp33_ASAP7_75t_L g761 ( 
.A(n_618),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_640),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_640),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_669),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_656),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_601),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_657),
.A2(n_496),
.B1(n_504),
.B2(n_465),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_669),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_596),
.A2(n_324),
.B1(n_337),
.B2(n_335),
.Y(n_769)
);

AO21x2_ASAP7_75t_L g770 ( 
.A1(n_591),
.A2(n_544),
.B(n_543),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

BUFx8_ASAP7_75t_SL g772 ( 
.A(n_630),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_669),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_582),
.B(n_536),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_656),
.B(n_543),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_607),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_616),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_649),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_669),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_669),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_601),
.B(n_472),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_647),
.A2(n_565),
.B1(n_568),
.B2(n_534),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_582),
.B(n_547),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_615),
.Y(n_785)
);

AND2x2_ASAP7_75t_SL g786 ( 
.A(n_651),
.B(n_264),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_614),
.Y(n_787)
);

HB1xp67_ASAP7_75t_SL g788 ( 
.A(n_664),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_646),
.B(n_554),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_660),
.B(n_572),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_660),
.B(n_578),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_660),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_616),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_660),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_673),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_649),
.B(n_477),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_651),
.B(n_271),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_619),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_646),
.Y(n_800)
);

BUFx4f_ASAP7_75t_L g801 ( 
.A(n_658),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_673),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_614),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_590),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_592),
.B(n_548),
.C(n_544),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_673),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_673),
.B(n_579),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_592),
.B(n_548),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_668),
.A2(n_571),
.B1(n_576),
.B2(n_338),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_594),
.B(n_528),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_668),
.B(n_484),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_590),
.B(n_532),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_581),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_619),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_651),
.B(n_551),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_581),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_587),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_587),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_590),
.B(n_486),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_590),
.A2(n_555),
.B1(n_559),
.B2(n_551),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_614),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_602),
.A2(n_559),
.B1(n_560),
.B2(n_555),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_619),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_602),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_589),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_674),
.B(n_560),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_602),
.A2(n_564),
.B1(n_570),
.B2(n_562),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_674),
.B(n_562),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_614),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_614),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_614),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_596),
.A2(n_343),
.B1(n_346),
.B2(n_345),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_668),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_589),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_804),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_681),
.B(n_668),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_786),
.A2(n_668),
.B1(n_602),
.B2(n_625),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_678),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_678),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_679),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_786),
.A2(n_605),
.B1(n_638),
.B2(n_625),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_785),
.B(n_594),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_687),
.A2(n_597),
.B(n_608),
.C(n_603),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_774),
.B(n_597),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_679),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_679),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_786),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_692),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_772),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_824),
.A2(n_608),
.B1(n_610),
.B2(n_603),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_692),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_789),
.B(n_605),
.Y(n_852)
);

XNOR2xp5_ASAP7_75t_L g853 ( 
.A(n_713),
.B(n_499),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_784),
.B(n_733),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_L g855 ( 
.A(n_682),
.B(n_610),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_813),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_733),
.B(n_735),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_735),
.B(n_613),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_729),
.B(n_613),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_681),
.B(n_464),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_739),
.B(n_605),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_739),
.B(n_605),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_729),
.B(n_617),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_795),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_719),
.B(n_480),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_804),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_725),
.A2(n_615),
.B(n_598),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_731),
.B(n_625),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_692),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_702),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_731),
.A2(n_625),
.B1(n_638),
.B2(n_674),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_717),
.B(n_622),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_800),
.A2(n_638),
.B1(n_674),
.B2(n_583),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_800),
.B(n_693),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_761),
.B(n_461),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_778),
.B(n_500),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_753),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_798),
.A2(n_638),
.B1(n_583),
.B2(n_620),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_684),
.B(n_617),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_676),
.B(n_677),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_695),
.B(n_620),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_741),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_702),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_810),
.B(n_525),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_813),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_816),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_702),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_798),
.A2(n_624),
.B1(n_628),
.B2(n_621),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_715),
.B(n_621),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_816),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_726),
.B(n_624),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_704),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_795),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_704),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_693),
.B(n_628),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_684),
.B(n_631),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_796),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_804),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_804),
.B(n_727),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_817),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_760),
.B(n_631),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_682),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_760),
.B(n_633),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_815),
.B(n_633),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_727),
.B(n_634),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_815),
.B(n_634),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_817),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_704),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_826),
.B(n_636),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_818),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_682),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_826),
.B(n_636),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_828),
.B(n_824),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_751),
.B(n_639),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_742),
.A2(n_648),
.B1(n_654),
.B2(n_639),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_727),
.B(n_648),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_682),
.A2(n_655),
.B1(n_659),
.B2(n_654),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_828),
.B(n_655),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_711),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_788),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_745),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_818),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_745),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_711),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_727),
.B(n_659),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_711),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_698),
.B(n_661),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_825),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_820),
.B(n_661),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_822),
.B(n_662),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_712),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_825),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_787),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_798),
.A2(n_682),
.B1(n_832),
.B2(n_769),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_745),
.Y(n_935)
);

O2A1O1Ixp5_ASAP7_75t_L g936 ( 
.A1(n_694),
.A2(n_665),
.B(n_671),
.C(n_662),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_798),
.A2(n_665),
.B1(n_671),
.B2(n_658),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_827),
.B(n_622),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_767),
.B(n_591),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_712),
.Y(n_940)
);

AO22x2_ASAP7_75t_L g941 ( 
.A1(n_713),
.A2(n_833),
.B1(n_811),
.B2(n_685),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_SL g942 ( 
.A(n_765),
.B(n_288),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_696),
.B(n_622),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_811),
.B(n_598),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_706),
.B(n_675),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_682),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_682),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_782),
.B(n_604),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_696),
.B(n_629),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_724),
.B(n_675),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_790),
.B(n_604),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_709),
.B(n_710),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_709),
.B(n_710),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_796),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_750),
.B(n_629),
.Y(n_955)
);

NAND3xp33_ASAP7_75t_L g956 ( 
.A(n_767),
.B(n_632),
.C(n_629),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_712),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_806),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_806),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_750),
.B(n_775),
.Y(n_960)
);

AND2x6_ASAP7_75t_SL g961 ( 
.A(n_808),
.B(n_250),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_791),
.B(n_632),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_834),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_797),
.B(n_690),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_690),
.B(n_672),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_775),
.B(n_632),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_770),
.B(n_644),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_770),
.B(n_644),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_682),
.A2(n_653),
.B1(n_667),
.B2(n_644),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_770),
.B(n_653),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_834),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_725),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_736),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_798),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_807),
.B(n_653),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_720),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_736),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_720),
.Y(n_978)
);

BUFx6f_ASAP7_75t_SL g979 ( 
.A(n_798),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_770),
.B(n_667),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_808),
.B(n_765),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_765),
.Y(n_982)
);

AND2x4_ASAP7_75t_SL g983 ( 
.A(n_766),
.B(n_244),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_792),
.A2(n_670),
.B1(n_667),
.B2(n_672),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_720),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_787),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_792),
.B(n_670),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_L g988 ( 
.A(n_798),
.B(n_658),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_792),
.A2(n_672),
.B(n_670),
.C(n_361),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_802),
.B(n_564),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_802),
.B(n_570),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_690),
.B(n_573),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_802),
.B(n_573),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_L g994 ( 
.A(n_798),
.B(n_658),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_787),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_812),
.B(n_352),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_722),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_787),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_L g999 ( 
.A(n_680),
.B(n_658),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_769),
.A2(n_658),
.B1(n_574),
.B2(n_577),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_809),
.B(n_263),
.C(n_250),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_819),
.B(n_362),
.Y(n_1002)
);

INVxp33_ASAP7_75t_L g1003 ( 
.A(n_783),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_902),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_902),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_952),
.A2(n_752),
.B(n_748),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_854),
.B(n_757),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_880),
.B(n_728),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_979),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_877),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_920),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_874),
.B(n_701),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_963),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_874),
.B(n_728),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_844),
.B(n_728),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_953),
.A2(n_752),
.B(n_748),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_960),
.A2(n_752),
.B(n_748),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_L g1018 ( 
.A1(n_942),
.A2(n_694),
.B(n_755),
.C(n_762),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_902),
.B(n_717),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_847),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_882),
.B(n_832),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_867),
.A2(n_752),
.B(n_748),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_879),
.B(n_734),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_934),
.A2(n_685),
.B1(n_805),
.B2(n_574),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_936),
.A2(n_683),
.B(n_680),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_951),
.A2(n_896),
.B(n_879),
.C(n_857),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_881),
.A2(n_847),
.B1(n_971),
.B2(n_963),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_847),
.A2(n_756),
.B1(n_758),
.B2(n_734),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_860),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_971),
.A2(n_805),
.B(n_577),
.C(n_361),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_847),
.A2(n_756),
.B1(n_758),
.B2(n_734),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_920),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_943),
.A2(n_758),
.B(n_756),
.Y(n_1033)
);

BUFx4f_ASAP7_75t_L g1034 ( 
.A(n_874),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_717),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_L g1036 ( 
.A(n_865),
.B(n_762),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_949),
.A2(n_758),
.B(n_756),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_942),
.A2(n_968),
.B(n_967),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_948),
.A2(n_762),
.B(n_272),
.C(n_278),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_911),
.B(n_717),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_856),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_903),
.B(n_694),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_955),
.A2(n_686),
.B(n_683),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_948),
.B(n_685),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_885),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_903),
.B(n_939),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_836),
.B(n_685),
.Y(n_1047)
);

BUFx4f_ASAP7_75t_L g1048 ( 
.A(n_944),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_972),
.B(n_694),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_852),
.B(n_755),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_886),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_966),
.A2(n_689),
.B(n_686),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1001),
.A2(n_705),
.B1(n_538),
.B2(n_801),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_981),
.A2(n_691),
.B(n_689),
.Y(n_1054)
);

AO21x1_ASAP7_75t_L g1055 ( 
.A1(n_970),
.A2(n_699),
.B(n_691),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_890),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_913),
.A2(n_272),
.B(n_292),
.C(n_278),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_972),
.B(n_755),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1003),
.A2(n_705),
.B1(n_801),
.B2(n_737),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_842),
.A2(n_700),
.B(n_699),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_944),
.B(n_688),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_980),
.A2(n_759),
.B(n_749),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_944),
.A2(n_763),
.B1(n_764),
.B2(n_749),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_884),
.B(n_292),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_876),
.B(n_320),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_911),
.B(n_801),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_973),
.A2(n_703),
.B(n_700),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_973),
.A2(n_707),
.B(n_703),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_838),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_983),
.B(n_320),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_849),
.B(n_875),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_895),
.A2(n_336),
.B(n_341),
.C(n_339),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_977),
.B(n_868),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_977),
.A2(n_716),
.B(n_707),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_836),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_965),
.A2(n_764),
.B(n_763),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_838),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_900),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_987),
.A2(n_718),
.B(n_716),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_946),
.B(n_801),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1003),
.A2(n_737),
.B1(n_738),
.B2(n_722),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_889),
.A2(n_773),
.B(n_768),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_946),
.B(n_688),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_891),
.A2(n_374),
.B(n_393),
.C(n_322),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_907),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_861),
.A2(n_723),
.B(n_718),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_910),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_947),
.B(n_688),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_864),
.A2(n_730),
.B(n_723),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_868),
.B(n_688),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_922),
.A2(n_708),
.B1(n_714),
.B2(n_697),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_864),
.A2(n_743),
.B(n_730),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_868),
.B(n_697),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_858),
.B(n_697),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_944),
.B(n_697),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_862),
.A2(n_773),
.B1(n_779),
.B2(n_768),
.Y(n_1096)
);

OAI321xp33_ASAP7_75t_L g1097 ( 
.A1(n_1000),
.A2(n_339),
.A3(n_336),
.B1(n_341),
.B2(n_363),
.C(n_369),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_964),
.B(n_708),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_893),
.A2(n_744),
.B(n_743),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_928),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_983),
.B(n_363),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_893),
.A2(n_747),
.B(n_744),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_921),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_932),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_841),
.A2(n_714),
.B1(n_732),
.B2(n_708),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_905),
.B(n_376),
.C(n_369),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_897),
.A2(n_747),
.B(n_779),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_914),
.B(n_708),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_916),
.B(n_714),
.Y(n_1109)
);

BUFx8_ASAP7_75t_L g1110 ( 
.A(n_979),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_947),
.B(n_714),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_897),
.A2(n_781),
.B(n_780),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_927),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_901),
.B(n_732),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_904),
.B(n_732),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_974),
.B(n_721),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_974),
.B(n_732),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_962),
.A2(n_781),
.B(n_780),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_941),
.B(n_374),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_906),
.B(n_722),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_954),
.A2(n_821),
.B(n_803),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_909),
.B(n_737),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_954),
.A2(n_831),
.B(n_829),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_912),
.B(n_738),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_958),
.A2(n_821),
.B(n_803),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_918),
.B(n_738),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_925),
.B(n_803),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_873),
.B(n_740),
.Y(n_1128)
);

OAI321xp33_ASAP7_75t_L g1129 ( 
.A1(n_996),
.A2(n_404),
.A3(n_403),
.B1(n_451),
.B2(n_445),
.C(n_388),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_839),
.Y(n_1130)
);

AND2x6_ASAP7_75t_L g1131 ( 
.A(n_917),
.B(n_829),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_835),
.B(n_787),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_958),
.A2(n_821),
.B(n_803),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_933),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_840),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_859),
.B(n_740),
.Y(n_1136)
);

INVx4_ASAP7_75t_L g1137 ( 
.A(n_979),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_959),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_863),
.B(n_740),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_837),
.B(n_376),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_843),
.A2(n_403),
.B(n_404),
.C(n_388),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_871),
.B(n_746),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_959),
.A2(n_830),
.B(n_821),
.Y(n_1143)
);

AO21x1_ASAP7_75t_L g1144 ( 
.A1(n_975),
.A2(n_313),
.B(n_271),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_855),
.A2(n_830),
.B(n_829),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_878),
.B(n_746),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_982),
.B(n_830),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_990),
.B(n_991),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1002),
.B(n_830),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_855),
.A2(n_831),
.B(n_787),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_993),
.A2(n_831),
.B(n_754),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_915),
.B(n_746),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_929),
.B(n_754),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_776),
.B(n_754),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_921),
.B(n_776),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_997),
.Y(n_1156)
);

O2A1O1Ixp5_ASAP7_75t_L g1157 ( 
.A1(n_850),
.A2(n_777),
.B(n_793),
.C(n_776),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_899),
.A2(n_293),
.B1(n_370),
.B2(n_371),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_930),
.B(n_777),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_835),
.B(n_866),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_933),
.A2(n_793),
.B(n_777),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_921),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_866),
.B(n_793),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_853),
.Y(n_1164)
);

AOI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_956),
.A2(n_799),
.B(n_794),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_898),
.B(n_794),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_969),
.A2(n_799),
.B(n_794),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_840),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_923),
.B(n_799),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_823),
.B(n_814),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_923),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_992),
.A2(n_445),
.B(n_429),
.C(n_454),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_933),
.A2(n_823),
.B(n_814),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_989),
.A2(n_823),
.B(n_814),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_845),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_898),
.B(n_393),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_923),
.A2(n_405),
.B1(n_384),
.B2(n_387),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_933),
.A2(n_771),
.B(n_721),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_935),
.B(n_393),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_935),
.A2(n_408),
.B1(n_381),
.B2(n_392),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_935),
.A2(n_454),
.B(n_451),
.C(n_438),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_L g1182 ( 
.A(n_945),
.B(n_288),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_872),
.A2(n_313),
.B(n_271),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_888),
.B(n_396),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_938),
.B(n_396),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_933),
.B(n_721),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_986),
.A2(n_771),
.B(n_721),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_950),
.B(n_375),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_872),
.A2(n_771),
.B(n_721),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_846),
.B(n_396),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_846),
.B(n_431),
.Y(n_1191)
);

NOR2xp67_ASAP7_75t_L g1192 ( 
.A(n_1029),
.B(n_1011),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1188),
.A2(n_988),
.B1(n_994),
.B2(n_941),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1008),
.A2(n_995),
.B(n_986),
.Y(n_1194)
);

CKINVDCx6p67_ASAP7_75t_R g1195 ( 
.A(n_1032),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1113),
.B(n_941),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1015),
.A2(n_995),
.B(n_986),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1041),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1034),
.B(n_986),
.Y(n_1199)
);

OAI21xp33_ASAP7_75t_L g1200 ( 
.A1(n_1064),
.A2(n_382),
.B(n_380),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1014),
.B(n_986),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1026),
.A2(n_431),
.B(n_429),
.C(n_421),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1010),
.Y(n_1203)
);

O2A1O1Ixp5_ASAP7_75t_L g1204 ( 
.A1(n_1118),
.A2(n_851),
.B(n_869),
.C(n_848),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1026),
.A2(n_988),
.B(n_994),
.C(n_999),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_1034),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1014),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1021),
.B(n_941),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1022),
.A2(n_998),
.B(n_995),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1023),
.A2(n_998),
.B1(n_995),
.B2(n_937),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1007),
.B(n_961),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1073),
.Y(n_1212)
);

OR2x6_ASAP7_75t_SL g1213 ( 
.A(n_1101),
.B(n_849),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1044),
.B(n_848),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1177),
.B(n_395),
.C(n_394),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1027),
.A2(n_998),
.B(n_995),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1044),
.B(n_998),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1188),
.B(n_853),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1075),
.B(n_851),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1045),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1046),
.B(n_869),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1071),
.B(n_870),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1051),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1032),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1065),
.B(n_870),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1140),
.B(n_883),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1149),
.A2(n_999),
.B(n_883),
.C(n_985),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1047),
.B(n_998),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1039),
.A2(n_421),
.B(n_437),
.C(n_438),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1141),
.A2(n_437),
.B(n_431),
.C(n_872),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1056),
.B(n_887),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1070),
.B(n_1012),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1012),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1149),
.A2(n_894),
.B(n_892),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1164),
.B(n_399),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1084),
.A2(n_293),
.B(n_370),
.C(n_976),
.Y(n_1236)
);

OAI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1182),
.A2(n_433),
.B1(n_400),
.B2(n_401),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1078),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1048),
.A2(n_448),
.B1(n_416),
.B2(n_417),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1047),
.B(n_892),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1055),
.A2(n_908),
.B(n_894),
.Y(n_1241)
);

NAND2xp33_ASAP7_75t_L g1242 ( 
.A(n_1160),
.B(n_908),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1048),
.B(n_919),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1006),
.A2(n_924),
.B(n_919),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1047),
.B(n_924),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1016),
.A2(n_931),
.B(n_926),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1017),
.A2(n_931),
.B(n_926),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1009),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1009),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1085),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1148),
.A2(n_957),
.B(n_940),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1087),
.B(n_413),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1050),
.A2(n_985),
.B(n_978),
.C(n_976),
.Y(n_1253)
);

CKINVDCx16_ASAP7_75t_R g1254 ( 
.A(n_1119),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1036),
.B(n_940),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1050),
.A2(n_978),
.B(n_957),
.C(n_422),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1100),
.B(n_1104),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1129),
.A2(n_385),
.B(n_313),
.C(n_351),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1119),
.B(n_419),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1119),
.A2(n_248),
.B1(n_386),
.B2(n_444),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1084),
.A2(n_351),
.B(n_383),
.C(n_385),
.Y(n_1261)
);

BUFx2_ASAP7_75t_SL g1262 ( 
.A(n_1137),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_SL g1263 ( 
.A(n_1057),
.B(n_423),
.C(n_420),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1137),
.B(n_351),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1131),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1120),
.A2(n_385),
.B(n_383),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1122),
.A2(n_402),
.B(n_383),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1013),
.B(n_424),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1138),
.B(n_428),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1061),
.B(n_721),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1042),
.B(n_434),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1124),
.A2(n_407),
.B(n_402),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1180),
.A2(n_447),
.B(n_317),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1156),
.B(n_12),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1024),
.A2(n_357),
.B1(n_317),
.B2(n_282),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1126),
.A2(n_407),
.B(n_402),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1024),
.B(n_13),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1061),
.B(n_721),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1190),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1162),
.B(n_14),
.Y(n_1281)
);

OA22x2_ASAP7_75t_L g1282 ( 
.A1(n_1063),
.A2(n_407),
.B1(n_422),
.B2(n_446),
.Y(n_1282)
);

O2A1O1Ixp5_ASAP7_75t_SL g1283 ( 
.A1(n_1132),
.A2(n_248),
.B(n_386),
.C(n_614),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1145),
.A2(n_446),
.B(n_422),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1191),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1162),
.B(n_15),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1110),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1095),
.B(n_239),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1020),
.B(n_1094),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1176),
.B(n_1184),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1134),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1020),
.B(n_15),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1095),
.B(n_240),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1090),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1033),
.A2(n_446),
.B(n_580),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1168),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1130),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1037),
.A2(n_606),
.B(n_580),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1181),
.A2(n_18),
.B(n_21),
.C(n_22),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1069),
.A2(n_248),
.B1(n_386),
.B2(n_771),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1108),
.A2(n_317),
.B1(n_357),
.B2(n_771),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1049),
.A2(n_317),
.B1(n_357),
.B2(n_771),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1116),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1106),
.B(n_248),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1028),
.A2(n_611),
.B(n_606),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1110),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1103),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1136),
.B(n_21),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1179),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1081),
.B(n_386),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1035),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_R g1312 ( 
.A(n_1082),
.B(n_771),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1098),
.A2(n_317),
.B(n_357),
.C(n_257),
.Y(n_1313)
);

OAI22x1_ASAP7_75t_L g1314 ( 
.A1(n_1158),
.A2(n_455),
.B1(n_304),
.B2(n_301),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1139),
.B(n_22),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1098),
.A2(n_317),
.B(n_357),
.C(n_258),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1171),
.B(n_255),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1004),
.B(n_267),
.Y(n_1318)
);

AND2x4_ASAP7_75t_SL g1319 ( 
.A(n_1116),
.B(n_357),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1114),
.B(n_1115),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1097),
.A2(n_1109),
.B(n_1127),
.C(n_1068),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1053),
.A2(n_1059),
.B1(n_1109),
.B2(n_1127),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1031),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1081),
.B(n_23),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1093),
.Y(n_1325)
);

INVx4_ASAP7_75t_SL g1326 ( 
.A(n_1131),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1077),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1035),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1004),
.B(n_270),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1043),
.A2(n_611),
.B(n_606),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1052),
.A2(n_611),
.B(n_606),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1005),
.B(n_1053),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1147),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1175),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1185),
.B(n_1142),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1135),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1131),
.Y(n_1337)
);

OR2x6_ASAP7_75t_L g1338 ( 
.A(n_1040),
.B(n_1066),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1005),
.B(n_274),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1105),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1131),
.A2(n_354),
.B1(n_275),
.B2(n_279),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1054),
.A2(n_611),
.B(n_606),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1131),
.A2(n_367),
.B1(n_281),
.B2(n_285),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1155),
.A2(n_1169),
.B(n_1133),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1128),
.A2(n_368),
.B1(n_287),
.B2(n_289),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_SL g1346 ( 
.A(n_1030),
.B(n_295),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1135),
.Y(n_1347)
);

AOI221x1_ASAP7_75t_L g1348 ( 
.A1(n_1277),
.A2(n_1030),
.B1(n_1152),
.B2(n_1165),
.C(n_1091),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1334),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1344),
.A2(n_1150),
.B(n_1102),
.Y(n_1350)
);

AOI221x1_ASAP7_75t_L g1351 ( 
.A1(n_1322),
.A2(n_1151),
.B1(n_1161),
.B2(n_1173),
.C(n_1067),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1344),
.A2(n_1125),
.B(n_1121),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1333),
.A2(n_1132),
.B(n_1058),
.C(n_1092),
.Y(n_1353)
);

AO32x2_ASAP7_75t_L g1354 ( 
.A1(n_1275),
.A2(n_1144),
.A3(n_1183),
.B1(n_1062),
.B2(n_1038),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1195),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1209),
.A2(n_1169),
.B(n_1155),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1218),
.B(n_1072),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1340),
.A2(n_1059),
.B1(n_1146),
.B2(n_1096),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1298),
.A2(n_1123),
.B(n_1076),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1224),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1079),
.B(n_1170),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1330),
.A2(n_1074),
.B(n_1154),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1203),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1202),
.A2(n_1172),
.B(n_1147),
.C(n_1060),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1202),
.A2(n_1157),
.B(n_1163),
.C(n_1166),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1213),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1330),
.A2(n_1089),
.B(n_1099),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1198),
.Y(n_1368)
);

NAND4xp25_ASAP7_75t_L g1369 ( 
.A(n_1299),
.B(n_1143),
.C(n_1025),
.D(n_1018),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1331),
.A2(n_1107),
.B(n_1112),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1331),
.A2(n_1342),
.B(n_1209),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1219),
.B(n_1153),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1342),
.A2(n_1174),
.B(n_1167),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_SL g1374 ( 
.A1(n_1289),
.A2(n_1086),
.B(n_1159),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1278),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1306),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1205),
.A2(n_1019),
.B(n_1040),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1211),
.B(n_1083),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1321),
.A2(n_1111),
.B(n_1088),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1232),
.B(n_25),
.Y(n_1380)
);

AO31x2_ASAP7_75t_L g1381 ( 
.A1(n_1197),
.A2(n_1187),
.A3(n_1178),
.B(n_1117),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1294),
.B(n_1208),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_1287),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1207),
.B(n_1117),
.Y(n_1384)
);

AOI21xp33_ASAP7_75t_L g1385 ( 
.A1(n_1310),
.A2(n_1200),
.B(n_1304),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1320),
.A2(n_1019),
.B(n_1080),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1252),
.B(n_26),
.Y(n_1387)
);

NOR2xp67_ASAP7_75t_L g1388 ( 
.A(n_1265),
.B(n_1186),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1323),
.A2(n_1186),
.B(n_1080),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1299),
.A2(n_1066),
.B(n_1189),
.C(n_29),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1278),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1216),
.A2(n_1197),
.B(n_1194),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_SL g1393 ( 
.A1(n_1281),
.A2(n_27),
.B(n_28),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1194),
.A2(n_325),
.A3(n_307),
.B(n_252),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1207),
.B(n_297),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1220),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_L g1397 ( 
.A(n_1265),
.B(n_112),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1216),
.A2(n_252),
.B(n_307),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1234),
.A2(n_325),
.A3(n_307),
.B(n_252),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1257),
.B(n_28),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1223),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1234),
.A2(n_252),
.B(n_307),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1325),
.B(n_1233),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1288),
.B(n_31),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1227),
.A2(n_252),
.B(n_307),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1238),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1244),
.A2(n_307),
.B(n_325),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1264),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1278),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1250),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1253),
.A2(n_325),
.A3(n_606),
.B(n_580),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1324),
.A2(n_1193),
.B1(n_1346),
.B2(n_1196),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1293),
.B(n_31),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1263),
.A2(n_411),
.B1(n_306),
.B2(n_308),
.Y(n_1414)
);

BUFx12f_ASAP7_75t_L g1415 ( 
.A(n_1264),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1201),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1292),
.A2(n_34),
.B(n_35),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1244),
.A2(n_1247),
.B(n_1246),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1291),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1235),
.A2(n_325),
.B1(n_299),
.B2(n_398),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1284),
.A2(n_425),
.B(n_316),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1222),
.A2(n_426),
.B1(n_340),
.B2(n_350),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1192),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1246),
.A2(n_325),
.B(n_312),
.Y(n_1424)
);

INVx3_ASAP7_75t_SL g1425 ( 
.A(n_1264),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1247),
.A2(n_443),
.B(n_355),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1291),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1229),
.A2(n_35),
.B(n_38),
.C(n_40),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1296),
.Y(n_1429)
);

INVx3_ASAP7_75t_SL g1430 ( 
.A(n_1201),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1305),
.A2(n_450),
.B(n_390),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1206),
.B(n_114),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1308),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.C(n_47),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1286),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1230),
.A2(n_452),
.B(n_391),
.C(n_415),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1305),
.A2(n_456),
.B(n_436),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1254),
.B(n_47),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1265),
.A2(n_353),
.B1(n_441),
.B2(n_51),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1228),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1245),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1236),
.A2(n_588),
.B(n_606),
.C(n_611),
.Y(n_1441)
);

AOI221x1_ASAP7_75t_L g1442 ( 
.A1(n_1258),
.A2(n_1284),
.B1(n_1316),
.B2(n_1313),
.C(n_1273),
.Y(n_1442)
);

OAI211xp5_ASAP7_75t_L g1443 ( 
.A1(n_1239),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1212),
.B(n_50),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1265),
.B(n_1243),
.Y(n_1445)
);

AO31x2_ASAP7_75t_L g1446 ( 
.A1(n_1251),
.A2(n_611),
.A3(n_580),
.B(n_588),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1291),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1327),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1228),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_L g1450 ( 
.A(n_1215),
.B(n_588),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1259),
.A2(n_588),
.B1(n_611),
.B2(n_580),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1307),
.B(n_53),
.Y(n_1452)
);

AO32x2_ASAP7_75t_L g1453 ( 
.A1(n_1210),
.A2(n_53),
.A3(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1225),
.B(n_58),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1251),
.A2(n_580),
.B(n_588),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1242),
.A2(n_1332),
.B(n_1214),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1256),
.A2(n_580),
.B(n_588),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1315),
.A2(n_136),
.B(n_229),
.Y(n_1458)
);

OAI22x1_ASAP7_75t_L g1459 ( 
.A1(n_1341),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_1459)
);

NOR2xp67_ASAP7_75t_L g1460 ( 
.A(n_1248),
.B(n_139),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1237),
.Y(n_1461)
);

AO21x1_ASAP7_75t_L g1462 ( 
.A1(n_1217),
.A2(n_62),
.B(n_64),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1266),
.A2(n_1267),
.A3(n_1272),
.B(n_1276),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1266),
.A2(n_151),
.B(n_226),
.Y(n_1464)
);

AO32x2_ASAP7_75t_L g1465 ( 
.A1(n_1301),
.A2(n_67),
.A3(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1297),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1337),
.A2(n_67),
.B1(n_68),
.B2(n_74),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1343),
.A2(n_74),
.B(n_76),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1295),
.A2(n_166),
.B(n_221),
.Y(n_1469)
);

BUFx12f_ASAP7_75t_L g1470 ( 
.A(n_1240),
.Y(n_1470)
);

NOR2xp67_ASAP7_75t_L g1471 ( 
.A(n_1248),
.B(n_157),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1295),
.A2(n_155),
.B(n_219),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1204),
.A2(n_140),
.B(n_217),
.Y(n_1473)
);

AO32x2_ASAP7_75t_L g1474 ( 
.A1(n_1302),
.A2(n_77),
.A3(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1303),
.B(n_79),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1303),
.B(n_81),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1221),
.A2(n_173),
.B(n_216),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1240),
.Y(n_1478)
);

AOI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1267),
.A2(n_168),
.B(n_212),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1241),
.A2(n_135),
.B(n_209),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1241),
.A2(n_134),
.B(n_207),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1272),
.A2(n_1276),
.B(n_1261),
.Y(n_1482)
);

AO31x2_ASAP7_75t_L g1483 ( 
.A1(n_1347),
.A2(n_231),
.A3(n_202),
.B(n_197),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1231),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1336),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1309),
.A2(n_192),
.B(n_190),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1262),
.B(n_82),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1271),
.B(n_82),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1280),
.A2(n_177),
.A3(n_87),
.B(n_88),
.Y(n_1489)
);

BUFx5_ASAP7_75t_L g1490 ( 
.A(n_1285),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1274),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1226),
.Y(n_1492)
);

CKINVDCx6p67_ASAP7_75t_R g1493 ( 
.A(n_1314),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1318),
.A2(n_86),
.B(n_90),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1268),
.B(n_1269),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1329),
.A2(n_95),
.B(n_97),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1260),
.B(n_95),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1249),
.Y(n_1498)
);

BUFx2_ASAP7_75t_R g1499 ( 
.A(n_1199),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1319),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1339),
.A2(n_1255),
.B(n_1338),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1338),
.A2(n_1335),
.B(n_1317),
.Y(n_1502)
);

OAI22x1_ASAP7_75t_L g1503 ( 
.A1(n_1249),
.A2(n_1290),
.B1(n_1282),
.B2(n_1326),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1338),
.A2(n_1236),
.B(n_1270),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_SL g1505 ( 
.A1(n_1279),
.A2(n_1261),
.B(n_1326),
.C(n_1283),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_R g1506 ( 
.A(n_1311),
.B(n_1328),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1345),
.B(n_1311),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_SL g1508 ( 
.A1(n_1326),
.A2(n_1312),
.B(n_1328),
.C(n_1300),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1203),
.B(n_884),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1202),
.A2(n_1188),
.B(n_1193),
.C(n_854),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1207),
.B(n_1206),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1218),
.B(n_681),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1344),
.A2(n_880),
.B(n_1113),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1211),
.B(n_1021),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1298),
.A2(n_1331),
.B(n_1330),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1218),
.A2(n_739),
.B1(n_884),
.B2(n_1188),
.Y(n_1516)
);

NAND2xp33_ASAP7_75t_L g1517 ( 
.A(n_1340),
.B(n_880),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1344),
.A2(n_880),
.B(n_1008),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1197),
.A2(n_1055),
.A3(n_1118),
.B(n_1144),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1287),
.Y(n_1520)
);

NOR2x1_ASAP7_75t_R g1521 ( 
.A(n_1287),
.B(n_849),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1344),
.A2(n_880),
.B(n_1008),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1516),
.A2(n_1357),
.B1(n_1385),
.B2(n_1517),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1516),
.A2(n_1514),
.B1(n_1404),
.B2(n_1413),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1467),
.A2(n_1468),
.B(n_1497),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1493),
.A2(n_1412),
.B1(n_1459),
.B2(n_1512),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1368),
.Y(n_1527)
);

INVx5_ASAP7_75t_L g1528 ( 
.A(n_1487),
.Y(n_1528)
);

BUFx2_ASAP7_75t_SL g1529 ( 
.A(n_1500),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1519),
.Y(n_1530)
);

BUFx8_ASAP7_75t_L g1531 ( 
.A(n_1520),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1418),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1355),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1396),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1412),
.A2(n_1387),
.B1(n_1467),
.B2(n_1495),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1443),
.A2(n_1509),
.B(n_1428),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1491),
.A2(n_1461),
.B1(n_1488),
.B2(n_1513),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1380),
.B(n_1363),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1360),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1437),
.B(n_1487),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1372),
.B(n_1378),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1376),
.Y(n_1542)
);

BUFx12f_ASAP7_75t_L g1543 ( 
.A(n_1383),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1434),
.A2(n_1487),
.B1(n_1444),
.B2(n_1408),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1358),
.A2(n_1382),
.B1(n_1366),
.B2(n_1492),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1358),
.A2(n_1400),
.B1(n_1415),
.B2(n_1503),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1454),
.A2(n_1502),
.B1(n_1484),
.B2(n_1448),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1401),
.A2(n_1406),
.B1(n_1410),
.B2(n_1429),
.Y(n_1548)
);

INVx6_ASAP7_75t_L g1549 ( 
.A(n_1478),
.Y(n_1549)
);

BUFx8_ASAP7_75t_L g1550 ( 
.A(n_1453),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1510),
.A2(n_1414),
.B1(n_1422),
.B2(n_1390),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1416),
.B(n_1439),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1427),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1425),
.A2(n_1422),
.B1(n_1414),
.B2(n_1476),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1462),
.A2(n_1379),
.B1(n_1485),
.B2(n_1403),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1375),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1438),
.A2(n_1478),
.B1(n_1470),
.B2(n_1466),
.Y(n_1557)
);

CKINVDCx11_ASAP7_75t_R g1558 ( 
.A(n_1383),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1423),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1507),
.A2(n_1417),
.B1(n_1440),
.B2(n_1432),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1391),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1430),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1440),
.B(n_1416),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1511),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1511),
.Y(n_1565)
);

BUFx10_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1475),
.A2(n_1348),
.B1(n_1369),
.B2(n_1442),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1391),
.Y(n_1568)
);

INVx8_ASAP7_75t_L g1569 ( 
.A(n_1432),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1490),
.A2(n_1449),
.B1(n_1420),
.B2(n_1496),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1490),
.A2(n_1494),
.B1(n_1421),
.B2(n_1369),
.Y(n_1571)
);

INVx4_ASAP7_75t_SL g1572 ( 
.A(n_1489),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1409),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1490),
.A2(n_1421),
.B1(n_1504),
.B2(n_1453),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1453),
.A2(n_1522),
.B1(n_1518),
.B2(n_1389),
.Y(n_1576)
);

CKINVDCx11_ASAP7_75t_R g1577 ( 
.A(n_1409),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1490),
.A2(n_1464),
.B1(n_1456),
.B2(n_1501),
.Y(n_1578)
);

CKINVDCx14_ASAP7_75t_R g1579 ( 
.A(n_1521),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1419),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1490),
.A2(n_1464),
.B1(n_1384),
.B2(n_1374),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1419),
.B(n_1447),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1451),
.A2(n_1388),
.B1(n_1450),
.B2(n_1433),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1435),
.A2(n_1364),
.B1(n_1395),
.B2(n_1498),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1365),
.A2(n_1386),
.B(n_1426),
.Y(n_1585)
);

BUFx2_ASAP7_75t_SL g1586 ( 
.A(n_1419),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1447),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1447),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1506),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1515),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1465),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1498),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1506),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1465),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1465),
.Y(n_1595)
);

INVx6_ASAP7_75t_L g1596 ( 
.A(n_1521),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1388),
.A2(n_1433),
.B1(n_1350),
.B2(n_1474),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1474),
.A2(n_1397),
.B1(n_1486),
.B2(n_1458),
.Y(n_1598)
);

INVx6_ASAP7_75t_L g1599 ( 
.A(n_1499),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1397),
.B(n_1471),
.Y(n_1600)
);

AOI21xp33_ASAP7_75t_L g1601 ( 
.A1(n_1431),
.A2(n_1436),
.B(n_1482),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1441),
.A2(n_1377),
.B1(n_1356),
.B2(n_1405),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1353),
.A2(n_1352),
.B(n_1392),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1460),
.A2(n_1471),
.B1(n_1457),
.B2(n_1469),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1460),
.A2(n_1457),
.B1(n_1477),
.B2(n_1424),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1472),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1474),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1398),
.A2(n_1407),
.B1(n_1473),
.B2(n_1402),
.Y(n_1608)
);

INVx4_ASAP7_75t_L g1609 ( 
.A(n_1473),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1479),
.A2(n_1393),
.B1(n_1455),
.B2(n_1505),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1480),
.A2(n_1481),
.B1(n_1373),
.B2(n_1508),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1359),
.A2(n_1370),
.B1(n_1367),
.B2(n_1361),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1362),
.A2(n_1371),
.B1(n_1351),
.B2(n_1354),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1483),
.A2(n_1354),
.B1(n_1519),
.B2(n_1463),
.Y(n_1614)
);

CKINVDCx11_ASAP7_75t_R g1615 ( 
.A(n_1483),
.Y(n_1615)
);

BUFx12f_ASAP7_75t_L g1616 ( 
.A(n_1519),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1354),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1463),
.A2(n_1381),
.B1(n_1411),
.B2(n_1446),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1463),
.A2(n_1381),
.B1(n_1411),
.B2(n_1394),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1399),
.B(n_1394),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1411),
.A2(n_1516),
.B1(n_1218),
.B2(n_1119),
.Y(n_1621)
);

BUFx8_ASAP7_75t_L g1622 ( 
.A(n_1381),
.Y(n_1622)
);

CKINVDCx14_ASAP7_75t_R g1623 ( 
.A(n_1446),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1368),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1368),
.Y(n_1625)
);

CKINVDCx6p67_ASAP7_75t_R g1626 ( 
.A(n_1366),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1514),
.B(n_1021),
.Y(n_1627)
);

BUFx4f_ASAP7_75t_SL g1628 ( 
.A(n_1383),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1357),
.A2(n_739),
.B1(n_1218),
.B2(n_713),
.Y(n_1629)
);

CKINVDCx11_ASAP7_75t_R g1630 ( 
.A(n_1383),
.Y(n_1630)
);

CKINVDCx12_ASAP7_75t_R g1631 ( 
.A(n_1521),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1360),
.Y(n_1632)
);

BUFx12f_ASAP7_75t_L g1633 ( 
.A(n_1383),
.Y(n_1633)
);

BUFx12f_ASAP7_75t_L g1634 ( 
.A(n_1383),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1478),
.Y(n_1635)
);

BUFx10_ASAP7_75t_L g1636 ( 
.A(n_1355),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1516),
.A2(n_1404),
.B1(n_1413),
.B2(n_1340),
.Y(n_1637)
);

INVx5_ASAP7_75t_L g1638 ( 
.A(n_1487),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1639)
);

CKINVDCx11_ASAP7_75t_R g1640 ( 
.A(n_1383),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1516),
.A2(n_1467),
.B(n_1468),
.Y(n_1641)
);

BUFx8_ASAP7_75t_L g1642 ( 
.A(n_1520),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1357),
.A2(n_739),
.B1(n_1218),
.B2(n_713),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1360),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1383),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1349),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1368),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1368),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1355),
.Y(n_1650)
);

BUFx4f_ASAP7_75t_SL g1651 ( 
.A(n_1383),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1517),
.B(n_1516),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1355),
.Y(n_1653)
);

NAND2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1445),
.B(n_1265),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1360),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1349),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1368),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1658)
);

INVx3_ASAP7_75t_SL g1659 ( 
.A(n_1355),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1516),
.A2(n_1404),
.B1(n_1413),
.B2(n_1340),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1368),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1368),
.Y(n_1662)
);

INVx6_ASAP7_75t_L g1663 ( 
.A(n_1478),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1368),
.Y(n_1664)
);

INVx6_ASAP7_75t_L g1665 ( 
.A(n_1478),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1514),
.B(n_1021),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1514),
.B(n_1021),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1514),
.B(n_1021),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1368),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1514),
.B(n_1382),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1514),
.B(n_1382),
.Y(n_1672)
);

CKINVDCx11_ASAP7_75t_R g1673 ( 
.A(n_1383),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1357),
.A2(n_739),
.B1(n_1218),
.B2(n_713),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1360),
.Y(n_1675)
);

BUFx8_ASAP7_75t_L g1676 ( 
.A(n_1520),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1418),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1678)
);

CKINVDCx11_ASAP7_75t_R g1679 ( 
.A(n_1383),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1516),
.A2(n_739),
.B1(n_884),
.B2(n_1218),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1516),
.A2(n_1404),
.B1(n_1413),
.B2(n_1340),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1516),
.A2(n_1218),
.B1(n_1119),
.B2(n_596),
.Y(n_1684)
);

INVx4_ASAP7_75t_L g1685 ( 
.A(n_1355),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1357),
.A2(n_739),
.B1(n_1218),
.B2(n_713),
.Y(n_1686)
);

INVx6_ASAP7_75t_L g1687 ( 
.A(n_1478),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1375),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1375),
.Y(n_1689)
);

BUFx10_ASAP7_75t_L g1690 ( 
.A(n_1355),
.Y(n_1690)
);

CKINVDCx6p67_ASAP7_75t_R g1691 ( 
.A(n_1366),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1368),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1516),
.A2(n_739),
.B1(n_1467),
.B2(n_1340),
.Y(n_1693)
);

BUFx8_ASAP7_75t_L g1694 ( 
.A(n_1520),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1355),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1516),
.A2(n_1404),
.B1(n_1413),
.B2(n_1340),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1375),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1622),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1528),
.B(n_1638),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1527),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1617),
.B(n_1534),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1632),
.B(n_1562),
.Y(n_1702)
);

INVx11_ASAP7_75t_L g1703 ( 
.A(n_1531),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1530),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1530),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1533),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1624),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1625),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1641),
.A2(n_1693),
.B(n_1603),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1618),
.A2(n_1610),
.B(n_1608),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1648),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1649),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1661),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1662),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1664),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1670),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1692),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1572),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1602),
.A2(n_1585),
.B(n_1620),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1569),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1572),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1617),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1681),
.A2(n_1646),
.B1(n_1680),
.B2(n_1682),
.C(n_1658),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1565),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1538),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1606),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1616),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1617),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_SL g1732 ( 
.A1(n_1652),
.A2(n_1525),
.B(n_1551),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1622),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1594),
.Y(n_1734)
);

AO31x2_ASAP7_75t_L g1735 ( 
.A1(n_1595),
.A2(n_1607),
.A3(n_1609),
.B(n_1605),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1619),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1613),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1671),
.B(n_1672),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1693),
.A2(n_1660),
.B(n_1637),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1623),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1592),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1548),
.B(n_1627),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1529),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1523),
.B(n_1667),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1539),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1590),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1548),
.B(n_1668),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1590),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1612),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1532),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1569),
.B(n_1654),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1532),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1669),
.B(n_1597),
.Y(n_1753)
);

AO21x2_ASAP7_75t_L g1754 ( 
.A1(n_1567),
.A2(n_1576),
.B(n_1601),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1604),
.A2(n_1576),
.B(n_1567),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1677),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1677),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1647),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1537),
.B(n_1524),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1537),
.B(n_1524),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1580),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1644),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1639),
.A2(n_1666),
.B1(n_1658),
.B2(n_1678),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1528),
.B(n_1638),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1580),
.Y(n_1765)
);

O2A1O1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1683),
.A2(n_1696),
.B(n_1536),
.C(n_1554),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1656),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1564),
.Y(n_1768)
);

OA21x2_ASAP7_75t_L g1769 ( 
.A1(n_1614),
.A2(n_1575),
.B(n_1597),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1615),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1578),
.A2(n_1581),
.B(n_1614),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1655),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1575),
.B(n_1621),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1545),
.B(n_1563),
.Y(n_1774)
);

AOI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1584),
.A2(n_1556),
.B(n_1582),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1621),
.B(n_1545),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1535),
.B(n_1547),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1565),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_SL g1779 ( 
.A1(n_1550),
.A2(n_1528),
.B1(n_1638),
.B2(n_1599),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1550),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1581),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1547),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1528),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1638),
.B(n_1573),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1535),
.B(n_1540),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1639),
.A2(n_1682),
.B1(n_1680),
.B2(n_1666),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1542),
.B(n_1566),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1675),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1578),
.A2(n_1571),
.B(n_1600),
.Y(n_1789)
);

AO21x2_ASAP7_75t_L g1790 ( 
.A1(n_1554),
.A2(n_1552),
.B(n_1587),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1571),
.A2(n_1600),
.B(n_1598),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1559),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1552),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1611),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1697),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1697),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1611),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1697),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1573),
.Y(n_1799)
);

AOI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1553),
.A2(n_1589),
.B(n_1593),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1688),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1689),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1598),
.A2(n_1555),
.B(n_1583),
.Y(n_1803)
);

INVx1_ASAP7_75t_SL g1804 ( 
.A(n_1577),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1568),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1526),
.B(n_1678),
.Y(n_1806)
);

NAND2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1574),
.B(n_1546),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1544),
.B(n_1646),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1555),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1684),
.A2(n_1643),
.B(n_1686),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1546),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1549),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1526),
.B(n_1684),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1560),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1561),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1549),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1560),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1596),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1586),
.Y(n_1819)
);

BUFx12f_ASAP7_75t_L g1820 ( 
.A(n_1558),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1583),
.Y(n_1821)
);

OAI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1599),
.A2(n_1691),
.B1(n_1626),
.B2(n_1663),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1570),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1588),
.B(n_1570),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1544),
.B(n_1566),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1635),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1635),
.Y(n_1827)
);

NAND4xp25_ASAP7_75t_SL g1828 ( 
.A(n_1629),
.B(n_1686),
.C(n_1674),
.D(n_1643),
.Y(n_1828)
);

BUFx2_ASAP7_75t_SL g1829 ( 
.A(n_1685),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1635),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1663),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1599),
.A2(n_1674),
.B1(n_1629),
.B2(n_1663),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1665),
.Y(n_1833)
);

AOI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1557),
.A2(n_1687),
.B(n_1665),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1665),
.B(n_1687),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1557),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1596),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1596),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1531),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1642),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1631),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1543),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1642),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1676),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1676),
.Y(n_1845)
);

OA21x2_ASAP7_75t_L g1846 ( 
.A1(n_1653),
.A2(n_1695),
.B(n_1628),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1728),
.B(n_1579),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_L g1848 ( 
.A(n_1766),
.B(n_1630),
.C(n_1679),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1780),
.B(n_1659),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1700),
.Y(n_1850)
);

OR2x6_ASAP7_75t_L g1851 ( 
.A(n_1699),
.B(n_1633),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1726),
.A2(n_1763),
.B(n_1786),
.C(n_1810),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_R g1853 ( 
.A(n_1846),
.B(n_1673),
.Y(n_1853)
);

BUFx4f_ASAP7_75t_SL g1854 ( 
.A(n_1707),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1739),
.A2(n_1685),
.B1(n_1650),
.B2(n_1659),
.C(n_1694),
.Y(n_1855)
);

OA21x2_ASAP7_75t_L g1856 ( 
.A1(n_1755),
.A2(n_1711),
.B(n_1722),
.Y(n_1856)
);

OA21x2_ASAP7_75t_L g1857 ( 
.A1(n_1711),
.A2(n_1628),
.B(n_1651),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1780),
.B(n_1636),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1745),
.B(n_1636),
.Y(n_1859)
);

A2O1A1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1806),
.A2(n_1694),
.B(n_1651),
.C(n_1640),
.Y(n_1860)
);

AO32x2_ASAP7_75t_L g1861 ( 
.A1(n_1783),
.A2(n_1634),
.A3(n_1645),
.B1(n_1690),
.B2(n_1727),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1738),
.B(n_1690),
.Y(n_1862)
);

OA21x2_ASAP7_75t_L g1863 ( 
.A1(n_1722),
.A2(n_1710),
.B(n_1771),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1806),
.A2(n_1813),
.B(n_1808),
.C(n_1832),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1699),
.B(n_1764),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1828),
.A2(n_1813),
.B1(n_1732),
.B2(n_1760),
.C(n_1759),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1805),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1761),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1704),
.B(n_1782),
.Y(n_1869)
);

INVx5_ASAP7_75t_L g1870 ( 
.A(n_1751),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1762),
.B(n_1772),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1743),
.B(n_1788),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1738),
.B(n_1742),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1699),
.B(n_1764),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1708),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1741),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1699),
.B(n_1764),
.Y(n_1877)
);

OAI21x1_ASAP7_75t_SL g1878 ( 
.A1(n_1732),
.A2(n_1834),
.B(n_1846),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1742),
.B(n_1747),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1803),
.A2(n_1777),
.B(n_1821),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1733),
.B(n_1698),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1820),
.A2(n_1846),
.B1(n_1804),
.B2(n_1840),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1708),
.Y(n_1883)
);

O2A1O1Ixp33_ASAP7_75t_SL g1884 ( 
.A1(n_1822),
.A2(n_1839),
.B(n_1840),
.C(n_1844),
.Y(n_1884)
);

OR2x6_ASAP7_75t_L g1885 ( 
.A(n_1698),
.B(n_1783),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1812),
.Y(n_1886)
);

AO32x2_ASAP7_75t_L g1887 ( 
.A1(n_1727),
.A2(n_1778),
.A3(n_1816),
.B1(n_1720),
.B2(n_1701),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1782),
.B(n_1713),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1733),
.B(n_1698),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1776),
.A2(n_1777),
.B1(n_1836),
.B2(n_1821),
.Y(n_1890)
);

O2A1O1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1809),
.A2(n_1792),
.B(n_1797),
.C(n_1794),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1776),
.A2(n_1773),
.B1(n_1809),
.B2(n_1811),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1803),
.A2(n_1825),
.B(n_1794),
.C(n_1797),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1735),
.Y(n_1894)
);

INVx4_ASAP7_75t_SL g1895 ( 
.A(n_1824),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1754),
.A2(n_1748),
.B(n_1746),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1753),
.B(n_1825),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1714),
.B(n_1716),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1773),
.A2(n_1791),
.B(n_1823),
.C(n_1836),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1771),
.A2(n_1789),
.B(n_1781),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1785),
.B(n_1815),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1744),
.A2(n_1811),
.B1(n_1823),
.B2(n_1779),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1785),
.B(n_1720),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1831),
.B(n_1833),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1714),
.B(n_1716),
.Y(n_1905)
);

O2A1O1Ixp33_ASAP7_75t_L g1906 ( 
.A1(n_1754),
.A2(n_1737),
.B(n_1749),
.C(n_1781),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1709),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1774),
.A2(n_1818),
.B1(n_1824),
.B2(n_1838),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1824),
.A2(n_1737),
.B(n_1749),
.C(n_1774),
.Y(n_1909)
);

AOI21xp33_ASAP7_75t_L g1910 ( 
.A1(n_1754),
.A2(n_1769),
.B(n_1737),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1824),
.A2(n_1814),
.B1(n_1817),
.B2(n_1837),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1768),
.B(n_1826),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1709),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1787),
.B(n_1845),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1845),
.B(n_1843),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1768),
.B(n_1826),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1843),
.B(n_1844),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1712),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1827),
.B(n_1830),
.Y(n_1919)
);

OAI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1775),
.A2(n_1769),
.B(n_1817),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1820),
.A2(n_1846),
.B1(n_1841),
.B2(n_1835),
.Y(n_1921)
);

CKINVDCx20_ASAP7_75t_R g1922 ( 
.A(n_1842),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1717),
.B(n_1718),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1793),
.B(n_1730),
.Y(n_1924)
);

NAND2xp33_ASAP7_75t_R g1925 ( 
.A(n_1818),
.B(n_1841),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1746),
.A2(n_1757),
.B(n_1752),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1795),
.B(n_1796),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1801),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1796),
.B(n_1798),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1816),
.B(n_1702),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1802),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1712),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1748),
.A2(n_1750),
.B(n_1752),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1793),
.B(n_1730),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1798),
.B(n_1715),
.Y(n_1935)
);

AO32x2_ASAP7_75t_L g1936 ( 
.A1(n_1778),
.A2(n_1735),
.A3(n_1814),
.B1(n_1734),
.B2(n_1790),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1703),
.Y(n_1937)
);

AND2x4_ASAP7_75t_SL g1938 ( 
.A(n_1723),
.B(n_1842),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1719),
.B(n_1770),
.Y(n_1939)
);

CKINVDCx20_ASAP7_75t_R g1940 ( 
.A(n_1842),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1784),
.B(n_1790),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1734),
.B(n_1705),
.Y(n_1942)
);

O2A1O1Ixp5_ASAP7_75t_SL g1943 ( 
.A1(n_1750),
.A2(n_1757),
.B(n_1756),
.C(n_1819),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1769),
.A2(n_1736),
.B(n_1705),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1873),
.B(n_1735),
.Y(n_1945)
);

INVxp67_ASAP7_75t_SL g1946 ( 
.A(n_1894),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1942),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1926),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1942),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1879),
.B(n_1735),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1903),
.B(n_1731),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1876),
.B(n_1850),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1904),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1926),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1928),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_1878),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1869),
.B(n_1735),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1875),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1871),
.B(n_1706),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1883),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1854),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1928),
.B(n_1706),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1887),
.B(n_1725),
.Y(n_1963)
);

INVx4_ASAP7_75t_L g1964 ( 
.A(n_1851),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1907),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1866),
.A2(n_1740),
.B1(n_1769),
.B2(n_1736),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1936),
.Y(n_1967)
);

NOR2x1p5_ASAP7_75t_L g1968 ( 
.A(n_1867),
.B(n_1834),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1860),
.B(n_1842),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1922),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1887),
.B(n_1897),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1936),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1936),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1900),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1914),
.B(n_1842),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1849),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1901),
.B(n_1939),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1900),
.Y(n_1978)
);

OAI222xp33_ASAP7_75t_L g1979 ( 
.A1(n_1892),
.A2(n_1740),
.B1(n_1807),
.B2(n_1800),
.C1(n_1767),
.C2(n_1758),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1931),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1866),
.A2(n_1736),
.B1(n_1807),
.B2(n_1724),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1913),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1918),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1932),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1863),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1892),
.A2(n_1807),
.B1(n_1721),
.B2(n_1724),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1863),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1931),
.B(n_1756),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1935),
.Y(n_1989)
);

INVx2_ASAP7_75t_SL g1990 ( 
.A(n_1885),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1862),
.B(n_1829),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1865),
.B(n_1729),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1865),
.B(n_1729),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1874),
.B(n_1877),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1898),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1852),
.A2(n_1829),
.B1(n_1819),
.B2(n_1723),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1898),
.Y(n_1997)
);

AND3x2_ASAP7_75t_L g1998 ( 
.A(n_1848),
.B(n_1784),
.C(n_1799),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1905),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1905),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1923),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1923),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1874),
.B(n_1729),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1885),
.Y(n_2004)
);

INVx4_ASAP7_75t_L g2005 ( 
.A(n_1851),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1912),
.B(n_1729),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1916),
.B(n_1927),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1888),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1888),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1994),
.B(n_1895),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1971),
.B(n_1859),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1995),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1957),
.B(n_1947),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1948),
.Y(n_2014)
);

AOI221xp5_ASAP7_75t_L g2015 ( 
.A1(n_1967),
.A2(n_1910),
.B1(n_1906),
.B2(n_1891),
.C(n_1902),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1971),
.B(n_1886),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1994),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1995),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1997),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1997),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1947),
.B(n_1896),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1950),
.B(n_1880),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1955),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_1966),
.B(n_1848),
.C(n_1896),
.Y(n_2024)
);

OAI321xp33_ASAP7_75t_L g2025 ( 
.A1(n_1981),
.A2(n_1902),
.A3(n_1864),
.B1(n_1880),
.B2(n_1893),
.C(n_1909),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1949),
.B(n_1933),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_2007),
.B(n_1856),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1977),
.B(n_1856),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1948),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1956),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1977),
.B(n_1857),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1949),
.B(n_1933),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1999),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1956),
.Y(n_2034)
);

AOI31xp33_ASAP7_75t_L g2035 ( 
.A1(n_1996),
.A2(n_1853),
.A3(n_1855),
.B(n_1884),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1994),
.B(n_1857),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1964),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1948),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2008),
.B(n_1943),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1956),
.Y(n_2040)
);

OAI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_1986),
.A2(n_1909),
.B1(n_1899),
.B2(n_1891),
.C(n_1890),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_1994),
.Y(n_2042)
);

INVxp67_ASAP7_75t_L g2043 ( 
.A(n_1980),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_2004),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1950),
.B(n_1944),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_1945),
.B(n_1944),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1948),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1954),
.Y(n_2048)
);

AOI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_1979),
.A2(n_1910),
.B1(n_1906),
.B2(n_1882),
.C(n_1855),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1999),
.Y(n_2050)
);

AO22x1_ASAP7_75t_L g2051 ( 
.A1(n_1970),
.A2(n_1881),
.B1(n_1889),
.B2(n_1870),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1954),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2000),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1954),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2000),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_2004),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1953),
.B(n_1917),
.Y(n_2057)
);

AOI211xp5_ASAP7_75t_L g2058 ( 
.A1(n_1969),
.A2(n_1921),
.B(n_1908),
.C(n_1920),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2001),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1964),
.Y(n_2060)
);

INVx5_ASAP7_75t_SL g2061 ( 
.A(n_1992),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1953),
.B(n_1872),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2008),
.B(n_1920),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_1970),
.Y(n_2064)
);

AOI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_1967),
.A2(n_1908),
.B1(n_1915),
.B2(n_1911),
.C(n_1930),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1967),
.A2(n_1934),
.B1(n_1924),
.B2(n_1941),
.Y(n_2066)
);

NAND3xp33_ASAP7_75t_L g2067 ( 
.A(n_1985),
.B(n_1858),
.C(n_1919),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_1976),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1951),
.B(n_1847),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2009),
.B(n_1929),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2001),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1968),
.B(n_1895),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2002),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2012),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_2026),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2042),
.B(n_1970),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2042),
.B(n_2006),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2039),
.B(n_1958),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2039),
.B(n_1958),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_2061),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2063),
.B(n_1960),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2012),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2031),
.B(n_2006),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2063),
.B(n_1960),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2018),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_2035),
.B(n_1975),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_2024),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2026),
.B(n_1965),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_2032),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2013),
.B(n_1945),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_2032),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2031),
.B(n_2017),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2048),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2017),
.B(n_1992),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2018),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2048),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_2064),
.B(n_1937),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2013),
.B(n_1988),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2070),
.B(n_1988),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_2010),
.B(n_1964),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2070),
.B(n_1962),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2036),
.B(n_1992),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2036),
.B(n_1992),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2019),
.B(n_1965),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2061),
.B(n_1993),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2061),
.B(n_1993),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2019),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_2064),
.B(n_1703),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2023),
.B(n_1959),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2020),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2020),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2061),
.B(n_1993),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2033),
.B(n_1982),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2033),
.B(n_1982),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2061),
.B(n_1993),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2048),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2011),
.B(n_2003),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2050),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_2010),
.B(n_2034),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_2050),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2053),
.B(n_1983),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_2010),
.B(n_1964),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2052),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2053),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2011),
.B(n_2003),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2045),
.B(n_1952),
.Y(n_2126)
);

AND2x4_ASAP7_75t_L g2127 ( 
.A(n_2010),
.B(n_2005),
.Y(n_2127)
);

NAND2xp33_ASAP7_75t_L g2128 ( 
.A(n_2068),
.B(n_1961),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2055),
.B(n_2059),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2045),
.B(n_1989),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2016),
.B(n_2003),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_2034),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2055),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2095),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2095),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_2087),
.B(n_2035),
.Y(n_2136)
);

NOR2x1p5_ASAP7_75t_L g2137 ( 
.A(n_2080),
.B(n_2024),
.Y(n_2137)
);

NAND3xp33_ASAP7_75t_L g2138 ( 
.A(n_2087),
.B(n_2049),
.C(n_2015),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2119),
.B(n_2034),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2120),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_2078),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2086),
.A2(n_2058),
.B1(n_2041),
.B2(n_2065),
.Y(n_2142)
);

INVx1_ASAP7_75t_SL g2143 ( 
.A(n_2128),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2075),
.B(n_2043),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2120),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2093),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2075),
.B(n_2089),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2089),
.B(n_2068),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2074),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2086),
.B(n_2030),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2093),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2126),
.B(n_2022),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2078),
.A2(n_2049),
.B1(n_2041),
.B2(n_2065),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2074),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2093),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2126),
.B(n_2022),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2091),
.Y(n_2157)
);

NOR2xp67_ASAP7_75t_L g2158 ( 
.A(n_2080),
.B(n_2067),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2119),
.B(n_2030),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2096),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2082),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2119),
.B(n_2040),
.Y(n_2162)
);

NAND2x1p5_ASAP7_75t_L g2163 ( 
.A(n_2080),
.B(n_2005),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2082),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2091),
.B(n_2028),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2079),
.B(n_2028),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2101),
.B(n_2046),
.Y(n_2167)
);

INVx6_ASAP7_75t_L g2168 ( 
.A(n_2119),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2105),
.B(n_2040),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2085),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2085),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2107),
.Y(n_2172)
);

OR2x2_ASAP7_75t_SL g2173 ( 
.A(n_2130),
.B(n_2067),
.Y(n_2173)
);

OAI21xp33_ASAP7_75t_L g2174 ( 
.A1(n_2079),
.A2(n_2027),
.B(n_2044),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2107),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2110),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2110),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2099),
.B(n_2021),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2111),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2111),
.Y(n_2180)
);

INVx4_ASAP7_75t_L g2181 ( 
.A(n_2132),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2101),
.B(n_2027),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2118),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2118),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2130),
.B(n_2046),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2105),
.B(n_2056),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2099),
.B(n_2044),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2124),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2124),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2109),
.B(n_2059),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2149),
.Y(n_2191)
);

NAND2xp33_ASAP7_75t_R g2192 ( 
.A(n_2150),
.B(n_2136),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2154),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2136),
.B(n_2081),
.Y(n_2194)
);

NAND2x1_ASAP7_75t_L g2195 ( 
.A(n_2168),
.B(n_2132),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2161),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2153),
.B(n_2081),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2164),
.Y(n_2198)
);

NAND4xp25_ASAP7_75t_L g2199 ( 
.A(n_2138),
.B(n_2132),
.C(n_2108),
.D(n_2076),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2167),
.B(n_2088),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2170),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2173),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2152),
.B(n_2088),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2171),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2172),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_2150),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_SL g2207 ( 
.A1(n_2142),
.A2(n_1973),
.B1(n_1972),
.B2(n_2072),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2141),
.B(n_2084),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2141),
.B(n_2084),
.Y(n_2209)
);

NAND3xp33_ASAP7_75t_L g2210 ( 
.A(n_2157),
.B(n_2147),
.C(n_2135),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2157),
.B(n_2098),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2175),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2146),
.Y(n_2213)
);

INVx1_ASAP7_75t_SL g2214 ( 
.A(n_2143),
.Y(n_2214)
);

NAND4xp25_ASAP7_75t_L g2215 ( 
.A(n_2158),
.B(n_2132),
.C(n_2076),
.D(n_2097),
.Y(n_2215)
);

NAND2x1p5_ASAP7_75t_L g2216 ( 
.A(n_2137),
.B(n_2080),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2139),
.B(n_2100),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2146),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2151),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2156),
.B(n_2098),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2139),
.B(n_2100),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2159),
.B(n_2100),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2159),
.B(n_2100),
.Y(n_2223)
);

NAND4xp75_ASAP7_75t_L g2224 ( 
.A(n_2148),
.B(n_2025),
.C(n_2092),
.D(n_2021),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2151),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2162),
.B(n_2122),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2185),
.B(n_2129),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2162),
.B(n_2122),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2176),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2169),
.B(n_2122),
.Y(n_2230)
);

NAND2xp33_ASAP7_75t_SL g2231 ( 
.A(n_2169),
.B(n_2106),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_2174),
.A2(n_2058),
.B1(n_2072),
.B2(n_1968),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2155),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2197),
.B(n_2144),
.Y(n_2234)
);

OAI21xp5_ASAP7_75t_L g2235 ( 
.A1(n_2224),
.A2(n_2025),
.B(n_2163),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2202),
.A2(n_2168),
.B1(n_2163),
.B2(n_2187),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2202),
.Y(n_2237)
);

OAI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_2224),
.A2(n_2140),
.B(n_2134),
.Y(n_2238)
);

AOI32xp33_ASAP7_75t_L g2239 ( 
.A1(n_2207),
.A2(n_2166),
.A3(n_2165),
.B1(n_2186),
.B2(n_2182),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2198),
.Y(n_2240)
);

NAND4xp25_ASAP7_75t_L g2241 ( 
.A(n_2192),
.B(n_2181),
.C(n_2145),
.D(n_2186),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2198),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_2195),
.Y(n_2243)
);

AOI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_2194),
.A2(n_2178),
.B1(n_1973),
.B2(n_1972),
.C(n_2155),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2216),
.B(n_2230),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2206),
.A2(n_2168),
.B1(n_2178),
.B2(n_2122),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2214),
.Y(n_2247)
);

CKINVDCx20_ASAP7_75t_R g2248 ( 
.A(n_2231),
.Y(n_2248)
);

OAI21xp33_ASAP7_75t_L g2249 ( 
.A1(n_2199),
.A2(n_2190),
.B(n_2179),
.Y(n_2249)
);

AOI221xp5_ASAP7_75t_L g2250 ( 
.A1(n_2210),
.A2(n_1973),
.B1(n_1972),
.B2(n_2160),
.C(n_2189),
.Y(n_2250)
);

INVx1_ASAP7_75t_SL g2251 ( 
.A(n_2231),
.Y(n_2251)
);

OAI221xp5_ASAP7_75t_SL g2252 ( 
.A1(n_2232),
.A2(n_2090),
.B1(n_2092),
.B2(n_2014),
.C(n_2038),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2216),
.B(n_2181),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2220),
.B(n_2177),
.Y(n_2254)
);

NOR2x1_ASAP7_75t_L g2255 ( 
.A(n_2215),
.B(n_2181),
.Y(n_2255)
);

OAI322xp33_ASAP7_75t_L g2256 ( 
.A1(n_2216),
.A2(n_2188),
.A3(n_2184),
.B1(n_2183),
.B2(n_2180),
.C1(n_2090),
.C2(n_2047),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2230),
.B(n_2127),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2208),
.A2(n_2129),
.B(n_2127),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2220),
.B(n_2133),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2201),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2217),
.B(n_2221),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_2217),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2211),
.B(n_2133),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2247),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2247),
.B(n_2200),
.Y(n_2265)
);

AOI21xp33_ASAP7_75t_SL g2266 ( 
.A1(n_2235),
.A2(n_2236),
.B(n_2239),
.Y(n_2266)
);

OAI322xp33_ASAP7_75t_L g2267 ( 
.A1(n_2234),
.A2(n_2209),
.A3(n_2200),
.B1(n_2203),
.B2(n_2227),
.C1(n_2204),
.C2(n_2201),
.Y(n_2267)
);

OAI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_2241),
.A2(n_2203),
.B1(n_2204),
.B2(n_2212),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2240),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2262),
.B(n_2191),
.Y(n_2270)
);

AOI222xp33_ASAP7_75t_L g2271 ( 
.A1(n_2244),
.A2(n_2233),
.B1(n_2213),
.B2(n_2218),
.C1(n_2219),
.C2(n_2225),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2262),
.B(n_2193),
.Y(n_2272)
);

AOI211xp5_ASAP7_75t_SL g2273 ( 
.A1(n_2248),
.A2(n_2223),
.B(n_2228),
.C(n_2222),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2238),
.A2(n_2195),
.B(n_2212),
.Y(n_2274)
);

NOR4xp25_ASAP7_75t_L g2275 ( 
.A(n_2237),
.B(n_2196),
.C(n_2229),
.D(n_2205),
.Y(n_2275)
);

AOI221xp5_ASAP7_75t_L g2276 ( 
.A1(n_2250),
.A2(n_2233),
.B1(n_2213),
.B2(n_2218),
.C(n_2225),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2242),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2237),
.A2(n_2219),
.B1(n_2160),
.B2(n_1985),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2261),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2260),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2248),
.A2(n_2221),
.B1(n_2228),
.B2(n_2226),
.Y(n_2281)
);

OAI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2251),
.A2(n_2227),
.B(n_2223),
.Y(n_2282)
);

INVx2_ASAP7_75t_SL g2283 ( 
.A(n_2261),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2256),
.A2(n_2226),
.B(n_2222),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2254),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2249),
.B(n_2083),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2283),
.B(n_2258),
.Y(n_2287)
);

XNOR2xp5_ASAP7_75t_L g2288 ( 
.A(n_2279),
.B(n_2245),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2279),
.B(n_2245),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2264),
.B(n_2259),
.Y(n_2290)
);

O2A1O1Ixp33_ASAP7_75t_L g2291 ( 
.A1(n_2266),
.A2(n_2252),
.B(n_2243),
.C(n_2246),
.Y(n_2291)
);

AOI221xp5_ASAP7_75t_L g2292 ( 
.A1(n_2275),
.A2(n_2263),
.B1(n_2257),
.B2(n_2243),
.C(n_2253),
.Y(n_2292)
);

INVx1_ASAP7_75t_SL g2293 ( 
.A(n_2265),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2268),
.B(n_2255),
.Y(n_2294)
);

A2O1A1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2274),
.A2(n_2276),
.B(n_2284),
.C(n_2273),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2268),
.A2(n_2257),
.B1(n_2253),
.B2(n_2014),
.C(n_2047),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2286),
.A2(n_2037),
.B1(n_2060),
.B2(n_2047),
.Y(n_2297)
);

AOI222xp33_ASAP7_75t_L g2298 ( 
.A1(n_2278),
.A2(n_2116),
.B1(n_2096),
.B2(n_2123),
.C1(n_2054),
.C2(n_2052),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2270),
.B(n_2109),
.Y(n_2299)
);

XNOR2x1_ASAP7_75t_L g2300 ( 
.A(n_2282),
.B(n_1998),
.Y(n_2300)
);

INVxp33_ASAP7_75t_L g2301 ( 
.A(n_2281),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_2293),
.B(n_2267),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2293),
.A2(n_2271),
.B1(n_2300),
.B2(n_2295),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2289),
.Y(n_2304)
);

NOR4xp25_ASAP7_75t_L g2305 ( 
.A(n_2294),
.B(n_2280),
.C(n_2277),
.D(n_2269),
.Y(n_2305)
);

NOR3xp33_ASAP7_75t_SL g2306 ( 
.A(n_2288),
.B(n_2272),
.C(n_2285),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2301),
.B(n_2102),
.Y(n_2307)
);

BUFx10_ASAP7_75t_L g2308 ( 
.A(n_2292),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2299),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2290),
.Y(n_2310)
);

HB1xp67_ASAP7_75t_L g2311 ( 
.A(n_2287),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2297),
.B(n_2278),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2291),
.B(n_2127),
.Y(n_2313)
);

NAND2xp33_ASAP7_75t_L g2314 ( 
.A(n_2296),
.B(n_2106),
.Y(n_2314)
);

OAI221xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2298),
.A2(n_2038),
.B1(n_2029),
.B2(n_2014),
.C(n_2056),
.Y(n_2315)
);

NAND3xp33_ASAP7_75t_L g2316 ( 
.A(n_2295),
.B(n_2060),
.C(n_2037),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2304),
.Y(n_2317)
);

AOI32xp33_ASAP7_75t_L g2318 ( 
.A1(n_2302),
.A2(n_2029),
.A3(n_2038),
.B1(n_2127),
.B2(n_2083),
.Y(n_2318)
);

NOR3xp33_ASAP7_75t_SL g2319 ( 
.A(n_2316),
.B(n_1991),
.C(n_1925),
.Y(n_2319)
);

AOI211xp5_ASAP7_75t_L g2320 ( 
.A1(n_2305),
.A2(n_2029),
.B(n_2112),
.C(n_2115),
.Y(n_2320)
);

AOI222xp33_ASAP7_75t_L g2321 ( 
.A1(n_2308),
.A2(n_2123),
.B1(n_2096),
.B2(n_2116),
.C1(n_2054),
.C2(n_2052),
.Y(n_2321)
);

OR2x2_ASAP7_75t_L g2322 ( 
.A(n_2309),
.B(n_2104),
.Y(n_2322)
);

OAI221xp5_ASAP7_75t_L g2323 ( 
.A1(n_2303),
.A2(n_2123),
.B1(n_2116),
.B2(n_1987),
.C(n_1985),
.Y(n_2323)
);

AOI221xp5_ASAP7_75t_L g2324 ( 
.A1(n_2306),
.A2(n_1987),
.B1(n_2054),
.B2(n_1974),
.C(n_1978),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2311),
.A2(n_2104),
.B1(n_2113),
.B2(n_2121),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2307),
.B(n_2102),
.Y(n_2326)
);

AOI321xp33_ASAP7_75t_L g2327 ( 
.A1(n_2313),
.A2(n_2072),
.A3(n_2066),
.B1(n_1987),
.B2(n_1946),
.C(n_1881),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2320),
.A2(n_2312),
.B1(n_2310),
.B2(n_2315),
.Y(n_2328)
);

OAI222xp33_ASAP7_75t_L g2329 ( 
.A1(n_2323),
.A2(n_2315),
.B1(n_2308),
.B2(n_2314),
.C1(n_1940),
.C2(n_2037),
.Y(n_2329)
);

OAI221xp5_ASAP7_75t_L g2330 ( 
.A1(n_2324),
.A2(n_2037),
.B1(n_2060),
.B2(n_2121),
.C(n_2113),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2317),
.A2(n_2114),
.B(n_2062),
.Y(n_2331)
);

O2A1O1Ixp33_ASAP7_75t_L g2332 ( 
.A1(n_2321),
.A2(n_2114),
.B(n_2071),
.C(n_2073),
.Y(n_2332)
);

OAI221xp5_ASAP7_75t_R g2333 ( 
.A1(n_2318),
.A2(n_2077),
.B1(n_2131),
.B2(n_2060),
.C(n_1861),
.Y(n_2333)
);

OAI211xp5_ASAP7_75t_L g2334 ( 
.A1(n_2322),
.A2(n_2112),
.B(n_2115),
.C(n_2077),
.Y(n_2334)
);

INVx2_ASAP7_75t_SL g2335 ( 
.A(n_2326),
.Y(n_2335)
);

NOR4xp25_ASAP7_75t_L g2336 ( 
.A(n_2327),
.B(n_2062),
.C(n_2071),
.D(n_2073),
.Y(n_2336)
);

NAND4xp75_ASAP7_75t_L g2337 ( 
.A(n_2335),
.B(n_2319),
.C(n_2325),
.D(n_2103),
.Y(n_2337)
);

INVxp33_ASAP7_75t_SL g2338 ( 
.A(n_2328),
.Y(n_2338)
);

XNOR2xp5_ASAP7_75t_L g2339 ( 
.A(n_2336),
.B(n_2072),
.Y(n_2339)
);

AOI22xp5_ASAP7_75t_L g2340 ( 
.A1(n_2330),
.A2(n_2103),
.B1(n_2016),
.B2(n_1978),
.Y(n_2340)
);

NAND4xp75_ASAP7_75t_L g2341 ( 
.A(n_2331),
.B(n_2333),
.C(n_2329),
.D(n_2334),
.Y(n_2341)
);

NOR2x1_ASAP7_75t_L g2342 ( 
.A(n_2332),
.B(n_2094),
.Y(n_2342)
);

NOR2x1_ASAP7_75t_L g2343 ( 
.A(n_2328),
.B(n_2094),
.Y(n_2343)
);

OAI32xp33_ASAP7_75t_L g2344 ( 
.A1(n_2338),
.A2(n_2341),
.A3(n_2337),
.B1(n_2343),
.B2(n_2339),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2342),
.B(n_2057),
.Y(n_2345)
);

OAI221xp5_ASAP7_75t_L g2346 ( 
.A1(n_2340),
.A2(n_2005),
.B1(n_1978),
.B2(n_1974),
.C(n_1861),
.Y(n_2346)
);

OAI211xp5_ASAP7_75t_SL g2347 ( 
.A1(n_2343),
.A2(n_1861),
.B(n_1990),
.C(n_1984),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2347),
.A2(n_1974),
.B1(n_1889),
.B2(n_1963),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_2345),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2349),
.Y(n_2350)
);

OAI22xp5_ASAP7_75t_SL g2351 ( 
.A1(n_2350),
.A2(n_2349),
.B1(n_2344),
.B2(n_2346),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_SL g2352 ( 
.A1(n_2350),
.A2(n_2348),
.B1(n_2005),
.B2(n_1990),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2351),
.A2(n_2069),
.B(n_2125),
.Y(n_2353)
);

AOI21xp33_ASAP7_75t_SL g2354 ( 
.A1(n_2352),
.A2(n_2051),
.B(n_2125),
.Y(n_2354)
);

OAI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2353),
.A2(n_2354),
.B1(n_2069),
.B2(n_2117),
.Y(n_2355)
);

NOR3xp33_ASAP7_75t_L g2356 ( 
.A(n_2353),
.B(n_2051),
.C(n_1800),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2355),
.A2(n_2356),
.B(n_2117),
.Y(n_2357)
);

OAI21xp5_ASAP7_75t_SL g2358 ( 
.A1(n_2357),
.A2(n_1938),
.B(n_2057),
.Y(n_2358)
);

XNOR2xp5_ASAP7_75t_L g2359 ( 
.A(n_2358),
.B(n_2131),
.Y(n_2359)
);

OAI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2359),
.A2(n_1723),
.B1(n_1765),
.B2(n_1761),
.C(n_1868),
.Y(n_2360)
);

AOI211xp5_ASAP7_75t_L g2361 ( 
.A1(n_2360),
.A2(n_1723),
.B(n_1765),
.C(n_1761),
.Y(n_2361)
);


endmodule