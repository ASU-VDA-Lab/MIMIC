module fake_jpeg_11917_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx10_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_5),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_2),
.B1(n_3),
.B2(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_24),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_11),
.B1(n_16),
.B2(n_10),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_16),
.Y(n_25)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_7),
.CI(n_13),
.CON(n_32),
.SN(n_32)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_36),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_29),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_28),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_42),
.B(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_32),
.B1(n_28),
.B2(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.C(n_38),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_41),
.B(n_38),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.A3(n_31),
.B1(n_17),
.B2(n_27),
.C1(n_21),
.C2(n_23),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_31),
.C(n_27),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_17),
.Y(n_49)
);


endmodule