module fake_jpeg_2855_n_74 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_23),
.B1(n_24),
.B2(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_22),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_29),
.B(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_27),
.C(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_33),
.B(n_24),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_24),
.B1(n_33),
.B2(n_27),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_11),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_7),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_2),
.C(n_6),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_10),
.B(n_11),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_61),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_62),
.C(n_52),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_7),
.B(n_8),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_15),
.C(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_65),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_60),
.C(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OAI322xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_64),
.A3(n_52),
.B1(n_17),
.B2(n_18),
.C1(n_20),
.C2(n_14),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_13),
.Y(n_74)
);


endmodule