module fake_jpeg_26687_n_204 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_12),
.B1(n_16),
.B2(n_21),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_11),
.B1(n_16),
.B2(n_22),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_24),
.A3(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_42)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_52),
.CI(n_15),
.CON(n_67),
.SN(n_67)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_40),
.B1(n_34),
.B2(n_16),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_48),
.B1(n_53),
.B2(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_51),
.Y(n_64)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_18),
.B1(n_23),
.B2(n_17),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_34),
.B1(n_39),
.B2(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_13),
.B1(n_21),
.B2(n_20),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_23),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_32),
.B(n_30),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_61),
.B1(n_63),
.B2(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_33),
.B(n_18),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_49),
.C(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_23),
.B1(n_36),
.B2(n_33),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_23),
.B1(n_36),
.B2(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_42),
.CI(n_51),
.CON(n_75),
.SN(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_63),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_62),
.B1(n_67),
.B2(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_57),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_58),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_65),
.C(n_67),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_74),
.C(n_75),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_73),
.B1(n_75),
.B2(n_61),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_62),
.B1(n_61),
.B2(n_57),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_68),
.B1(n_66),
.B2(n_49),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_63),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_83),
.B1(n_79),
.B2(n_72),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_108),
.B1(n_120),
.B2(n_18),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_78),
.B1(n_61),
.B2(n_76),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_117),
.B(n_90),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_0),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_19),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_73),
.B1(n_61),
.B2(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_70),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_69),
.B(n_58),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_86),
.C(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_125),
.C(n_140),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_86),
.C(n_94),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_111),
.B(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_106),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_131),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_32),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_135),
.B1(n_102),
.B2(n_110),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_19),
.B1(n_17),
.B2(n_2),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_0),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_0),
.C(n_1),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_119),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_149),
.B1(n_151),
.B2(n_132),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_113),
.B1(n_110),
.B2(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_140),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_128),
.C(n_125),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_1),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_163),
.B(n_1),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_130),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_161),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_134),
.C(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_139),
.C(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_143),
.B1(n_142),
.B2(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_160),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_148),
.B1(n_144),
.B2(n_154),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_176),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_153),
.B(n_2),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_173),
.B(n_3),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_3),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_165),
.B1(n_159),
.B2(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_183),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_3),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_4),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_4),
.B(n_5),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_10),
.C(n_5),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_172),
.B(n_175),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_6),
.B(n_7),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_189),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_184),
.A2(n_181),
.B1(n_175),
.B2(n_8),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_6),
.C(n_7),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_8),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_194),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_201),
.A3(n_188),
.B1(n_199),
.B2(n_190),
.C1(n_8),
.C2(n_9),
.Y(n_202)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_192),
.B(n_187),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_8),
.B(n_9),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_9),
.Y(n_204)
);


endmodule