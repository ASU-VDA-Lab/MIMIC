module fake_jpeg_31833_n_100 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_10),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_17),
.B1(n_14),
.B2(n_21),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_28),
.B1(n_27),
.B2(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_21),
.B1(n_25),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_46),
.B1(n_19),
.B2(n_26),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_25),
.C(n_28),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_26),
.Y(n_59)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_52),
.B1(n_42),
.B2(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_27),
.B1(n_26),
.B2(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_0),
.Y(n_64)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_12),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_26),
.B1(n_23),
.B2(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_7),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_62),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_63),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_12),
.C(n_19),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_40),
.Y(n_71)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_55),
.B1(n_58),
.B2(n_63),
.C(n_52),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_59),
.C(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_57),
.B1(n_50),
.B2(n_52),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_78),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_76),
.C(n_75),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_89),
.C(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_66),
.B1(n_82),
.B2(n_81),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_66),
.C(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_73),
.B1(n_51),
.B2(n_41),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_52),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_94),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_3),
.B(n_5),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g98 ( 
.A(n_97),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_8),
.Y(n_100)
);


endmodule