module fake_jpeg_10753_n_476 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_476);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_133;
wire n_419;
wire n_132;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_26),
.B(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_54),
.B(n_58),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_91),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_66),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g118 ( 
.A(n_67),
.Y(n_118)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_94),
.Y(n_107)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_78),
.Y(n_109)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_80),
.Y(n_151)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_85),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_11),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_89),
.B(n_92),
.Y(n_134)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_23),
.B1(n_38),
.B2(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_11),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_29),
.B(n_0),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_100),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_24),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_20),
.B1(n_15),
.B2(n_34),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_103),
.A2(n_117),
.B1(n_127),
.B2(n_141),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_20),
.B1(n_34),
.B2(n_43),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_104),
.A2(n_158),
.B1(n_93),
.B2(n_88),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_34),
.B1(n_14),
.B2(n_41),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_117),
.A2(n_127),
.B1(n_141),
.B2(n_67),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_126),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_14),
.B1(n_41),
.B2(n_43),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_61),
.A2(n_14),
.B1(n_41),
.B2(n_43),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_90),
.A2(n_37),
.B(n_29),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_155),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_51),
.A2(n_37),
.B1(n_24),
.B2(n_44),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_153),
.B1(n_157),
.B2(n_67),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_56),
.A2(n_24),
.B1(n_44),
.B2(n_23),
.Y(n_153)
);

AO22x2_ASAP7_75t_L g157 ( 
.A1(n_49),
.A2(n_38),
.B1(n_33),
.B2(n_32),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_63),
.A2(n_32),
.B1(n_13),
.B2(n_25),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_171),
.B1(n_177),
.B2(n_156),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_0),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_167),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_0),
.Y(n_167)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_69),
.B1(n_99),
.B2(n_74),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_92),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_175),
.A2(n_59),
.B1(n_55),
.B2(n_156),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_176),
.A2(n_188),
.B1(n_197),
.B2(n_203),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_66),
.B1(n_64),
.B2(n_91),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_118),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_179),
.A2(n_170),
.B1(n_196),
.B2(n_190),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_116),
.Y(n_180)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_100),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_182),
.B(n_123),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_128),
.A2(n_100),
.B1(n_61),
.B2(n_72),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g186 ( 
.A(n_118),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_79),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_190),
.Y(n_210)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_0),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_108),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_0),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_2),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_82),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_196),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_201),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_60),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_2),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_2),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_223),
.B1(n_113),
.B2(n_130),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_165),
.B(n_139),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_145),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_236),
.B1(n_180),
.B2(n_109),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_154),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_189),
.A2(n_144),
.B1(n_115),
.B2(n_106),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_124),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_182),
.Y(n_247)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_209),
.B1(n_234),
.B2(n_200),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_239),
.A2(n_258),
.B1(n_266),
.B2(n_229),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_181),
.B(n_193),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_246),
.B(n_216),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_181),
.C(n_173),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_249),
.C(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_200),
.B1(n_175),
.B2(n_171),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_245),
.B1(n_259),
.B2(n_261),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_164),
.B(n_200),
.C(n_236),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_248),
.Y(n_279)
);

NOR2x1p5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_182),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_166),
.C(n_167),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_172),
.B(n_194),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_265),
.B(n_221),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_161),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_163),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_220),
.A2(n_191),
.B1(n_184),
.B2(n_110),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_177),
.B1(n_144),
.B2(n_115),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_211),
.B(n_169),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_106),
.B1(n_140),
.B2(n_86),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_160),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_262),
.Y(n_293)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_208),
.B(n_198),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_210),
.B1(n_230),
.B2(n_218),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_269),
.B1(n_282),
.B2(n_284),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_216),
.B1(n_228),
.B2(n_208),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_273),
.A2(n_290),
.B(n_257),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_246),
.A2(n_203),
.B1(n_226),
.B2(n_147),
.Y(n_282)
);

OAI22x1_ASAP7_75t_SL g285 ( 
.A1(n_246),
.A2(n_232),
.B1(n_235),
.B2(n_180),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_248),
.Y(n_311)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_292),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_226),
.B1(n_147),
.B2(n_238),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_289),
.A2(n_243),
.B1(n_261),
.B2(n_262),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_245),
.A2(n_235),
.B1(n_232),
.B2(n_214),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_240),
.A2(n_214),
.B(n_229),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_291),
.B(n_248),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_265),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_241),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_272),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_257),
.C(n_249),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_286),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_304),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_253),
.B(n_256),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_299),
.A2(n_309),
.B(n_312),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_250),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_305),
.C(n_310),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_260),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_302),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_277),
.A2(n_239),
.B1(n_252),
.B2(n_244),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_303),
.A2(n_289),
.B1(n_285),
.B2(n_282),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_279),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_279),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_268),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_307),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_255),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_311),
.A2(n_315),
.B(n_318),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_247),
.B(n_244),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_259),
.B1(n_293),
.B2(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_219),
.B(n_224),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_263),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_295),
.B(n_274),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_334),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_306),
.B(n_217),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_327),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_325),
.A2(n_309),
.B1(n_315),
.B2(n_316),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_308),
.A2(n_319),
.B1(n_277),
.B2(n_299),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_328),
.A2(n_330),
.B1(n_332),
.B2(n_270),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_290),
.B1(n_293),
.B2(n_285),
.Y(n_330)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_312),
.B1(n_303),
.B2(n_302),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_267),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_281),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_339),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_271),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_217),
.Y(n_340)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_314),
.B(n_280),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_271),
.C(n_288),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_346),
.C(n_317),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_280),
.C(n_224),
.Y(n_346)
);

AO22x2_ASAP7_75t_L g347 ( 
.A1(n_304),
.A2(n_270),
.B1(n_212),
.B2(n_215),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_347),
.B(n_307),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_348),
.A2(n_357),
.B1(n_370),
.B2(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_355),
.C(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_320),
.Y(n_353)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_318),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_321),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_317),
.C(n_301),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_301),
.C(n_207),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_325),
.A2(n_336),
.B1(n_329),
.B2(n_345),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_270),
.Y(n_359)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_360),
.A2(n_215),
.B1(n_135),
.B2(n_101),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_212),
.Y(n_363)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_345),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_364),
.B(n_368),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_365),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_328),
.B(n_332),
.Y(n_367)
);

XOR2x2_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_347),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_322),
.B(n_335),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_335),
.A2(n_212),
.B1(n_168),
.B2(n_188),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_207),
.C(n_159),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_151),
.C(n_205),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_372),
.B(n_347),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_362),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_382),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_360),
.A2(n_330),
.B(n_344),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_381),
.B(n_351),
.Y(n_407)
);

XOR2x2_ASAP7_75t_SL g379 ( 
.A(n_348),
.B(n_337),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_386),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_380),
.A2(n_385),
.B1(n_391),
.B2(n_351),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_349),
.A2(n_331),
.B(n_338),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_353),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_219),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_331),
.B1(n_346),
.B2(n_347),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_347),
.Y(n_387)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_352),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_367),
.A2(n_188),
.B1(n_168),
.B2(n_215),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_393),
.A2(n_370),
.B1(n_365),
.B2(n_369),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_359),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_358),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_355),
.C(n_350),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_395),
.B(n_398),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_354),
.C(n_356),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_366),
.C(n_378),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_399),
.B(n_400),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_366),
.C(n_388),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_413),
.Y(n_426)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_402),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_372),
.C(n_371),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_403),
.B(n_410),
.Y(n_427)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_368),
.CI(n_352),
.CON(n_404),
.SN(n_404)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_385),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_407),
.A2(n_389),
.B(n_383),
.Y(n_422)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_408),
.Y(n_428)
);

OAI221xp5_ASAP7_75t_L g410 ( 
.A1(n_377),
.A2(n_361),
.B1(n_363),
.B2(n_219),
.C(n_205),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_412),
.Y(n_414)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_396),
.A2(n_390),
.B(n_387),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_422),
.B(n_423),
.Y(n_434)
);

OAI21x1_ASAP7_75t_SL g438 ( 
.A1(n_418),
.A2(n_429),
.B(n_118),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_386),
.C(n_380),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_420),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_389),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_399),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_421),
.B(n_397),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_383),
.C(n_391),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_377),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_400),
.C(n_401),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_432),
.Y(n_447)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_397),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_437),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_435),
.B(n_436),
.Y(n_454)
);

OAI221xp5_ASAP7_75t_L g436 ( 
.A1(n_428),
.A2(n_404),
.B1(n_413),
.B2(n_393),
.C(n_201),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_192),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_438),
.A2(n_36),
.B(n_25),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_424),
.A2(n_122),
.B(n_111),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_439),
.A2(n_425),
.B(n_132),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_120),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_442),
.Y(n_453)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_444),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_84),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_109),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_455),
.Y(n_462)
);

OAI21x1_ASAP7_75t_SL g446 ( 
.A1(n_434),
.A2(n_429),
.B(n_415),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_449),
.B(n_450),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_431),
.A2(n_422),
.B(n_416),
.Y(n_449)
);

AOI21xp33_ASAP7_75t_L g450 ( 
.A1(n_443),
.A2(n_430),
.B(n_3),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_444),
.A2(n_433),
.B(n_442),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_452),
.B(n_437),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_457),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_2),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_458),
.B(n_459),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_2),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_450),
.B(n_3),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_460),
.A2(n_461),
.B(n_463),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_3),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_453),
.C(n_36),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_456),
.A2(n_36),
.B(n_25),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_466),
.A2(n_462),
.B(n_4),
.Y(n_469)
);

A2O1A1O1Ixp25_ASAP7_75t_L g468 ( 
.A1(n_461),
.A2(n_25),
.B(n_36),
.C(n_5),
.D(n_6),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_468),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_470),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_465),
.A2(n_36),
.B(n_7),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

O2A1O1Ixp33_ASAP7_75t_SL g474 ( 
.A1(n_473),
.A2(n_467),
.B(n_464),
.C(n_9),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_474),
.B(n_5),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_475),
.A2(n_472),
.B1(n_5),
.B2(n_8),
.Y(n_476)
);


endmodule