module fake_jpeg_9592_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

OR2x2_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_19),
.B1(n_23),
.B2(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_58),
.B(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_34),
.B1(n_20),
.B2(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_30),
.B(n_31),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_18),
.B(n_31),
.C(n_21),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_81),
.Y(n_101)
);

NAND2x1_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_45),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_89),
.B(n_16),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_89),
.B1(n_97),
.B2(n_81),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_41),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_30),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_97),
.Y(n_114)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_19),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_88),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_112),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_80),
.B1(n_75),
.B2(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_126),
.B1(n_128),
.B2(n_108),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_47),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_26),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_61),
.B1(n_53),
.B2(n_65),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_127),
.B1(n_77),
.B2(n_96),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_46),
.C(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_62),
.C(n_44),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_110),
.Y(n_132)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_28),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_56),
.B1(n_48),
.B2(n_53),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_98),
.B1(n_90),
.B2(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_60),
.B1(n_45),
.B2(n_67),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_72),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_132),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_134),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_118),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_95),
.B1(n_93),
.B2(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_141),
.B1(n_148),
.B2(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_108),
.B1(n_126),
.B2(n_114),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_95),
.B1(n_84),
.B2(n_57),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_156),
.C(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_155),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_23),
.B(n_32),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_149),
.B(n_152),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_45),
.B1(n_66),
.B2(n_95),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_19),
.B(n_23),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_87),
.B1(n_92),
.B2(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_44),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_149),
.B(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_26),
.B(n_28),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_87),
.B1(n_102),
.B2(n_129),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_70),
.B(n_152),
.Y(n_197)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_177),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_166),
.B(n_176),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_175),
.C(n_178),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_189),
.B(n_193),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_106),
.B1(n_122),
.B2(n_120),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_187),
.B1(n_190),
.B2(n_165),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_105),
.C(n_62),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_105),
.C(n_17),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_186),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_17),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_27),
.C(n_82),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_106),
.B1(n_118),
.B2(n_87),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_192),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_135),
.B1(n_148),
.B2(n_154),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_131),
.A2(n_21),
.B(n_24),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_201),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_196),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_184),
.B(n_193),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_130),
.B1(n_153),
.B2(n_157),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_204),
.B1(n_210),
.B2(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_171),
.B1(n_179),
.B2(n_188),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_157),
.A3(n_145),
.B1(n_160),
.B2(n_24),
.C1(n_71),
.C2(n_134),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_12),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_134),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_211),
.C(n_161),
.Y(n_244)
);

OAI22x1_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_25),
.B1(n_27),
.B2(n_102),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_121),
.B1(n_24),
.B2(n_72),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_8),
.C(n_15),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_222),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_27),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_8),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_225),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_209),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_227),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_171),
.B1(n_184),
.B2(n_161),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_234),
.A2(n_246),
.B1(n_247),
.B2(n_0),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_162),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_237),
.C(n_238),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_183),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_199),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_182),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_169),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_239),
.A2(n_15),
.B(n_12),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_200),
.B1(n_206),
.B2(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_249),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_196),
.C(n_208),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_170),
.B1(n_27),
.B2(n_72),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_262),
.Y(n_284)
);

XOR2x2_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_210),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_264),
.C(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_203),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_257),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_207),
.B1(n_216),
.B2(n_195),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_265),
.B1(n_247),
.B2(n_241),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_271),
.C(n_238),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_197),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_227),
.C(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

AOI211xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_213),
.B(n_212),
.C(n_197),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_223),
.B1(n_240),
.B2(n_228),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_219),
.B1(n_15),
.B2(n_12),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_229),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_231),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_241),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_1),
.C(n_2),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_9),
.Y(n_301)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.C(n_256),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_235),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_234),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

AO221x1_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_246),
.B1(n_260),
.B2(n_271),
.C(n_257),
.Y(n_289)
);

INVx11_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_259),
.B(n_256),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_293),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_251),
.B1(n_248),
.B2(n_255),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_295),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_11),
.C(n_10),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_9),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_2),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_279),
.C(n_284),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_302),
.B1(n_277),
.B2(n_283),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_308),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_279),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_302),
.Y(n_317)
);

BUFx4f_ASAP7_75t_SL g312 ( 
.A(n_296),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_296),
.B(n_292),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_277),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_292),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_323),
.C(n_312),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_300),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_290),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_327),
.B(n_326),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_312),
.B1(n_309),
.B2(n_5),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_325),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_316),
.B(n_315),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_332),
.C(n_4),
.Y(n_334)
);

AOI221xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_335)
);

AOI221xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_301),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule