module fake_netlist_5_1400_n_1809 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1809);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1809;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_93),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_3),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_3),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_56),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_7),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_16),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_76),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_52),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_25),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_29),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_31),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_103),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx4_ASAP7_75t_R g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_97),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_36),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_41),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_11),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_70),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_40),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_7),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_108),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_94),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_143),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_79),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_42),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_77),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_50),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_16),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_132),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_52),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_89),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_60),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_37),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_100),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_57),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_49),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_129),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_153),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_139),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_39),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_23),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_148),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_21),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_9),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_88),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_61),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_55),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_86),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_27),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_85),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_44),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_40),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_118),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_125),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_112),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_141),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_109),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_154),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_18),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_24),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_33),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_159),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_99),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_13),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_136),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_35),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_65),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_115),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_6),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_68),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_46),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_66),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_110),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_27),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_21),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_63),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_15),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_78),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_34),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_4),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_104),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_142),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_35),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_53),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_60),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_74),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_95),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_137),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_45),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_51),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_105),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_98),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_101),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_45),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_38),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_31),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_54),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_146),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_51),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_75),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_15),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_102),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_164),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_55),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_33),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_67),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_64),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_43),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_1),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_120),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_71),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_22),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_124),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_20),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_152),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_46),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_151),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_59),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_117),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_126),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_22),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_96),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_203),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_209),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_235),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_178),
.B(n_1),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_178),
.B(n_2),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_170),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_262),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_205),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_262),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_212),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_262),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_219),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_262),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_171),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_222),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_220),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_220),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_223),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_180),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_193),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_206),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_230),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_210),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_327),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_230),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_197),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_225),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_226),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_229),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_259),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_230),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_233),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_261),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_265),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_238),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_208),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_295),
.Y(n_375)
);

BUFx2_ASAP7_75t_SL g376 ( 
.A(n_206),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_195),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_241),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_246),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_248),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_240),
.B(n_5),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_249),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_221),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_234),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_250),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_242),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_247),
.B(n_5),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_287),
.B(n_8),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_252),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_253),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_254),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_255),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_240),
.B(n_8),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_260),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_263),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_272),
.B(n_10),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_264),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_270),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_178),
.B(n_11),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_279),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_269),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_199),
.B(n_12),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_280),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_288),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_273),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_337),
.B(n_235),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_345),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_328),
.A2(n_245),
.B(n_199),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_337),
.B(n_327),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_360),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_245),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_336),
.B(n_276),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_330),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_347),
.Y(n_428)
);

NAND2x1_ASAP7_75t_L g429 ( 
.A(n_339),
.B(n_188),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_399),
.B(n_276),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_177),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_369),
.B(n_230),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_331),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_334),
.A2(n_285),
.B(n_275),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_388),
.B(n_327),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_334),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

CKINVDCx6p67_ASAP7_75t_R g443 ( 
.A(n_400),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_338),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_369),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_393),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_393),
.B(n_196),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_340),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_340),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_341),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_347),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_350),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_341),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_336),
.B(n_179),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_185),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_353),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_187),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_358),
.B(n_189),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_358),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_364),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_376),
.B(n_202),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_374),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_374),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_384),
.B(n_230),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_386),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_381),
.B(n_272),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_390),
.B(n_251),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_449),
.A2(n_299),
.B1(n_282),
.B2(n_236),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_381),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_449),
.B(n_332),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_432),
.A2(n_194),
.B1(n_217),
.B2(n_174),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_446),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_454),
.B(n_335),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_346),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_440),
.B(n_348),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_440),
.B(n_352),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_355),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_446),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_434),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_453),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_454),
.B(n_365),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_366),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_453),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_454),
.B(n_367),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_424),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_447),
.B(n_370),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_450),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_419),
.B(n_373),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_456),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_416),
.A2(n_216),
.B(n_215),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_419),
.B(n_378),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g517 ( 
.A(n_459),
.B(n_387),
.C(n_390),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_454),
.B(n_379),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_456),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_424),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_424),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_426),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_478),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_436),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_455),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_432),
.A2(n_459),
.B1(n_477),
.B2(n_463),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_436),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_436),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_432),
.A2(n_333),
.B1(n_387),
.B2(n_376),
.Y(n_535)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_455),
.B(n_391),
.C(n_333),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_432),
.B(n_380),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_455),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_443),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_382),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_426),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_432),
.B(n_385),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_439),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_439),
.B(n_251),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_426),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_443),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_459),
.A2(n_302),
.B1(n_314),
.B2(n_326),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_447),
.B(n_389),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_392),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_450),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_L g557 ( 
.A1(n_478),
.A2(n_391),
.B1(n_277),
.B2(n_218),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_412),
.B(n_395),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_468),
.B(n_397),
.Y(n_559)
);

OAI22xp33_ASAP7_75t_L g560 ( 
.A1(n_429),
.A2(n_278),
.B1(n_257),
.B2(n_244),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_427),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_468),
.B(n_398),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_457),
.B(n_362),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_450),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_412),
.B(n_403),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_437),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_450),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_450),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_404),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_429),
.A2(n_283),
.B1(n_232),
.B2(n_231),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_423),
.A2(n_291),
.B1(n_168),
.B2(n_169),
.Y(n_580)
);

BUFx4f_ASAP7_75t_L g581 ( 
.A(n_450),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_434),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_437),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_463),
.B(n_375),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_412),
.B(n_204),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_437),
.Y(n_586)
);

NOR2x1p5_ASAP7_75t_L g587 ( 
.A(n_443),
.B(n_166),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_428),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_412),
.B(n_271),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_437),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

INVxp33_ASAP7_75t_L g592 ( 
.A(n_457),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_438),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_438),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_438),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_434),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_441),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_428),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_443),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_435),
.B(n_342),
.Y(n_601)
);

INVx6_ASAP7_75t_L g602 ( 
.A(n_434),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_434),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_428),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_412),
.B(n_165),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_463),
.B(n_251),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_441),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_428),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_441),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_457),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_412),
.B(n_224),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_213),
.C(n_359),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_412),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_441),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_457),
.B(n_165),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g616 ( 
.A1(n_416),
.A2(n_320),
.B(n_267),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_423),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_237),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_423),
.B(n_359),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_441),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_423),
.B(n_405),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_444),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_444),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_435),
.B(n_344),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_444),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_444),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_435),
.B(n_251),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_428),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_429),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_470),
.B(n_357),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_617),
.B(n_470),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_531),
.B(n_251),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_538),
.B(n_311),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_507),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_L g635 ( 
.A(n_495),
.B(n_464),
.C(n_214),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_617),
.B(n_470),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_482),
.A2(n_472),
.B1(n_470),
.B2(n_451),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_526),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_630),
.B(n_470),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_537),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_546),
.B(n_470),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_538),
.A2(n_464),
.B(n_422),
.C(n_475),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_227),
.C(n_211),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_482),
.A2(n_472),
.B1(n_470),
.B2(n_451),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_482),
.A2(n_472),
.B1(n_444),
.B2(n_451),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_554),
.B(n_356),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_543),
.A2(n_416),
.B(n_448),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_482),
.A2(n_472),
.B1(n_448),
.B2(n_451),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_521),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_543),
.B(n_311),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_613),
.B(n_311),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_521),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_507),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_548),
.B(n_472),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_548),
.B(n_472),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_480),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_548),
.B(n_522),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_578),
.B(n_361),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_522),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_480),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_530),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_621),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_524),
.B(n_472),
.Y(n_663)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_547),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_628),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_547),
.B(n_311),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_588),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_529),
.B(n_532),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_482),
.A2(n_368),
.B1(n_371),
.B2(n_372),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_532),
.B(n_448),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_533),
.B(n_448),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_629),
.B(n_422),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_533),
.B(n_451),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_534),
.B(n_452),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_629),
.B(n_422),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_610),
.B(n_488),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_600),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_484),
.B(n_167),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_559),
.B(n_167),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g681 ( 
.A(n_600),
.B(n_172),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_534),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_570),
.B(n_584),
.Y(n_683)
);

AOI221xp5_ASAP7_75t_L g684 ( 
.A1(n_485),
.A2(n_296),
.B1(n_200),
.B2(n_198),
.C(n_192),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_530),
.B(n_394),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_514),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_514),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_561),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_619),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_519),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_489),
.B(n_452),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_499),
.B(n_452),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_628),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_519),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_491),
.B(n_172),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_610),
.A2(n_183),
.B1(n_182),
.B2(n_186),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_608),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_502),
.B(n_452),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_621),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_506),
.B(n_452),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_486),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_518),
.B(n_474),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_542),
.B(n_474),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_486),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_585),
.B(n_474),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_549),
.B(n_258),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_487),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_589),
.B(n_474),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_549),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_562),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_539),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_619),
.B(n_592),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_492),
.B(n_175),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_558),
.B(n_474),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_541),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_601),
.A2(n_624),
.B1(n_168),
.B2(n_169),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_562),
.A2(n_479),
.B1(n_474),
.B2(n_416),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_564),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_564),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_573),
.B(n_474),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_487),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_496),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_496),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_611),
.B(n_467),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_498),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_535),
.A2(n_324),
.B1(n_274),
.B2(n_284),
.Y(n_727)
);

NOR2x1p5_ASAP7_75t_L g728 ( 
.A(n_517),
.B(n_166),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_498),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_517),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_512),
.B(n_175),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_588),
.B(n_479),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_503),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_605),
.A2(n_182),
.B1(n_183),
.B2(n_186),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_SL g735 ( 
.A(n_552),
.B(n_190),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_608),
.Y(n_736)
);

OR2x2_ASAP7_75t_SL g737 ( 
.A(n_481),
.B(n_289),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_571),
.B(n_465),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_465),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_599),
.B(n_479),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_599),
.B(n_604),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_516),
.B(n_190),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_599),
.B(n_467),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_560),
.B(n_191),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_503),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_604),
.B(n_479),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_505),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_505),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_604),
.B(n_467),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_618),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_580),
.B(n_465),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_579),
.B(n_191),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_483),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_557),
.B(n_615),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_608),
.B(n_467),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_483),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_596),
.A2(n_445),
.B(n_442),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_481),
.B(n_394),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_606),
.B(n_290),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_608),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_490),
.B(n_479),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_566),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_485),
.B(n_268),
.C(n_286),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_490),
.B(n_479),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_608),
.B(n_467),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_580),
.B(n_201),
.Y(n_766)
);

NOR2x1p5_ASAP7_75t_L g767 ( 
.A(n_587),
.B(n_173),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_490),
.B(n_511),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_511),
.B(n_467),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_493),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_561),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_561),
.B(n_467),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_566),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_493),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_511),
.B(n_467),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_612),
.B(n_624),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_536),
.B(n_405),
.C(n_401),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_551),
.B(n_556),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_494),
.A2(n_305),
.B1(n_293),
.B2(n_318),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_601),
.B(n_401),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_561),
.B(n_577),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_567),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_551),
.B(n_467),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_551),
.B(n_556),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_556),
.B(n_467),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_500),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_567),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_553),
.A2(n_323),
.B(n_313),
.C(n_298),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_561),
.B(n_410),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_577),
.B(n_410),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_576),
.B(n_410),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_568),
.B(n_201),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_576),
.B(n_410),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_500),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_576),
.B(n_410),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_528),
.B(n_469),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_577),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_574),
.Y(n_798)
);

AO22x2_ASAP7_75t_L g799 ( 
.A1(n_587),
.A2(n_297),
.B1(n_312),
.B2(n_303),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_750),
.B(n_574),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_640),
.B(n_683),
.Y(n_801)
);

AOI21x1_ASAP7_75t_L g802 ( 
.A1(n_673),
.A2(n_590),
.B(n_575),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_730),
.B(n_568),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_673),
.A2(n_596),
.B(n_581),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_726),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_676),
.A2(n_596),
.B(n_581),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_676),
.A2(n_581),
.B(n_497),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_754),
.A2(n_307),
.B(n_582),
.C(n_603),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_741),
.A2(n_582),
.B(n_497),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_667),
.A2(n_603),
.B(n_540),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_738),
.B(n_575),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_739),
.B(n_590),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_633),
.A2(n_540),
.B(n_528),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_662),
.B(n_469),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_633),
.A2(n_666),
.B(n_650),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_712),
.B(n_469),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_739),
.B(n_704),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_650),
.A2(n_568),
.B(n_577),
.Y(n_819)
);

AOI21xp33_ASAP7_75t_L g820 ( 
.A1(n_766),
.A2(n_239),
.B(n_228),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_689),
.B(n_568),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_704),
.B(n_733),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_679),
.A2(n_594),
.B(n_626),
.C(n_625),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_712),
.B(n_471),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_733),
.B(n_594),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_666),
.A2(n_703),
.B(n_702),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_677),
.A2(n_699),
.B1(n_635),
.B2(n_689),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_664),
.B(n_597),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_654),
.A2(n_598),
.B(n_597),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_665),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_659),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_677),
.A2(n_606),
.B1(n_494),
.B2(n_602),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_662),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_659),
.Y(n_835)
);

OAI21xp33_ASAP7_75t_L g836 ( 
.A1(n_684),
.A2(n_680),
.B(n_695),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_634),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_664),
.B(n_598),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_665),
.B(n_577),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_732),
.A2(n_572),
.B(n_504),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_655),
.A2(n_609),
.B(n_607),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_740),
.A2(n_572),
.B(n_508),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_657),
.A2(n_494),
.B1(n_602),
.B2(n_325),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_643),
.B(n_515),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_681),
.B(n_294),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_632),
.A2(n_609),
.B(n_626),
.C(n_625),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_660),
.B(n_614),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_746),
.A2(n_572),
.B(n_508),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_717),
.A2(n_572),
.B(n_509),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_664),
.B(n_501),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_665),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_664),
.B(n_614),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_685),
.B(n_515),
.Y(n_853)
);

INVx8_ASAP7_75t_L g854 ( 
.A(n_665),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_713),
.A2(n_620),
.B(n_623),
.C(n_622),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_664),
.B(n_709),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_698),
.A2(n_550),
.B(n_501),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_701),
.B(n_620),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_647),
.A2(n_623),
.B(n_527),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_691),
.A2(n_700),
.B(n_692),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_661),
.B(n_513),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_751),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_707),
.B(n_513),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_711),
.B(n_520),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_758),
.B(n_520),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_632),
.A2(n_602),
.B1(n_494),
.B2(n_322),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_714),
.A2(n_544),
.B(n_622),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_720),
.A2(n_544),
.B(n_527),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_693),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_780),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_693),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_771),
.A2(n_563),
.B(n_545),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_744),
.A2(n_563),
.B(n_523),
.C(n_525),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_781),
.A2(n_765),
.B(n_755),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_642),
.A2(n_591),
.B(n_523),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_641),
.A2(n_639),
.B(n_636),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_705),
.A2(n_565),
.B(n_550),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_723),
.B(n_525),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_747),
.B(n_545),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_708),
.A2(n_591),
.B(n_565),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_752),
.A2(n_569),
.B(n_583),
.C(n_586),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_653),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_638),
.B(n_569),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_631),
.A2(n_583),
.B(n_595),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_797),
.A2(n_595),
.B(n_586),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_638),
.B(n_593),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_646),
.B(n_471),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_715),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_748),
.B(n_593),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_693),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_706),
.A2(n_606),
.B(n_627),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_653),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_728),
.B(n_473),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_693),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_709),
.B(n_606),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_763),
.B(n_776),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_710),
.B(n_606),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_697),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_710),
.B(n_606),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_718),
.B(n_719),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_797),
.A2(n_616),
.B(n_433),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_721),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_737),
.B(n_735),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_718),
.B(n_606),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_686),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_688),
.A2(n_616),
.B(n_442),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_L g907 ( 
.A1(n_731),
.A2(n_192),
.B(n_200),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_722),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_719),
.B(n_627),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_697),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_649),
.A2(n_602),
.B1(n_627),
.B2(n_294),
.Y(n_911)
);

CKINVDCx16_ASAP7_75t_R g912 ( 
.A(n_669),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_668),
.A2(n_325),
.B1(n_308),
.B2(n_315),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_652),
.Y(n_914)
);

NOR2x2_ASAP7_75t_L g915 ( 
.A(n_716),
.B(n_173),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_688),
.A2(n_442),
.B(n_445),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_688),
.A2(n_445),
.B(n_433),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_670),
.A2(n_627),
.B1(n_322),
.B2(n_316),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_688),
.A2(n_433),
.B(n_417),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_696),
.B(n_243),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_715),
.B(n_473),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_682),
.B(n_473),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_742),
.B(n_475),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_722),
.B(n_627),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_688),
.A2(n_420),
.B(n_425),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_706),
.A2(n_420),
.B(n_425),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_725),
.B(n_627),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_761),
.A2(n_420),
.B(n_425),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_725),
.B(n_627),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_796),
.B(n_308),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_663),
.A2(n_420),
.B(n_410),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_729),
.B(n_466),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_745),
.B(n_466),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_745),
.B(n_466),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_764),
.A2(n_417),
.B(n_420),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_767),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_781),
.A2(n_417),
.B(n_420),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_686),
.B(n_466),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_768),
.A2(n_417),
.B(n_420),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_777),
.B(n_476),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_734),
.B(n_256),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_778),
.A2(n_784),
.B(n_736),
.Y(n_942)
);

BUFx8_ASAP7_75t_L g943 ( 
.A(n_687),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_796),
.A2(n_316),
.B1(n_315),
.B2(n_466),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_796),
.B(n_476),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_687),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_690),
.B(n_266),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_690),
.B(n_176),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_637),
.B(n_410),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_645),
.A2(n_417),
.B(n_425),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_694),
.B(n_792),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_697),
.A2(n_417),
.B(n_425),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_727),
.B(n_475),
.C(n_476),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_697),
.A2(n_417),
.B(n_425),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_648),
.A2(n_425),
.B(n_406),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_SL g956 ( 
.A(n_678),
.B(n_176),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_694),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_762),
.B(n_406),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_736),
.A2(n_406),
.B(n_408),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_644),
.A2(n_408),
.B(n_414),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_678),
.B(n_181),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_736),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_736),
.A2(n_418),
.B(n_408),
.Y(n_963)
);

NOR2x2_ASAP7_75t_L g964 ( 
.A(n_799),
.B(n_181),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_773),
.B(n_413),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_760),
.A2(n_421),
.B(n_413),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_760),
.B(n_462),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_799),
.B(n_184),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_788),
.B(n_184),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_760),
.A2(n_421),
.B(n_413),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_782),
.B(n_414),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_760),
.B(n_414),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_788),
.B(n_458),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_799),
.B(n_198),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_753),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_671),
.A2(n_415),
.B(n_418),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_672),
.A2(n_415),
.B1(n_418),
.B2(n_421),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_798),
.B(n_415),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_759),
.B(n_674),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_787),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_675),
.A2(n_461),
.B(n_460),
.C(n_458),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_801),
.B(n_756),
.Y(n_982)
);

NAND2x2_ASAP7_75t_L g983 ( 
.A(n_936),
.B(n_291),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_816),
.A2(n_743),
.B(n_749),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_887),
.B(n_292),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_912),
.B(n_759),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_854),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_801),
.A2(n_651),
.B1(n_743),
.B2(n_749),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_836),
.B(n_651),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_827),
.A2(n_755),
.B(n_765),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_914),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_923),
.B(n_770),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_SL g993 ( 
.A1(n_903),
.A2(n_296),
.B1(n_300),
.B2(n_304),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_854),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_837),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_862),
.B(n_870),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_805),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_901),
.A2(n_724),
.B(n_783),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_882),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_892),
.Y(n_1000)
);

INVx6_ASAP7_75t_L g1001 ( 
.A(n_943),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_962),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_SL g1003 ( 
.A(n_941),
.B(n_300),
.C(n_304),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_820),
.A2(n_779),
.B(n_790),
.C(n_789),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_834),
.B(n_770),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_860),
.A2(n_795),
.B(n_793),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_888),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_905),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_920),
.A2(n_791),
.B(n_790),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_910),
.A2(n_769),
.B(n_785),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_SL g1011 ( 
.A1(n_809),
.A2(n_772),
.B(n_789),
.C(n_775),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_896),
.B(n_306),
.C(n_309),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_910),
.A2(n_772),
.B(n_757),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_SL g1015 ( 
.A1(n_903),
.A2(n_319),
.B1(n_309),
.B2(n_310),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_SL g1016 ( 
.A(n_896),
.B(n_306),
.C(n_310),
.Y(n_1016)
);

INVxp33_ASAP7_75t_SL g1017 ( 
.A(n_956),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_862),
.A2(n_794),
.B1(n_786),
.B2(n_774),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_941),
.A2(n_794),
.B(n_786),
.C(n_774),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_920),
.A2(n_317),
.B(n_319),
.C(n_321),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_853),
.A2(n_321),
.B(n_317),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_910),
.A2(n_814),
.B(n_951),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_SL g1023 ( 
.A1(n_803),
.A2(n_430),
.B(n_461),
.C(n_460),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_818),
.B(n_822),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_828),
.B(n_462),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_943),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_947),
.A2(n_461),
.B(n_460),
.C(n_458),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_808),
.B(n_12),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_961),
.B(n_461),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_921),
.B(n_13),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_940),
.A2(n_430),
.B1(n_460),
.B2(n_458),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_910),
.A2(n_838),
.B(n_829),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_947),
.A2(n_462),
.B(n_431),
.C(n_411),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_817),
.B(n_462),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_823),
.B(n_462),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_893),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_SL g1037 ( 
.A(n_907),
.B(n_845),
.C(n_969),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_946),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_945),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_852),
.A2(n_431),
.B(n_411),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_957),
.A2(n_462),
.B1(n_431),
.B2(n_411),
.Y(n_1041)
);

OAI22x1_ASAP7_75t_L g1042 ( 
.A1(n_968),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_930),
.A2(n_913),
.B(n_948),
.C(n_865),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_SL g1044 ( 
.A1(n_856),
.A2(n_162),
.B(n_161),
.C(n_147),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_803),
.A2(n_462),
.B(n_431),
.C(n_411),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_815),
.B(n_462),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_930),
.A2(n_14),
.B(n_17),
.C(n_20),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_957),
.A2(n_462),
.B1(n_431),
.B2(n_411),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_854),
.B(n_462),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_902),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_908),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_865),
.A2(n_431),
.B(n_411),
.C(n_407),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_802),
.A2(n_431),
.B(n_411),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_804),
.A2(n_431),
.B(n_411),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_825),
.A2(n_431),
.B1(n_411),
.B2(n_407),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_980),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_974),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_806),
.A2(n_900),
.B(n_819),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_815),
.B(n_407),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_883),
.B(n_23),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_948),
.A2(n_407),
.B(n_25),
.C(n_26),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_883),
.B(n_24),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_SL g1063 ( 
.A1(n_915),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_886),
.B(n_407),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_886),
.B(n_407),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_812),
.A2(n_407),
.B1(n_134),
.B2(n_131),
.Y(n_1066)
);

AOI22x1_ASAP7_75t_L g1067 ( 
.A1(n_807),
.A2(n_407),
.B1(n_121),
.B2(n_119),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_906),
.A2(n_407),
.B(n_113),
.Y(n_1068)
);

XNOR2xp5_ASAP7_75t_L g1069 ( 
.A(n_944),
.B(n_111),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_847),
.B(n_407),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_813),
.A2(n_106),
.B1(n_91),
.B2(n_90),
.Y(n_1071)
);

AOI33xp33_ASAP7_75t_L g1072 ( 
.A1(n_922),
.A2(n_28),
.A3(n_30),
.B1(n_32),
.B2(n_34),
.B3(n_37),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_876),
.A2(n_87),
.B(n_84),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_962),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_844),
.A2(n_32),
.B(n_38),
.C(n_41),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_847),
.A2(n_42),
.B(n_43),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_861),
.B(n_864),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_831),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_964),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_962),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_831),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_861),
.A2(n_44),
.B(n_47),
.C(n_48),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_831),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_864),
.B(n_47),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_922),
.B(n_48),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_975),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_975),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_973),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_953),
.B(n_49),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_832),
.Y(n_1090)
);

INVx3_ASAP7_75t_SL g1091 ( 
.A(n_894),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_800),
.B(n_50),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_856),
.A2(n_83),
.B(n_82),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_894),
.B(n_72),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_958),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_821),
.B(n_54),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_973),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_894),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_851),
.B(n_81),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_821),
.A2(n_61),
.B(n_841),
.C(n_830),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_826),
.B(n_835),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_894),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_L g1103 ( 
.A1(n_824),
.A2(n_875),
.B(n_855),
.C(n_976),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_965),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_851),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_942),
.A2(n_850),
.B(n_811),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_953),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_869),
.B(n_871),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_962),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_918),
.A2(n_949),
.B1(n_979),
.B2(n_843),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_932),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_979),
.A2(n_909),
.B1(n_858),
.B2(n_899),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_869),
.B(n_871),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_890),
.B(n_971),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_898),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_890),
.B(n_978),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_891),
.A2(n_928),
.B(n_935),
.C(n_846),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_977),
.A2(n_972),
.B(n_879),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_898),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_850),
.A2(n_849),
.B(n_949),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_863),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_839),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_833),
.B(n_924),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_933),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_873),
.A2(n_881),
.B(n_889),
.C(n_878),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_839),
.B(n_866),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_859),
.A2(n_810),
.B(n_929),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_950),
.B(n_874),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_1100),
.A2(n_927),
.B(n_904),
.C(n_897),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_997),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1056),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1007),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_1061),
.A2(n_895),
.B(n_967),
.C(n_981),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1118),
.A2(n_868),
.A3(n_867),
.B(n_877),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_987),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1051),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_997),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1103),
.A2(n_880),
.B(n_857),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1039),
.B(n_967),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_985),
.B(n_960),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1058),
.A2(n_872),
.B(n_885),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1050),
.Y(n_1142)
);

INVx5_ASAP7_75t_L g1143 ( 
.A(n_1083),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_991),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1077),
.B(n_938),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1036),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1039),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1095),
.B(n_934),
.Y(n_1148)
);

OAI22x1_ASAP7_75t_L g1149 ( 
.A1(n_1069),
.A2(n_972),
.B1(n_911),
.B2(n_955),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1091),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1106),
.A2(n_884),
.B(n_931),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1043),
.A2(n_939),
.B(n_926),
.C(n_842),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_987),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1054),
.A2(n_840),
.B(n_848),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_990),
.A2(n_937),
.B(n_952),
.Y(n_1155)
);

CKINVDCx8_ASAP7_75t_R g1156 ( 
.A(n_1057),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_1103),
.A2(n_970),
.B(n_966),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1090),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1090),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1001),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1088),
.A2(n_954),
.B1(n_917),
.B2(n_916),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1006),
.A2(n_959),
.B(n_963),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1120),
.A2(n_919),
.B(n_925),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_998),
.A2(n_984),
.B(n_1010),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1033),
.A2(n_1052),
.A3(n_1045),
.B(n_1117),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1001),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1112),
.A2(n_1127),
.A3(n_1019),
.B(n_989),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1022),
.A2(n_1125),
.B(n_1049),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1032),
.A2(n_992),
.B(n_1011),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_1025),
.A2(n_1110),
.B(n_1068),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1123),
.A2(n_988),
.B(n_1009),
.Y(n_1171)
);

AOI211x1_ASAP7_75t_L g1172 ( 
.A1(n_1076),
.A2(n_1104),
.B(n_1021),
.C(n_1089),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1040),
.A2(n_1005),
.B(n_1014),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1123),
.A2(n_1024),
.B(n_1126),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1024),
.A2(n_982),
.B(n_1128),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1001),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_989),
.A2(n_1027),
.A3(n_1066),
.B(n_1096),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1023),
.A2(n_1025),
.B(n_1070),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1084),
.A2(n_1062),
.B(n_1060),
.C(n_1037),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1029),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1128),
.A2(n_1064),
.B(n_1065),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1091),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_995),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1084),
.A2(n_1088),
.B1(n_1107),
.B2(n_1060),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1107),
.A2(n_1062),
.B1(n_1121),
.B2(n_1030),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1121),
.A2(n_1030),
.B1(n_1092),
.B2(n_1020),
.Y(n_1186)
);

AO32x2_ASAP7_75t_L g1187 ( 
.A1(n_1071),
.A2(n_993),
.A3(n_1015),
.B1(n_1063),
.B2(n_1048),
.Y(n_1187)
);

INVx3_ASAP7_75t_SL g1188 ( 
.A(n_1026),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_996),
.B(n_1003),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1004),
.A2(n_1073),
.B(n_1047),
.C(n_1082),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1034),
.A2(n_1005),
.B(n_1116),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_996),
.B(n_1124),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1111),
.B(n_1101),
.Y(n_1193)
);

BUFx4f_ASAP7_75t_L g1194 ( 
.A(n_1122),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_994),
.A2(n_1114),
.B(n_1074),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1085),
.B(n_1038),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_SL g1197 ( 
.A1(n_1075),
.A2(n_1094),
.B(n_1023),
.C(n_1035),
.Y(n_1197)
);

INVx3_ASAP7_75t_SL g1198 ( 
.A(n_1079),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1031),
.A2(n_1018),
.B(n_1093),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1067),
.A2(n_1035),
.B(n_1041),
.Y(n_1200)
);

AOI211xp5_ASAP7_75t_L g1201 ( 
.A1(n_1028),
.A2(n_986),
.B(n_1044),
.C(n_1017),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1109),
.A2(n_1059),
.B(n_1087),
.Y(n_1202)
);

AO32x2_ASAP7_75t_L g1203 ( 
.A1(n_1072),
.A2(n_1098),
.A3(n_1115),
.B1(n_1097),
.B2(n_1016),
.Y(n_1203)
);

BUFx2_ASAP7_75t_SL g1204 ( 
.A(n_994),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_999),
.B(n_1008),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1108),
.A2(n_1113),
.B(n_1046),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1109),
.A2(n_1086),
.B(n_1099),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1042),
.A2(n_1000),
.A3(n_1105),
.B(n_1081),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1102),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1028),
.B(n_1013),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1115),
.A2(n_1016),
.A3(n_1055),
.B(n_983),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1055),
.A2(n_983),
.A3(n_1109),
.B(n_1078),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1002),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_SL g1214 ( 
.A1(n_1013),
.A2(n_1078),
.B(n_1119),
.C(n_986),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1119),
.A2(n_1109),
.B(n_1074),
.C(n_1080),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_1002),
.A2(n_727),
.A3(n_1112),
.B1(n_988),
.B2(n_1066),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1002),
.A2(n_836),
.B1(n_1012),
.B2(n_801),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1002),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1074),
.B(n_836),
.C(n_683),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1074),
.A2(n_1103),
.B(n_1100),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1080),
.A2(n_801),
.B1(n_1077),
.B2(n_531),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1080),
.A2(n_836),
.B1(n_1012),
.B2(n_801),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_997),
.B(n_870),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_SL g1226 ( 
.A(n_1001),
.B(n_678),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1077),
.A2(n_801),
.B1(n_531),
.B2(n_862),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1043),
.A2(n_836),
.B(n_801),
.C(n_754),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1043),
.B(n_836),
.C(n_683),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1083),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1100),
.A2(n_632),
.B(n_1061),
.C(n_836),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_L g1237 ( 
.A(n_986),
.B(n_836),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_997),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1017),
.B(n_342),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1012),
.A2(n_836),
.B1(n_1076),
.B2(n_1100),
.C(n_1061),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1017),
.B(n_715),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1017),
.B(n_342),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1103),
.A2(n_1100),
.B(n_801),
.Y(n_1243)
);

NAND2x1_ASAP7_75t_L g1244 ( 
.A(n_1119),
.B(n_898),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1077),
.B(n_801),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1043),
.A2(n_836),
.B(n_801),
.C(n_754),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1083),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1077),
.B(n_801),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1118),
.A2(n_1033),
.A3(n_1052),
.B(n_1100),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1003),
.A2(n_836),
.B(n_820),
.C(n_440),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1043),
.A2(n_836),
.B(n_801),
.C(n_754),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1026),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1056),
.Y(n_1261)
);

AOI221x1_ASAP7_75t_L g1262 ( 
.A1(n_1012),
.A2(n_836),
.B1(n_1076),
.B2(n_1100),
.C(n_1061),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1001),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_997),
.Y(n_1265)
);

NAND3x1_ASAP7_75t_L g1266 ( 
.A(n_1012),
.B(n_481),
.C(n_485),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1054),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1003),
.A2(n_836),
.B(n_820),
.C(n_440),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1103),
.A2(n_1100),
.B(n_801),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1103),
.A2(n_1100),
.B(n_801),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_997),
.B(n_870),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_997),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1058),
.A2(n_816),
.B(n_827),
.Y(n_1273)
);

CKINVDCx6p67_ASAP7_75t_R g1274 ( 
.A(n_1188),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1266),
.A2(n_1237),
.B1(n_1242),
.B2(n_1239),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1130),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1245),
.A2(n_1250),
.B1(n_1189),
.B2(n_1185),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1260),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1231),
.A2(n_1184),
.B1(n_1149),
.B2(n_1185),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1131),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1231),
.A2(n_1140),
.B1(n_1184),
.B2(n_1269),
.Y(n_1281)
);

INVx8_ASAP7_75t_L g1282 ( 
.A(n_1143),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1179),
.A2(n_1228),
.B1(n_1246),
.B2(n_1259),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1261),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1186),
.A2(n_1243),
.B1(n_1270),
.B2(n_1269),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1136),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1132),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1227),
.B(n_1221),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1186),
.A2(n_1270),
.B1(n_1243),
.B2(n_1219),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1144),
.Y(n_1290)
);

INVx4_ASAP7_75t_SL g1291 ( 
.A(n_1208),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1264),
.Y(n_1292)
);

BUFx8_ASAP7_75t_SL g1293 ( 
.A(n_1194),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1219),
.A2(n_1222),
.B1(n_1217),
.B2(n_1227),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1217),
.A2(n_1222),
.B1(n_1146),
.B2(n_1241),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1171),
.A2(n_1221),
.B1(n_1139),
.B2(n_1265),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1150),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_1143),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1143),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1150),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1226),
.A2(n_1201),
.B1(n_1198),
.B2(n_1180),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1142),
.Y(n_1302)
);

CKINVDCx6p67_ASAP7_75t_R g1303 ( 
.A(n_1232),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1240),
.A2(n_1262),
.B1(n_1156),
.B2(n_1192),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1139),
.A2(n_1180),
.B1(n_1199),
.B2(n_1174),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1199),
.A2(n_1137),
.B1(n_1272),
.B2(n_1238),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1193),
.B(n_1172),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1183),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1166),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1232),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1196),
.A2(n_1210),
.B1(n_1220),
.B2(n_1147),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1225),
.A2(n_1271),
.B1(n_1194),
.B2(n_1247),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1172),
.B(n_1145),
.Y(n_1314)
);

BUFx8_ASAP7_75t_L g1315 ( 
.A(n_1160),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1176),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1209),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1182),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1232),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1247),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1247),
.A2(n_1148),
.B1(n_1159),
.B2(n_1158),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1220),
.A2(n_1187),
.B1(n_1268),
.B2(n_1255),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1135),
.Y(n_1323)
);

CKINVDCx6p67_ASAP7_75t_R g1324 ( 
.A(n_1204),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1208),
.B(n_1203),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1205),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1187),
.A2(n_1168),
.B1(n_1170),
.B2(n_1151),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1187),
.A2(n_1170),
.B1(n_1233),
.B2(n_1203),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1175),
.A2(n_1206),
.B1(n_1161),
.B2(n_1181),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1213),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1191),
.A2(n_1169),
.B1(n_1218),
.B2(n_1202),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1190),
.A2(n_1215),
.B1(n_1201),
.B2(n_1195),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1153),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1214),
.A2(n_1153),
.B1(n_1129),
.B2(n_1197),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1207),
.A2(n_1244),
.B1(n_1133),
.B2(n_1152),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1157),
.B(n_1155),
.Y(n_1336)
);

CKINVDCx6p67_ASAP7_75t_R g1337 ( 
.A(n_1211),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1178),
.A2(n_1138),
.B1(n_1273),
.B2(n_1252),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1178),
.A2(n_1138),
.B1(n_1223),
.B2(n_1229),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1208),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1212),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1234),
.A2(n_1235),
.B1(n_1249),
.B2(n_1263),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1248),
.A2(n_1256),
.B1(n_1163),
.B2(n_1164),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1212),
.Y(n_1345)
);

OAI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1200),
.A2(n_1173),
.B(n_1141),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1162),
.A2(n_1154),
.B1(n_1258),
.B2(n_1230),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1211),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1216),
.A2(n_1177),
.B1(n_1165),
.B2(n_1251),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1224),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1167),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1251),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1216),
.A2(n_1177),
.B1(n_1165),
.B2(n_1134),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1134),
.B(n_1253),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1216),
.Y(n_1355)
);

BUFx4f_ASAP7_75t_SL g1356 ( 
.A(n_1236),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1254),
.A2(n_1185),
.B1(n_440),
.B2(n_1184),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1257),
.B(n_1267),
.Y(n_1358)
);

CKINVDCx11_ASAP7_75t_R g1359 ( 
.A(n_1260),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1264),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1130),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1131),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1231),
.A2(n_836),
.B1(n_1012),
.B2(n_1003),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1131),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1131),
.Y(n_1365)
);

INVx6_ASAP7_75t_L g1366 ( 
.A(n_1264),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1266),
.A2(n_646),
.B1(n_836),
.B2(n_658),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1260),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1264),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1231),
.A2(n_836),
.B1(n_1012),
.B2(n_1003),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1231),
.A2(n_912),
.B1(n_766),
.B2(n_1063),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1260),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1266),
.A2(n_646),
.B1(n_836),
.B2(n_658),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_1150),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1260),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1131),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1130),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1150),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_1150),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1131),
.Y(n_1380)
);

BUFx2_ASAP7_75t_SL g1381 ( 
.A(n_1143),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1150),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1150),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1245),
.B(n_1250),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_1260),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1231),
.A2(n_836),
.B1(n_1012),
.B2(n_1003),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1231),
.A2(n_912),
.B1(n_766),
.B2(n_1063),
.Y(n_1387)
);

OAI22x1_ASAP7_75t_L g1388 ( 
.A1(n_1217),
.A2(n_1222),
.B1(n_1231),
.B2(n_1084),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1231),
.A2(n_836),
.B1(n_1012),
.B2(n_1003),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1131),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1231),
.A2(n_836),
.B1(n_1012),
.B2(n_1003),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1179),
.A2(n_801),
.B1(n_1250),
.B2(n_1245),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1260),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1264),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1150),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1340),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1346),
.A2(n_1354),
.B(n_1285),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1342),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1361),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1332),
.A2(n_1308),
.B(n_1334),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1291),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1361),
.Y(n_1402)
);

AO21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1289),
.A2(n_1341),
.B(n_1355),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1291),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1291),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1336),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1282),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1336),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1325),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1277),
.B(n_1392),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1359),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1282),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1322),
.B(n_1281),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1377),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1377),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1345),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1351),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1276),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1352),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1356),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1322),
.B(n_1281),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1352),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_R g1423 ( 
.A(n_1385),
.B(n_1393),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1317),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1288),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1294),
.B(n_1328),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1305),
.B(n_1296),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1327),
.B(n_1279),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1392),
.B(n_1384),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1358),
.A2(n_1343),
.B(n_1347),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1290),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1354),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1349),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1388),
.B(n_1337),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1338),
.A2(n_1339),
.B(n_1344),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1317),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1349),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1348),
.B(n_1280),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1353),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1367),
.A2(n_1373),
.B1(n_1275),
.B2(n_1301),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1353),
.B(n_1283),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1284),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1286),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1283),
.A2(n_1391),
.B(n_1363),
.Y(n_1445)
);

AO21x1_ASAP7_75t_SL g1446 ( 
.A1(n_1329),
.A2(n_1335),
.B(n_1314),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1358),
.A2(n_1343),
.B(n_1314),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1362),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1364),
.B(n_1365),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1350),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1350),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1370),
.A2(n_1386),
.B(n_1389),
.C(n_1387),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1333),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1376),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1380),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1308),
.B(n_1307),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1295),
.B(n_1312),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1390),
.B(n_1330),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1384),
.B(n_1326),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1309),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1304),
.A2(n_1332),
.B(n_1321),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1371),
.A2(n_1387),
.B1(n_1313),
.B2(n_1302),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1357),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1331),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1333),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1333),
.A2(n_1371),
.B(n_1323),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1299),
.Y(n_1467)
);

NOR2x1_ASAP7_75t_SL g1468 ( 
.A(n_1381),
.B(n_1297),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1299),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1278),
.A2(n_1375),
.B(n_1368),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1311),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1311),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1319),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1274),
.A2(n_1287),
.B1(n_1306),
.B2(n_1318),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1319),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1320),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1320),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1300),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1298),
.A2(n_1303),
.B(n_1324),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1300),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1382),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1432),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1463),
.A2(n_1395),
.B(n_1378),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1450),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1401),
.B(n_1404),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1454),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1445),
.A2(n_1383),
.B(n_1369),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1445),
.A2(n_1360),
.B1(n_1316),
.B2(n_1372),
.C(n_1310),
.Y(n_1488)
);

AOI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1452),
.A2(n_1315),
.B1(n_1374),
.B2(n_1379),
.C(n_1366),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1418),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1413),
.A2(n_1293),
.B(n_1395),
.C(n_1378),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1411),
.Y(n_1492)
);

OAI211xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1463),
.A2(n_1315),
.B(n_1374),
.C(n_1379),
.Y(n_1493)
);

AO21x1_ASAP7_75t_L g1494 ( 
.A1(n_1462),
.A2(n_1378),
.B(n_1395),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1450),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1409),
.B(n_1366),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1430),
.B(n_1394),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1441),
.B(n_1394),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1462),
.A2(n_1292),
.B1(n_1427),
.B2(n_1410),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1399),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1401),
.B(n_1292),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1430),
.B(n_1459),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1402),
.B(n_1414),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1439),
.B(n_1435),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1439),
.B(n_1435),
.Y(n_1505)
);

NOR2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1407),
.B(n_1412),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1404),
.B(n_1405),
.Y(n_1507)
);

AO32x2_ASAP7_75t_L g1508 ( 
.A1(n_1403),
.A2(n_1437),
.A3(n_1428),
.B1(n_1438),
.B2(n_1434),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1470),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1415),
.B(n_1425),
.Y(n_1510)
);

OAI211xp5_ASAP7_75t_L g1511 ( 
.A1(n_1413),
.A2(n_1421),
.B(n_1457),
.C(n_1429),
.Y(n_1511)
);

AO32x1_ASAP7_75t_L g1512 ( 
.A1(n_1421),
.A2(n_1429),
.A3(n_1426),
.B1(n_1419),
.B2(n_1422),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1449),
.Y(n_1513)
);

O2A1O1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1400),
.A2(n_1457),
.B(n_1461),
.C(n_1464),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1458),
.B(n_1466),
.Y(n_1515)
);

NAND4xp25_ASAP7_75t_L g1516 ( 
.A(n_1418),
.B(n_1456),
.C(n_1424),
.D(n_1425),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1458),
.B(n_1466),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1431),
.A2(n_1464),
.B(n_1400),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_R g1519 ( 
.A(n_1466),
.B(n_1420),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1426),
.A2(n_1461),
.B1(n_1427),
.B2(n_1442),
.C(n_1440),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1455),
.B(n_1460),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1451),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1424),
.A2(n_1427),
.B1(n_1456),
.B2(n_1437),
.Y(n_1523)
);

INVx6_ASAP7_75t_L g1524 ( 
.A(n_1478),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1461),
.A2(n_1427),
.B(n_1469),
.C(n_1477),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1461),
.A2(n_1471),
.B(n_1469),
.C(n_1477),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1440),
.B(n_1443),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1431),
.B(n_1466),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1471),
.B(n_1472),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1436),
.A2(n_1468),
.B1(n_1420),
.B2(n_1453),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1467),
.Y(n_1531)
);

AOI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1405),
.A2(n_1408),
.B(n_1406),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1417),
.B(n_1460),
.Y(n_1533)
);

AO32x2_ASAP7_75t_L g1534 ( 
.A1(n_1403),
.A2(n_1433),
.A3(n_1447),
.B1(n_1398),
.B2(n_1396),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1444),
.B(n_1448),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1515),
.B(n_1447),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1510),
.B(n_1447),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1494),
.A2(n_1446),
.B1(n_1470),
.B2(n_1436),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1499),
.A2(n_1446),
.B1(n_1470),
.B2(n_1436),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1517),
.B(n_1447),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1486),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1484),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1534),
.B(n_1397),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_SL g1545 ( 
.A(n_1509),
.B(n_1423),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1520),
.A2(n_1470),
.B1(n_1436),
.B2(n_1472),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1502),
.B(n_1482),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1483),
.Y(n_1548)
);

INVx5_ASAP7_75t_L g1549 ( 
.A(n_1528),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1535),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1498),
.A2(n_1473),
.B1(n_1476),
.B2(n_1416),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_SL g1552 ( 
.A(n_1513),
.B(n_1465),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1521),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1533),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1498),
.A2(n_1473),
.B1(n_1476),
.B2(n_1416),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1495),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_SL g1557 ( 
.A(n_1509),
.B(n_1423),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1533),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1511),
.A2(n_1453),
.B1(n_1397),
.B2(n_1468),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1533),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1544),
.Y(n_1561)
);

AOI33xp33_ASAP7_75t_L g1562 ( 
.A1(n_1559),
.A2(n_1514),
.A3(n_1525),
.B1(n_1490),
.B2(n_1489),
.B3(n_1526),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1547),
.B(n_1497),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1528),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1538),
.B(n_1527),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1538),
.B(n_1527),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1547),
.B(n_1516),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1544),
.B(n_1528),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1543),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1552),
.A2(n_1532),
.B(n_1518),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1545),
.A2(n_1523),
.B1(n_1487),
.B2(n_1488),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1559),
.A2(n_1530),
.B1(n_1528),
.B2(n_1501),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1534),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1522),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1549),
.B(n_1485),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1537),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1549),
.B(n_1507),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1552),
.Y(n_1580)
);

AOI322xp5_ASAP7_75t_L g1581 ( 
.A1(n_1545),
.A2(n_1491),
.A3(n_1505),
.B1(n_1504),
.B2(n_1474),
.C1(n_1501),
.C2(n_1508),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1536),
.B(n_1534),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1534),
.Y(n_1583)
);

AND2x2_ASAP7_75t_SL g1584 ( 
.A(n_1557),
.B(n_1483),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1541),
.B(n_1556),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1548),
.B(n_1522),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1549),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1549),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1573),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1588),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1573),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1587),
.B(n_1558),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1587),
.B(n_1558),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1576),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1567),
.B(n_1550),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1586),
.B(n_1575),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1571),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1587),
.B(n_1560),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1550),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1563),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1588),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1571),
.A2(n_1546),
.B1(n_1557),
.B2(n_1540),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1569),
.Y(n_1610)
);

OAI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1581),
.A2(n_1539),
.B(n_1555),
.C(n_1551),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1577),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1577),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1588),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1553),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1587),
.B(n_1560),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1569),
.Y(n_1619)
);

CKINVDCx16_ASAP7_75t_R g1620 ( 
.A(n_1572),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1581),
.B(n_1531),
.Y(n_1621)
);

INVx6_ASAP7_75t_L g1622 ( 
.A(n_1591),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1579),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1579),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1560),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1589),
.B(n_1590),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1593),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1592),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1581),
.B(n_1531),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1579),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1563),
.B(n_1492),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1594),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1626),
.B(n_1564),
.Y(n_1633)
);

AOI32xp33_ASAP7_75t_L g1634 ( 
.A1(n_1602),
.A2(n_1629),
.A3(n_1621),
.B1(n_1620),
.B2(n_1580),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1622),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1597),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1606),
.B(n_1562),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1631),
.B(n_1492),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1597),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1594),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1596),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1600),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1596),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1622),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1626),
.B(n_1564),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1601),
.B(n_1565),
.Y(n_1647)
);

OAI321xp33_ASAP7_75t_L g1648 ( 
.A1(n_1609),
.A2(n_1572),
.A3(n_1571),
.B1(n_1580),
.B2(n_1493),
.C(n_1565),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1627),
.B(n_1564),
.Y(n_1649)
);

AND2x4_ASAP7_75t_SL g1650 ( 
.A(n_1610),
.B(n_1576),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1603),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1598),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1627),
.B(n_1593),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1605),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1598),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1599),
.B(n_1564),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1599),
.B(n_1568),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1611),
.A2(n_1572),
.B(n_1584),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1601),
.B(n_1565),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1620),
.B(n_1591),
.C(n_1585),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1662)
);

OR2x6_ASAP7_75t_L g1663 ( 
.A(n_1622),
.B(n_1591),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1609),
.B(n_1591),
.C(n_1585),
.Y(n_1664)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1665 ( 
.A1(n_1619),
.A2(n_1491),
.B(n_1566),
.C(n_1575),
.D(n_1580),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1613),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1613),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1628),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1595),
.B(n_1585),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_1605),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1617),
.B(n_1608),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1622),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1604),
.B(n_1506),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1663),
.B(n_1622),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1668),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1641),
.B(n_1566),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1642),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1663),
.B(n_1568),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1659),
.A2(n_1584),
.B(n_1503),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1643),
.B(n_1617),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1637),
.B(n_1566),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1642),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1638),
.B(n_1500),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1648),
.A2(n_1584),
.B(n_1512),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1663),
.Y(n_1687)
);

AND2x2_ASAP7_75t_SL g1688 ( 
.A(n_1671),
.B(n_1584),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1654),
.B(n_1501),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1634),
.B(n_1589),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1664),
.A2(n_1584),
.B(n_1512),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1644),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1673),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1655),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1661),
.B(n_1593),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1663),
.B(n_1568),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1653),
.B(n_1672),
.Y(n_1697)
);

NOR3xp33_ASAP7_75t_SL g1698 ( 
.A(n_1674),
.B(n_1519),
.C(n_1529),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1672),
.B(n_1595),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1635),
.B(n_1593),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1655),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1666),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1653),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1653),
.B(n_1589),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1633),
.B(n_1625),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1647),
.B(n_1590),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1633),
.B(n_1646),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1647),
.B(n_1660),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1678),
.Y(n_1711)
);

OAI32xp33_ASAP7_75t_L g1712 ( 
.A1(n_1690),
.A2(n_1665),
.A3(n_1669),
.B1(n_1674),
.B2(n_1660),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1684),
.B(n_1635),
.Y(n_1713)
);

AOI222xp33_ASAP7_75t_L g1714 ( 
.A1(n_1688),
.A2(n_1650),
.B1(n_1583),
.B2(n_1574),
.C1(n_1582),
.C2(n_1646),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1693),
.Y(n_1715)
);

AOI32xp33_ASAP7_75t_L g1716 ( 
.A1(n_1695),
.A2(n_1650),
.A3(n_1645),
.B1(n_1657),
.B2(n_1658),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1680),
.A2(n_1669),
.B(n_1645),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1676),
.B(n_1662),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1703),
.B(n_1662),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1709),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1688),
.A2(n_1549),
.B1(n_1669),
.B2(n_1591),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1685),
.A2(n_1549),
.B1(n_1591),
.B2(n_1585),
.Y(n_1723)
);

NOR3xp33_ASAP7_75t_L g1724 ( 
.A(n_1691),
.B(n_1479),
.C(n_1591),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1687),
.A2(n_1585),
.B1(n_1593),
.B2(n_1639),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1689),
.A2(n_1585),
.B1(n_1519),
.B2(n_1578),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1697),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1675),
.B(n_1576),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1687),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1677),
.A2(n_1570),
.B(n_1666),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1683),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1682),
.A2(n_1576),
.B1(n_1578),
.B2(n_1656),
.Y(n_1732)
);

NAND5xp2_ASAP7_75t_SL g1733 ( 
.A(n_1675),
.B(n_1658),
.C(n_1657),
.D(n_1582),
.E(n_1574),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1710),
.B(n_1608),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1698),
.A2(n_1640),
.B(n_1632),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1681),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1729),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1711),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1736),
.B(n_1681),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1715),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1727),
.B(n_1709),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1720),
.A2(n_1705),
.B1(n_1696),
.B2(n_1679),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1719),
.A2(n_1713),
.B1(n_1724),
.B2(n_1728),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1700),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1721),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1731),
.Y(n_1746)
);

OAI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1717),
.A2(n_1699),
.B1(n_1696),
.B2(n_1679),
.C(n_1692),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1718),
.B(n_1704),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1716),
.A2(n_1724),
.B(n_1735),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1734),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1722),
.A2(n_1700),
.B1(n_1704),
.B2(n_1706),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1714),
.B(n_1706),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1712),
.A2(n_1683),
.B(n_1694),
.C(n_1702),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1733),
.A2(n_1700),
.B1(n_1699),
.B2(n_1707),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1732),
.B(n_1707),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1740),
.B(n_1726),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1737),
.Y(n_1758)
);

XNOR2xp5_ASAP7_75t_L g1759 ( 
.A(n_1743),
.B(n_1723),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1749),
.A2(n_1730),
.B(n_1686),
.C(n_1702),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1749),
.A2(n_1730),
.B1(n_1701),
.B2(n_1694),
.C(n_1686),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1753),
.B(n_1701),
.C(n_1479),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1750),
.B(n_1708),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1739),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1755),
.A2(n_1639),
.B1(n_1636),
.B2(n_1656),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1744),
.B(n_1636),
.Y(n_1766)
);

AOI322xp5_ASAP7_75t_L g1767 ( 
.A1(n_1752),
.A2(n_1583),
.A3(n_1574),
.B1(n_1582),
.B2(n_1652),
.C1(n_1561),
.C2(n_1590),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1758),
.Y(n_1768)
);

NOR4xp25_ASAP7_75t_L g1769 ( 
.A(n_1764),
.B(n_1760),
.C(n_1761),
.D(n_1757),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1766),
.Y(n_1770)
);

NOR3xp33_ASAP7_75t_L g1771 ( 
.A(n_1763),
.B(n_1747),
.C(n_1741),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1759),
.A2(n_1751),
.B(n_1748),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1762),
.B(n_1742),
.C(n_1738),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1765),
.A2(n_1744),
.B1(n_1756),
.B2(n_1754),
.Y(n_1774)
);

NOR2x1_ASAP7_75t_L g1775 ( 
.A(n_1767),
.B(n_1745),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1759),
.B(n_1746),
.Y(n_1776)
);

INVxp33_ASAP7_75t_SL g1777 ( 
.A(n_1764),
.Y(n_1777)
);

NAND4xp25_ASAP7_75t_SL g1778 ( 
.A(n_1775),
.B(n_1652),
.C(n_1667),
.D(n_1670),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1772),
.A2(n_1651),
.B(n_1475),
.C(n_1607),
.Y(n_1779)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1780 ( 
.A1(n_1769),
.A2(n_1630),
.B(n_1615),
.C(n_1623),
.D(n_1614),
.Y(n_1780)
);

NAND4xp75_ASAP7_75t_L g1781 ( 
.A(n_1768),
.B(n_1607),
.C(n_1595),
.D(n_1616),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1776),
.A2(n_1529),
.B1(n_1616),
.B2(n_1607),
.C(n_1583),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1778),
.B(n_1773),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1782),
.A2(n_1771),
.B1(n_1777),
.B2(n_1774),
.C(n_1770),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1779),
.A2(n_1616),
.B1(n_1582),
.B2(n_1583),
.C(n_1574),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1780),
.Y(n_1786)
);

NOR3xp33_ASAP7_75t_L g1787 ( 
.A(n_1781),
.B(n_1475),
.C(n_1467),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1780),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1783),
.B(n_1612),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1788),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1784),
.A2(n_1576),
.B1(n_1578),
.B2(n_1496),
.Y(n_1791)
);

NOR2xp67_ASAP7_75t_L g1792 ( 
.A(n_1787),
.B(n_1475),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1786),
.A2(n_1576),
.B1(n_1578),
.B2(n_1496),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1790),
.B(n_1785),
.C(n_1467),
.Y(n_1794)
);

O2A1O1Ixp33_ASAP7_75t_L g1795 ( 
.A1(n_1789),
.A2(n_1475),
.B(n_1592),
.C(n_1630),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1792),
.A2(n_1624),
.B(n_1623),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1794),
.Y(n_1797)
);

OAI22x1_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1791),
.B1(n_1793),
.B2(n_1795),
.Y(n_1798)
);

AO211x2_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1796),
.B(n_1624),
.C(n_1615),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1798),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1800),
.Y(n_1801)
);

AOI22x1_ASAP7_75t_L g1802 ( 
.A1(n_1799),
.A2(n_1480),
.B1(n_1531),
.B2(n_1453),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1801),
.A2(n_1407),
.B1(n_1412),
.B2(n_1524),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1802),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1804),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1805),
.B(n_1803),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1806),
.Y(n_1807)
);

OAI221xp5_ASAP7_75t_R g1808 ( 
.A1(n_1807),
.A2(n_1407),
.B1(n_1412),
.B2(n_1612),
.C(n_1478),
.Y(n_1808)
);

AOI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1808),
.A2(n_1480),
.B(n_1531),
.C(n_1481),
.Y(n_1809)
);


endmodule