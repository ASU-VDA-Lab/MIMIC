module real_jpeg_6488_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_0),
.B(n_213),
.Y(n_212)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_2),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_2),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_66),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_2),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_2),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_3),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_3),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_206),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_4),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_5),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_5),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_6),
.B(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_13),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_14),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_15),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_15),
.B(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_160),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_158),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_19),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_72),
.B2(n_138),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_42),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.C(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_23),
.A2(n_24),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_25),
.B(n_27),
.Y(n_157)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_26),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g153 ( 
.A(n_29),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_145)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_35),
.Y(n_149)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_51),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_54),
.B(n_132),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_54),
.B(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_115),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_91),
.C(n_106),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_74),
.B(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_87),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_82),
.C(n_87),
.Y(n_137)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_84),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_106),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_93),
.B1(n_101),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_97),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_102),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_102),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_114),
.Y(n_135)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_133),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_128),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_124),
.B2(n_127),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_146),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_140),
.A2(n_141),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_143),
.B(n_146),
.Y(n_244)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.C(n_157),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_157),
.Y(n_165)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_240),
.B(n_245),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_200),
.B(n_239),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_181),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_163),
.B(n_181),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_164),
.B(n_167),
.C(n_178),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_178),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_176),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_183),
.Y(n_182)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_198),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_185),
.B1(n_198),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_194),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_187),
.B1(n_194),
.B2(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_233),
.B(n_238),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_219),
.B(n_232),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_207),
.C(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_226),
.B(n_231),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_230),
.Y(n_231)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);


endmodule