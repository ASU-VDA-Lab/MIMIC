module real_jpeg_12644_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_238, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_238;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_57),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_20),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_4),
.A2(n_29),
.B1(n_54),
.B2(n_58),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_4),
.A2(n_29),
.B1(n_51),
.B2(n_52),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_37),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_37),
.B1(n_54),
.B2(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_7),
.B(n_64),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_7),
.B(n_21),
.C(n_41),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_7),
.B(n_96),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_7),
.B(n_42),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_7),
.A2(n_52),
.B(n_66),
.C(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_7),
.B(n_48),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_10),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_99)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

XNOR2x2_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_128),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_126),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_101),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_15),
.B(n_101),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_74),
.C(n_91),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_16),
.B(n_91),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_45),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_17),
.B(n_63),
.C(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_30),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_18),
.B(n_30),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_24),
.B(n_26),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_19),
.A2(n_25),
.B(n_90),
.Y(n_89)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_20),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_21),
.B(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_28),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_24),
.A2(n_25),
.B(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_24),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_24),
.B(n_95),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_25),
.B(n_138),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_27),
.B(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_27),
.B(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_43),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_31),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_32),
.B(n_42),
.Y(n_189)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_33),
.A2(n_98),
.B(n_123),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_34),
.A2(n_37),
.B(n_67),
.Y(n_182)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_35),
.B(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_49),
.C(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_38),
.B(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_38),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_42),
.B(n_143),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_43),
.A2(n_99),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_43),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_59),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_47),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_48),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_58),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_60),
.Y(n_77)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B(n_71),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_64),
.B(n_83),
.Y(n_178)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_68),
.B(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_69),
.B(n_115),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_74),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.C(n_84),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_75),
.B(n_78),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_81),
.B(n_114),
.Y(n_197)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_84),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_206)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_153),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_125),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_118),
.B2(n_119),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_111),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_120),
.A2(n_121),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI321xp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_221),
.A3(n_230),
.B1(n_235),
.B2(n_236),
.C(n_238),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_201),
.B(n_220),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_185),
.B(n_200),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_173),
.B(n_184),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_154),
.B(n_172),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_148),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_148),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_147),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.C(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_166),
.B(n_171),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_162),
.B(n_165),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_169),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_179),
.C(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_199),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_199),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_193),
.B1(n_194),
.B2(n_198),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_191),
.C(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_206),
.C(n_207),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.CI(n_197),
.CON(n_194),
.SN(n_194)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_215),
.C(n_218),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);


endmodule