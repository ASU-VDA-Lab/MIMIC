module fake_jpeg_11449_n_550 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_550);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_62),
.Y(n_119)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_96),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_27),
.Y(n_77)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_0),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_89),
.Y(n_136)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_103),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_132),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_48),
.B1(n_36),
.B2(n_21),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_107),
.A2(n_144),
.B1(n_28),
.B2(n_30),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_58),
.A2(n_50),
.B1(n_43),
.B2(n_42),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_109),
.A2(n_124),
.B1(n_73),
.B2(n_70),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_20),
.B1(n_29),
.B2(n_35),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_114),
.A2(n_167),
.B1(n_121),
.B2(n_46),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_20),
.B1(n_29),
.B2(n_35),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_115),
.A2(n_122),
.B1(n_46),
.B2(n_40),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_66),
.A2(n_29),
.B1(n_35),
.B2(n_43),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_85),
.A2(n_43),
.B1(n_50),
.B2(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_63),
.B(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_19),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_30),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_137),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_72),
.A2(n_26),
.B1(n_50),
.B2(n_42),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_26),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_60),
.A2(n_43),
.B1(n_50),
.B2(n_46),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_169),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_105),
.B(n_97),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_170),
.Y(n_261)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_124),
.A2(n_74),
.B1(n_101),
.B2(n_100),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_174),
.A2(n_180),
.B1(n_193),
.B2(n_215),
.Y(n_253)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_192),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_179),
.B(n_181),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_95),
.B1(n_90),
.B2(n_98),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_28),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_28),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_182),
.B(n_190),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_185),
.A2(n_196),
.B1(n_201),
.B2(n_120),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_186),
.Y(n_282)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_187),
.Y(n_252)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_51),
.Y(n_190)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_152),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_51),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_116),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_51),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_203),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_209),
.Y(n_279)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_213),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_211),
.Y(n_281)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_216),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_99),
.B1(n_41),
.B2(n_40),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_150),
.B(n_41),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_227),
.B1(n_151),
.B2(n_166),
.Y(n_246)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_220),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_138),
.A2(n_155),
.B1(n_129),
.B2(n_143),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_219),
.A2(n_226),
.B1(n_31),
.B2(n_32),
.Y(n_273)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_138),
.A2(n_40),
.B1(n_30),
.B2(n_41),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_222),
.A2(n_119),
.B1(n_121),
.B2(n_155),
.Y(n_229)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_224),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_225),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_129),
.A2(n_76),
.B1(n_52),
.B2(n_96),
.Y(n_226)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_76),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_228),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_229),
.A2(n_237),
.B1(n_269),
.B2(n_272),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_153),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_245),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_174),
.A2(n_136),
.B1(n_166),
.B2(n_151),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_240),
.A2(n_227),
.B1(n_210),
.B2(n_218),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_162),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_161),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_168),
.B(n_118),
.C(n_160),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_250),
.C(n_260),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_160),
.Y(n_250)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_173),
.B(n_126),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_260),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_196),
.B(n_52),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_262),
.B(n_212),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_185),
.A2(n_125),
.B1(n_31),
.B2(n_32),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_180),
.A2(n_125),
.B1(n_31),
.B2(n_102),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_175),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_222),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_178),
.B(n_0),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_191),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_184),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g290 ( 
.A(n_280),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_202),
.B(n_223),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_283),
.A2(n_291),
.B(n_308),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_284),
.Y(n_372)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_287),
.B(n_297),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_253),
.B(n_242),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_236),
.B(n_211),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_293),
.B(n_299),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_189),
.C(n_177),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_309),
.C(n_324),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_229),
.A2(n_215),
.B1(n_226),
.B2(n_207),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_295),
.A2(n_322),
.B1(n_268),
.B2(n_255),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_248),
.B(n_220),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_329),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_301),
.A2(n_310),
.B1(n_318),
.B2(n_325),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_169),
.B1(n_208),
.B2(n_183),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_312),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_231),
.B(n_205),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_304),
.B(n_328),
.Y(n_369)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_307),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_253),
.A2(n_242),
.B(n_233),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_245),
.B(n_264),
.C(n_232),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_261),
.A2(n_217),
.B1(n_198),
.B2(n_186),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_314),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_315),
.B(n_316),
.Y(n_344)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_234),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_269),
.A2(n_224),
.B(n_188),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_265),
.B(n_243),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_235),
.A2(n_32),
.B1(n_3),
.B2(n_4),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_251),
.A2(n_2),
.B(n_3),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_320),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_275),
.A2(n_4),
.B(n_5),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_321),
.B(n_241),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_280),
.A2(n_32),
.B1(n_6),
.B2(n_7),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_323),
.A2(n_328),
.B1(n_330),
.B2(n_267),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_249),
.B(n_8),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_273),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_260),
.A2(n_14),
.B(n_9),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_260),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_277),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_233),
.A2(n_11),
.B(n_12),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_267),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_263),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_331),
.A2(n_268),
.B1(n_239),
.B2(n_257),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_278),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_257),
.C(n_270),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_342),
.B(n_366),
.C(n_287),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_347),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_258),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_345),
.B(n_362),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_346),
.A2(n_358),
.B1(n_325),
.B2(n_303),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_258),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_243),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_355),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_290),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_356),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_292),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_291),
.A2(n_255),
.B1(n_282),
.B2(n_239),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_307),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_360),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_288),
.B(n_243),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_361),
.B(n_317),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_270),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_364),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_285),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_307),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_365),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_296),
.B(n_241),
.C(n_230),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_316),
.B(n_321),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_367),
.B(n_368),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_288),
.B(n_308),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_369),
.B(n_370),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_259),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_317),
.A2(n_259),
.B1(n_266),
.B2(n_238),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_371),
.A2(n_357),
.B1(n_360),
.B2(n_340),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_312),
.B(n_266),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_373),
.B(n_326),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_339),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_376),
.B(n_380),
.Y(n_428)
);

XOR2x2_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_324),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_339),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_298),
.B(n_283),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_SL g435 ( 
.A1(n_385),
.A2(n_410),
.B(n_386),
.C(n_400),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_363),
.A2(n_313),
.B1(n_298),
.B2(n_326),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_386),
.A2(n_395),
.B1(n_346),
.B2(n_337),
.Y(n_415)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_391),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g392 ( 
.A1(n_368),
.A2(n_313),
.A3(n_311),
.B1(n_294),
.B2(n_315),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_314),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_396),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_356),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_402),
.C(n_378),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_334),
.B(n_297),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_353),
.A2(n_327),
.B(n_320),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_403),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_355),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_406),
.B(n_407),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_351),
.B(n_286),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_408),
.A2(n_409),
.B1(n_357),
.B2(n_371),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_358),
.A2(n_318),
.B1(n_300),
.B2(n_284),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_349),
.A2(n_329),
.B(n_274),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_336),
.C(n_342),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_400),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_384),
.A2(n_373),
.B1(n_354),
.B2(n_372),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_412),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_435),
.B1(n_376),
.B2(n_380),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_422),
.C(n_431),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_415),
.A2(n_423),
.B1(n_426),
.B2(n_429),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_336),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_434),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_388),
.B(n_333),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_421),
.B(n_430),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_366),
.C(n_361),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_395),
.A2(n_346),
.B1(n_343),
.B2(n_353),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_401),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_442),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_377),
.A2(n_346),
.B1(n_337),
.B2(n_374),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_337),
.B1(n_374),
.B2(n_369),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_381),
.B(n_333),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_350),
.C(n_332),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_332),
.C(n_335),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_397),
.C(n_405),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_338),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_383),
.B1(n_379),
.B2(n_390),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_440),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_396),
.Y(n_437)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_375),
.C(n_404),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_387),
.A2(n_393),
.B1(n_406),
.B2(n_389),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_401),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_438),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_444),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_438),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_458),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_392),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_452),
.Y(n_471)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_375),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_453),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_454),
.A2(n_408),
.B1(n_435),
.B2(n_409),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_455),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_428),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_460),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_382),
.Y(n_458)
);

XOR2x2_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_461),
.Y(n_481)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_417),
.Y(n_462)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_394),
.Y(n_463)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_463),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_391),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_466),
.C(n_467),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_407),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_364),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_405),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_403),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_432),
.C(n_416),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_448),
.A2(n_433),
.B1(n_423),
.B2(n_415),
.Y(n_475)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_482),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_434),
.C(n_427),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_480),
.C(n_483),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_452),
.C(n_445),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_457),
.A2(n_447),
.B(n_433),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_426),
.C(n_435),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_451),
.A2(n_413),
.B1(n_418),
.B2(n_424),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_486),
.B1(n_490),
.B2(n_244),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_451),
.A2(n_404),
.B1(n_435),
.B2(n_429),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_465),
.B1(n_463),
.B2(n_467),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_447),
.A2(n_397),
.B1(n_338),
.B2(n_385),
.Y(n_490)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_468),
.Y(n_492)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_492),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_487),
.B(n_464),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_497),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_486),
.A2(n_454),
.B(n_457),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_494),
.A2(n_482),
.B(n_483),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_495),
.A2(n_496),
.B1(n_490),
.B2(n_481),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_489),
.A2(n_449),
.B1(n_466),
.B2(n_469),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_476),
.B(n_446),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_410),
.C(n_460),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_507),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_458),
.Y(n_499)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_472),
.B(n_323),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_502),
.C(n_509),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_335),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_485),
.A2(n_372),
.B1(n_244),
.B2(n_238),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_506),
.Y(n_521)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_508),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_256),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_519),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_480),
.C(n_479),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_517),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_478),
.C(n_477),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_518),
.A2(n_501),
.B1(n_521),
.B2(n_514),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_504),
.A2(n_484),
.B(n_474),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_503),
.A2(n_471),
.B(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_520),
.B(n_522),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_503),
.C(n_471),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_525),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_511),
.B(n_495),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_526),
.A2(n_506),
.B1(n_510),
.B2(n_519),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_494),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_528),
.B(n_530),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_502),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_470),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_532),
.B(n_533),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_523),
.B(n_499),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_522),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_535),
.A2(n_538),
.B(n_529),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_515),
.C(n_521),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_539),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_541),
.A2(n_542),
.B(n_534),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_536),
.A2(n_529),
.B1(n_510),
.B2(n_533),
.Y(n_542)
);

OAI221xp5_ASAP7_75t_L g543 ( 
.A1(n_534),
.A2(n_496),
.B1(n_500),
.B2(n_230),
.C(n_274),
.Y(n_543)
);

OAI211xp5_ASAP7_75t_SL g545 ( 
.A1(n_543),
.A2(n_274),
.B(n_537),
.C(n_256),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_544),
.A2(n_545),
.B(n_540),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_274),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_547),
.A2(n_12),
.B(n_13),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_13),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_549),
.B(n_14),
.Y(n_550)
);


endmodule