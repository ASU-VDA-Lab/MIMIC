module fake_jpeg_0_n_353 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_75),
.Y(n_80)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_54),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_14),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_11),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_73),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_28),
.A2(n_13),
.B(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_0),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_10),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_23),
.B(n_37),
.C(n_31),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_67),
.B(n_16),
.C(n_24),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_37),
.B1(n_26),
.B2(n_31),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_87),
.A2(n_114),
.B1(n_115),
.B2(n_1),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_97),
.B(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_20),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_20),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_34),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_105),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_25),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_111),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_51),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_18),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_127),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_18),
.B(n_33),
.C(n_25),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_109),
.A2(n_96),
.B(n_125),
.C(n_124),
.D(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_33),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_26),
.B1(n_35),
.B2(n_41),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_63),
.A2(n_35),
.B1(n_41),
.B2(n_40),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_41),
.C(n_24),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_115),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_68),
.A2(n_24),
.B1(n_16),
.B2(n_36),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_40),
.B1(n_36),
.B2(n_4),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_10),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_85),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_129),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_162),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_93),
.B(n_124),
.C(n_110),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_61),
.B1(n_72),
.B2(n_36),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_144),
.B1(n_154),
.B2(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_149),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_80),
.A2(n_40),
.B1(n_36),
.B2(n_4),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_40),
.B1(n_3),
.B2(n_5),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_161),
.B1(n_92),
.B2(n_118),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_90),
.B(n_94),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_1),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_165),
.B1(n_166),
.B2(n_170),
.Y(n_204)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_154)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_82),
.B(n_6),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_150),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_84),
.A2(n_6),
.B1(n_7),
.B2(n_88),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_83),
.A2(n_89),
.B1(n_104),
.B2(n_120),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_119),
.B(n_89),
.C(n_96),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_113),
.B1(n_86),
.B2(n_126),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_113),
.B1(n_86),
.B2(n_126),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_92),
.A2(n_104),
.B1(n_120),
.B2(n_95),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_84),
.A2(n_96),
.B1(n_118),
.B2(n_125),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_174),
.B1(n_165),
.B2(n_131),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_92),
.B1(n_95),
.B2(n_117),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_179),
.A2(n_155),
.B(n_200),
.C(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_93),
.C(n_117),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_192),
.C(n_195),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_100),
.A3(n_112),
.B1(n_116),
.B2(n_139),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_200),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_100),
.B(n_170),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_134),
.B(n_149),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_207),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_163),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_157),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_134),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_194),
.B(n_205),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_204),
.A2(n_140),
.B1(n_142),
.B2(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_217),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_213),
.A2(n_214),
.B1(n_220),
.B2(n_238),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_137),
.B1(n_166),
.B2(n_144),
.Y(n_214)
);

AO22x2_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_145),
.B1(n_167),
.B2(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_185),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_129),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_231),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_225),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_169),
.B1(n_143),
.B2(n_133),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_143),
.B1(n_132),
.B2(n_128),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_224),
.Y(n_241)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx10_ASAP7_75t_R g244 ( 
.A(n_222),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_233),
.B(n_177),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_155),
.A3(n_184),
.B1(n_179),
.B2(n_180),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_178),
.Y(n_225)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_237),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_196),
.C(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_172),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_190),
.B(n_189),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_186),
.A2(n_171),
.B1(n_174),
.B2(n_190),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_176),
.CI(n_197),
.CON(n_240),
.SN(n_240)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_240),
.B(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_176),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.Y(n_266)
);

AND2x6_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_189),
.Y(n_245)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_248),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_194),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_255),
.B(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_209),
.A2(n_182),
.B1(n_238),
.B2(n_213),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_262),
.B1(n_239),
.B2(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_182),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_260),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_231),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_208),
.C(n_227),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_223),
.B1(n_212),
.B2(n_221),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_223),
.B(n_233),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_271),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_241),
.A2(n_216),
.B(n_214),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_244),
.Y(n_297)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_216),
.B1(n_236),
.B2(n_234),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_211),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_278),
.C(n_284),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_216),
.B(n_237),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_261),
.B1(n_250),
.B2(n_247),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_239),
.A2(n_227),
.B(n_226),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_244),
.B(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_234),
.C(n_222),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_240),
.C(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_253),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_240),
.C(n_255),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_269),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_287),
.B(n_302),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_274),
.B1(n_277),
.B2(n_272),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_250),
.B1(n_242),
.B2(n_248),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_291),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_245),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_300),
.C(n_301),
.Y(n_306)
);

NAND4xp25_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.C(n_266),
.D(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_273),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_285),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_303),
.A2(n_312),
.B1(n_309),
.B2(n_314),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_266),
.B1(n_268),
.B2(n_275),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_267),
.C(n_282),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_293),
.C(n_300),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_299),
.B(n_292),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_307),
.C(n_305),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_301),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_306),
.B(n_287),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_326),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_323),
.A2(n_316),
.B1(n_299),
.B2(n_315),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_286),
.C(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_303),
.Y(n_333)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_328),
.B(n_330),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_280),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_323),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_332),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_308),
.B(n_312),
.C(n_275),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_319),
.B(n_333),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_321),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_340),
.B(n_341),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_321),
.B1(n_280),
.B2(n_335),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

AOI322xp5_ASAP7_75t_L g344 ( 
.A1(n_339),
.A2(n_304),
.A3(n_324),
.B1(n_335),
.B2(n_326),
.C1(n_318),
.C2(n_265),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_344),
.Y(n_347)
);

AOI21x1_ASAP7_75t_L g348 ( 
.A1(n_345),
.A2(n_346),
.B(n_341),
.Y(n_348)
);

NOR4xp25_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_317),
.C(n_307),
.D(n_265),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_343),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_349),
.B(n_347),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_304),
.B(n_270),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_270),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_270),
.Y(n_353)
);


endmodule