module fake_ariane_2945_n_4773 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_913, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_1008, n_581, n_294, n_1020, n_646, n_197, n_640, n_463, n_1024, n_830, n_176, n_691, n_34, n_404, n_172, n_943, n_678, n_651, n_987, n_936, n_347, n_423, n_961, n_183, n_469, n_479, n_726, n_603, n_878, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_908, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_1029, n_985, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_906, n_416, n_969, n_283, n_919, n_50, n_187, n_525, n_806, n_367, n_970, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_924, n_927, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_864, n_952, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_940, n_346, n_1016, n_214, n_764, n_979, n_348, n_552, n_2, n_462, n_607, n_670, n_897, n_32, n_949, n_956, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_891, n_737, n_137, n_885, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_917, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_960, n_520, n_980, n_870, n_87, n_714, n_279, n_905, n_702, n_945, n_958, n_207, n_790, n_857, n_898, n_363, n_720, n_968, n_354, n_41, n_813, n_926, n_140, n_725, n_419, n_151, n_28, n_146, n_1009, n_230, n_270, n_194, n_633, n_900, n_154, n_883, n_338, n_142, n_995, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_871, n_315, n_903, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_879, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_1018, n_855, n_158, n_69, n_259, n_835, n_95, n_808, n_953, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_1003, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_858, n_242, n_645, n_989, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_928, n_3, n_271, n_465, n_486, n_507, n_901, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_971, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_894, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_868, n_326, n_681, n_778, n_227, n_48, n_874, n_188, n_323, n_550, n_1023, n_988, n_635, n_707, n_997, n_330, n_914, n_400, n_689, n_694, n_884, n_11, n_129, n_126, n_983, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_1015, n_536, n_644, n_293, n_823, n_921, n_620, n_228, n_325, n_276, n_93, n_688, n_859, n_636, n_427, n_108, n_587, n_497, n_693, n_863, n_303, n_671, n_442, n_777, n_929, n_168, n_81, n_1, n_206, n_352, n_538, n_899, n_920, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_1013, n_986, n_638, n_136, n_334, n_192, n_729, n_887, n_661, n_488, n_775, n_667, n_300, n_533, n_904, n_505, n_14, n_163, n_88, n_869, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_957, n_977, n_512, n_715, n_889, n_935, n_579, n_844, n_1012, n_459, n_685, n_221, n_321, n_911, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_861, n_175, n_950, n_1017, n_711, n_877, n_1021, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_942, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_907, n_235, n_1006, n_881, n_660, n_464, n_735, n_575, n_546, n_1019, n_297, n_962, n_662, n_641, n_1005, n_503, n_941, n_700, n_910, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_939, n_371, n_845, n_888, n_199, n_918, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_865, n_10, n_414, n_571, n_680, n_287, n_302, n_993, n_380, n_6, n_948, n_582, n_94, n_284, n_922, n_1004, n_4, n_448, n_593, n_755, n_710, n_860, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_255, n_560, n_450, n_890, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_1022, n_135, n_896, n_409, n_171, n_947, n_930, n_519, n_902, n_384, n_468, n_853, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_872, n_933, n_13, n_27, n_916, n_254, n_596, n_954, n_912, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_982, n_915, n_215, n_252, n_629, n_664, n_161, n_454, n_966, n_992, n_298, n_955, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_984, n_537, n_223, n_403, n_25, n_750, n_834, n_991, n_83, n_389, n_1007, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_951, n_1026, n_213, n_938, n_862, n_110, n_304, n_895, n_659, n_67, n_509, n_583, n_1014, n_724, n_306, n_666, n_1000, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_946, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_875, n_669, n_785, n_827, n_931, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_967, n_998, n_999, n_472, n_937, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_880, n_793, n_852, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_1027, n_996, n_521, n_963, n_873, n_51, n_496, n_739, n_1028, n_76, n_342, n_866, n_26, n_246, n_517, n_925, n_530, n_0, n_792, n_1001, n_824, n_428, n_159, n_1002, n_358, n_105, n_580, n_892, n_608, n_959, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_975, n_563, n_229, n_394, n_923, n_250, n_932, n_773, n_165, n_144, n_981, n_1010, n_882, n_990, n_317, n_867, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_944, n_749, n_994, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_973, n_523, n_268, n_972, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_856, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_876, n_618, n_411, n_484, n_712, n_849, n_909, n_976, n_353, n_22, n_736, n_767, n_1025, n_241, n_29, n_357, n_412, n_687, n_447, n_964, n_191, n_382, n_797, n_489, n_80, n_480, n_978, n_211, n_642, n_1011, n_97, n_408, n_828, n_595, n_322, n_251, n_974, n_506, n_893, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_854, n_471, n_351, n_886, n_965, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_934, n_783, n_675, n_4773);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_913;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_1008;
input n_581;
input n_294;
input n_1020;
input n_646;
input n_197;
input n_640;
input n_463;
input n_1024;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_943;
input n_678;
input n_651;
input n_987;
input n_936;
input n_347;
input n_423;
input n_961;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_878;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_908;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_1029;
input n_985;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_906;
input n_416;
input n_969;
input n_283;
input n_919;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_970;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_924;
input n_927;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_864;
input n_952;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_940;
input n_346;
input n_1016;
input n_214;
input n_764;
input n_979;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_897;
input n_32;
input n_949;
input n_956;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_891;
input n_737;
input n_137;
input n_885;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_917;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_960;
input n_520;
input n_980;
input n_870;
input n_87;
input n_714;
input n_279;
input n_905;
input n_702;
input n_945;
input n_958;
input n_207;
input n_790;
input n_857;
input n_898;
input n_363;
input n_720;
input n_968;
input n_354;
input n_41;
input n_813;
input n_926;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_1009;
input n_230;
input n_270;
input n_194;
input n_633;
input n_900;
input n_154;
input n_883;
input n_338;
input n_142;
input n_995;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_871;
input n_315;
input n_903;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_879;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_1018;
input n_855;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_953;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_1003;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_858;
input n_242;
input n_645;
input n_989;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_928;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_901;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_971;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_894;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_868;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_874;
input n_188;
input n_323;
input n_550;
input n_1023;
input n_988;
input n_635;
input n_707;
input n_997;
input n_330;
input n_914;
input n_400;
input n_689;
input n_694;
input n_884;
input n_11;
input n_129;
input n_126;
input n_983;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_1015;
input n_536;
input n_644;
input n_293;
input n_823;
input n_921;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_859;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_863;
input n_303;
input n_671;
input n_442;
input n_777;
input n_929;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_899;
input n_920;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_1013;
input n_986;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_887;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_904;
input n_505;
input n_14;
input n_163;
input n_88;
input n_869;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_957;
input n_977;
input n_512;
input n_715;
input n_889;
input n_935;
input n_579;
input n_844;
input n_1012;
input n_459;
input n_685;
input n_221;
input n_321;
input n_911;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_861;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_877;
input n_1021;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_942;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_907;
input n_235;
input n_1006;
input n_881;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_1019;
input n_297;
input n_962;
input n_662;
input n_641;
input n_1005;
input n_503;
input n_941;
input n_700;
input n_910;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_939;
input n_371;
input n_845;
input n_888;
input n_199;
input n_918;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_865;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_993;
input n_380;
input n_6;
input n_948;
input n_582;
input n_94;
input n_284;
input n_922;
input n_1004;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_860;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_255;
input n_560;
input n_450;
input n_890;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_1022;
input n_135;
input n_896;
input n_409;
input n_171;
input n_947;
input n_930;
input n_519;
input n_902;
input n_384;
input n_468;
input n_853;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_872;
input n_933;
input n_13;
input n_27;
input n_916;
input n_254;
input n_596;
input n_954;
input n_912;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_982;
input n_915;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_966;
input n_992;
input n_298;
input n_955;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_984;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_991;
input n_83;
input n_389;
input n_1007;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_951;
input n_1026;
input n_213;
input n_938;
input n_862;
input n_110;
input n_304;
input n_895;
input n_659;
input n_67;
input n_509;
input n_583;
input n_1014;
input n_724;
input n_306;
input n_666;
input n_1000;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_875;
input n_669;
input n_785;
input n_827;
input n_931;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_967;
input n_998;
input n_999;
input n_472;
input n_937;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_880;
input n_793;
input n_852;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_1027;
input n_996;
input n_521;
input n_963;
input n_873;
input n_51;
input n_496;
input n_739;
input n_1028;
input n_76;
input n_342;
input n_866;
input n_26;
input n_246;
input n_517;
input n_925;
input n_530;
input n_0;
input n_792;
input n_1001;
input n_824;
input n_428;
input n_159;
input n_1002;
input n_358;
input n_105;
input n_580;
input n_892;
input n_608;
input n_959;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_975;
input n_563;
input n_229;
input n_394;
input n_923;
input n_250;
input n_932;
input n_773;
input n_165;
input n_144;
input n_981;
input n_1010;
input n_882;
input n_990;
input n_317;
input n_867;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_944;
input n_749;
input n_994;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_973;
input n_523;
input n_268;
input n_972;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_856;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_876;
input n_618;
input n_411;
input n_484;
input n_712;
input n_849;
input n_909;
input n_976;
input n_353;
input n_22;
input n_736;
input n_767;
input n_1025;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_964;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_978;
input n_211;
input n_642;
input n_1011;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_974;
input n_506;
input n_893;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_854;
input n_471;
input n_351;
input n_886;
input n_965;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_934;
input n_783;
input n_675;

output n_4773;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4688;
wire n_3432;
wire n_2163;
wire n_1681;
wire n_4030;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_4770;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_4586;
wire n_1469;
wire n_4342;
wire n_4692;
wire n_4557;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_4475;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_4403;
wire n_4602;
wire n_1713;
wire n_2818;
wire n_1436;
wire n_2407;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_4626;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_1837;
wire n_4178;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4547;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_4058;
wire n_2006;
wire n_4090;
wire n_2446;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_2461;
wire n_2207;
wire n_2702;
wire n_1706;
wire n_3719;
wire n_4363;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_2238;
wire n_2529;
wire n_1503;
wire n_4103;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_4683;
wire n_1298;
wire n_2653;
wire n_2873;
wire n_1745;
wire n_4610;
wire n_1366;
wire n_4674;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_4416;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4439;
wire n_2547;
wire n_4600;
wire n_3382;
wire n_1453;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_4575;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_4660;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4653;
wire n_4106;
wire n_4589;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_4581;
wire n_2960;
wire n_4260;
wire n_4625;
wire n_3270;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_4148;
wire n_1062;
wire n_3679;
wire n_4702;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_1736;
wire n_4512;
wire n_2342;
wire n_4590;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_4038;
wire n_4132;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_4500;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_4734;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_4722;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_4515;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_2878;
wire n_1284;
wire n_1428;
wire n_1241;
wire n_3890;
wire n_4741;
wire n_3830;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_2782;
wire n_3879;
wire n_4136;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_4567;
wire n_4176;
wire n_1207;
wire n_4760;
wire n_4124;
wire n_3606;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_3474;
wire n_2232;
wire n_4488;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_3552;
wire n_1542;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3324;
wire n_3209;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_4608;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_4597;
wire n_4560;
wire n_3482;
wire n_1900;
wire n_3948;
wire n_4621;
wire n_1074;
wire n_3230;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_4546;
wire n_1889;
wire n_1977;
wire n_4768;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4454;
wire n_4147;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_2332;
wire n_1703;
wire n_3975;
wire n_3828;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_3571;
wire n_2004;
wire n_3183;
wire n_3883;
wire n_1850;
wire n_4032;
wire n_4018;
wire n_4576;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_4117;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_2341;
wire n_1654;
wire n_2899;
wire n_1560;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_4572;
wire n_4505;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1230;
wire n_2739;
wire n_3739;
wire n_1840;
wire n_3962;
wire n_1597;
wire n_4082;
wire n_4476;
wire n_2942;
wire n_4680;
wire n_1771;
wire n_2902;
wire n_4541;
wire n_4360;
wire n_1544;
wire n_3271;
wire n_4540;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_1267;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_2956;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_4443;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_4665;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_4593;
wire n_4562;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_2909;
wire n_1121;
wire n_1416;
wire n_1378;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_4747;
wire n_1830;
wire n_3850;
wire n_4529;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_4498;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_2969;
wire n_1669;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_4432;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_4495;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_4737;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_2806;
wire n_1935;
wire n_4109;
wire n_3191;
wire n_1716;
wire n_4108;
wire n_3777;
wire n_4530;
wire n_4502;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_4740;
wire n_3588;
wire n_1108;
wire n_1590;
wire n_3280;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3900;
wire n_4115;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_2134;
wire n_3862;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_4513;
wire n_1179;
wire n_4311;
wire n_3284;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_2791;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_4378;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_4459;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_2855;
wire n_1182;
wire n_2166;
wire n_2848;
wire n_4594;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_4709;
wire n_1562;
wire n_3306;
wire n_2748;
wire n_2185;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4642;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_1972;
wire n_1178;
wire n_2015;
wire n_2925;
wire n_1292;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_4718;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_4130;
wire n_1083;
wire n_3937;
wire n_2161;
wire n_1418;
wire n_4763;
wire n_4175;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_4587;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_4456;
wire n_1312;
wire n_4508;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_3651;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_2365;
wire n_1880;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_3559;
wire n_3792;
wire n_1903;
wire n_1623;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_2224;
wire n_1226;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_4410;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_3567;
wire n_4003;
wire n_1392;
wire n_2795;
wire n_1832;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_4438;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_3884;
wire n_4492;
wire n_1147;
wire n_2829;
wire n_4367;
wire n_4433;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_4445;
wire n_3673;
wire n_1563;
wire n_3052;
wire n_4254;
wire n_4462;
wire n_2507;
wire n_4219;
wire n_4484;
wire n_3438;
wire n_4723;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_4451;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1234;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_2681;
wire n_1363;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_2632;
wire n_1255;
wire n_3179;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_4613;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_2980;
wire n_1095;
wire n_3699;
wire n_3078;
wire n_1728;
wire n_2335;
wire n_3971;
wire n_4315;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_4442;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_4494;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_4207;
wire n_3711;
wire n_4201;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_4725;
wire n_2312;
wire n_2677;
wire n_4296;
wire n_3171;
wire n_1826;
wire n_4719;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_4751;
wire n_3994;
wire n_4636;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_2996;
wire n_3660;
wire n_2812;
wire n_1496;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_4049;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_3589;
wire n_1869;
wire n_3623;
wire n_1743;
wire n_4522;
wire n_2718;
wire n_4263;
wire n_4707;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_4426;
wire n_3876;
wire n_4588;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2178;
wire n_1802;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_4634;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_4658;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4089;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_4699;
wire n_1198;
wire n_4096;
wire n_4506;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_4728;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_4138;
wire n_4643;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_2476;
wire n_1365;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_4713;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_2122;
wire n_3572;
wire n_1611;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_4543;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_4555;
wire n_1901;
wire n_2055;
wire n_4486;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_3118;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4441;
wire n_1906;
wire n_4323;
wire n_1899;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_4447;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_4640;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_4458;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_4523;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3983;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3286;
wire n_4480;
wire n_3734;
wire n_3370;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_4583;
wire n_3788;
wire n_3939;
wire n_2075;
wire n_3542;
wire n_1726;
wire n_3263;
wire n_3569;
wire n_3837;
wire n_2523;
wire n_1945;
wire n_3835;
wire n_2418;
wire n_2496;
wire n_1614;
wire n_1162;
wire n_1377;
wire n_2031;
wire n_3260;
wire n_3761;
wire n_3349;
wire n_3819;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_1602;
wire n_4348;
wire n_4616;
wire n_4771;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_3403;
wire n_4261;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_4661;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_2254;
wire n_3290;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_1402;
wire n_1242;
wire n_3957;
wire n_2774;
wire n_2707;
wire n_2754;
wire n_4580;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_3995;
wire n_1119;
wire n_4460;
wire n_3713;
wire n_4670;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_4648;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_4481;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4461;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_2660;
wire n_1859;
wire n_3426;
wire n_1502;
wire n_4615;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_3737;
wire n_3931;
wire n_2516;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_2949;
wire n_2661;
wire n_1294;
wire n_2894;
wire n_2300;
wire n_1667;
wire n_3896;
wire n_4067;
wire n_2452;
wire n_1649;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_4551;
wire n_3214;
wire n_3551;
wire n_4521;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_4677;
wire n_1844;
wire n_4525;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_4387;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_3186;
wire n_1791;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_2594;
wire n_1460;
wire n_1239;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_4324;
wire n_3626;
wire n_1898;
wire n_4428;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_4598;
wire n_4729;
wire n_4464;
wire n_4463;
wire n_1793;
wire n_4446;
wire n_3180;
wire n_3648;
wire n_4662;
wire n_3423;
wire n_1081;
wire n_1975;
wire n_1373;
wire n_1388;
wire n_2119;
wire n_1266;
wire n_1540;
wire n_2742;
wire n_1719;
wire n_3671;
wire n_4396;
wire n_4440;
wire n_2366;
wire n_1797;
wire n_2493;
wire n_4425;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_4565;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_1800;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_4652;
wire n_3016;
wire n_4114;
wire n_2460;
wire n_4552;
wire n_2840;
wire n_1580;
wire n_3135;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_4482;
wire n_2480;
wire n_3024;
wire n_4528;
wire n_2772;
wire n_3564;
wire n_1700;
wire n_2637;
wire n_3795;
wire n_1332;
wire n_2306;
wire n_4328;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4568;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2916;
wire n_1394;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4351;
wire n_4424;
wire n_3340;
wire n_4429;
wire n_4192;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_2581;
wire n_1527;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_4524;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_4646;
wire n_4657;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_4436;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_3836;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_4545;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_2489;
wire n_1161;
wire n_4758;
wire n_3685;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_2492;
wire n_3864;
wire n_4694;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_1215;
wire n_4664;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_2265;
wire n_4633;
wire n_4708;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_4050;
wire n_3173;
wire n_3732;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_1804;
wire n_1406;
wire n_4717;
wire n_4306;
wire n_4739;
wire n_3174;
wire n_2684;
wire n_1405;
wire n_3314;
wire n_2726;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_4671;
wire n_2272;
wire n_3266;
wire n_4766;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_4558;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4511;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_4675;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_4289;
wire n_1137;
wire n_1873;
wire n_1856;
wire n_1258;
wire n_1476;
wire n_2723;
wire n_2016;
wire n_2725;
wire n_2667;
wire n_1524;
wire n_3925;
wire n_2928;
wire n_4651;
wire n_4689;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_3167;
wire n_2850;
wire n_3746;
wire n_1293;
wire n_1874;
wire n_4748;
wire n_4537;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_4618;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_2307;
wire n_1488;
wire n_1330;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_4704;
wire n_3129;
wire n_2720;
wire n_1561;
wire n_1556;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_2064;
wire n_2353;
wire n_1429;
wire n_1324;
wire n_2528;
wire n_3543;
wire n_3640;
wire n_1778;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_1154;
wire n_4330;
wire n_1557;
wire n_1759;
wire n_2325;
wire n_1829;
wire n_1130;
wire n_4635;
wire n_4724;
wire n_1450;
wire n_4152;
wire n_4744;
wire n_3718;
wire n_4706;
wire n_2022;
wire n_3390;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_4666;
wire n_4764;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_2546;
wire n_2890;
wire n_2454;
wire n_2911;
wire n_3455;
wire n_3381;
wire n_1493;
wire n_3736;
wire n_4466;
wire n_3313;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_2760;
wire n_3907;
wire n_1864;
wire n_4603;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_4419;
wire n_1151;
wire n_4595;
wire n_4420;
wire n_4703;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3605;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_4721;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4404;
wire n_4742;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_4630;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_4377;
wire n_4617;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_4563;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4732;
wire n_4301;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_4727;
wire n_1303;
wire n_4561;
wire n_1547;
wire n_1438;
wire n_3291;
wire n_1541;
wire n_4188;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_4641;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_2610;
wire n_3715;
wire n_1593;
wire n_4140;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_4712;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_3982;
wire n_4715;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_2665;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_4755;
wire n_2771;
wire n_3755;
wire n_1090;
wire n_2403;
wire n_3842;
wire n_2947;
wire n_1367;
wire n_4202;
wire n_4536;
wire n_2044;
wire n_4534;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_3769;
wire n_4078;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_4437;
wire n_1192;
wire n_3738;
wire n_3098;
wire n_1380;
wire n_4503;
wire n_1624;
wire n_3055;
wire n_2854;
wire n_1801;
wire n_1291;
wire n_4070;
wire n_2020;
wire n_3987;
wire n_2310;
wire n_4249;
wire n_4418;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_3386;
wire n_4139;
wire n_4769;
wire n_4582;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_2177;
wire n_3695;
wire n_1511;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_4450;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_4412;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4368;
wire n_3444;
wire n_4370;
wire n_4682;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_4091;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_2343;
wire n_1048;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_4184;
wire n_4430;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_4631;
wire n_1356;
wire n_2234;
wire n_3189;
wire n_2309;
wire n_1341;
wire n_3233;
wire n_1955;
wire n_1504;
wire n_2431;
wire n_2110;
wire n_3289;
wire n_3175;
wire n_1440;
wire n_1773;
wire n_2666;
wire n_3322;
wire n_4544;
wire n_4538;
wire n_1370;
wire n_1603;
wire n_4191;
wire n_4478;
wire n_4409;
wire n_2935;
wire n_2401;
wire n_4246;
wire n_3822;
wire n_4355;
wire n_3255;
wire n_3818;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_4061;
wire n_2658;
wire n_3587;
wire n_3509;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_4601;
wire n_3344;
wire n_4754;
wire n_1403;
wire n_1065;
wire n_1948;
wire n_3006;
wire n_1534;
wire n_2767;
wire n_4518;
wire n_4155;
wire n_3376;
wire n_4278;
wire n_4531;
wire n_4710;
wire n_1959;
wire n_1290;
wire n_3497;
wire n_3770;
wire n_4375;
wire n_4542;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_4532;
wire n_4685;
wire n_2692;
wire n_3927;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_4684;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_2645;
wire n_2553;
wire n_1420;
wire n_3790;
wire n_4711;
wire n_2749;
wire n_2592;
wire n_1454;
wire n_3490;
wire n_2459;
wire n_4413;
wire n_3396;
wire n_1210;
wire n_4241;
wire n_2751;
wire n_1135;
wire n_2566;
wire n_3113;
wire n_1622;
wire n_4183;
wire n_3101;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_3251;
wire n_3288;
wire n_1885;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3904;
wire n_3887;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_4650;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_3409;
wire n_1653;
wire n_1749;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_4469;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_4455;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_4384;
wire n_1157;
wire n_1584;
wire n_4366;
wire n_4639;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_4733;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_1814;
wire n_4210;
wire n_4577;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_4623;
wire n_2315;
wire n_1857;
wire n_3926;
wire n_4209;
wire n_1687;
wire n_4457;
wire n_2073;
wire n_2150;
wire n_4509;
wire n_4004;
wire n_1552;
wire n_2938;
wire n_3630;
wire n_2498;
wire n_1612;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_3106;
wire n_2977;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_4669;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_3786;
wire n_2455;
wire n_3092;
wire n_2600;
wire n_1617;
wire n_3437;
wire n_2231;
wire n_4270;
wire n_2828;
wire n_4212;
wire n_4620;
wire n_1626;
wire n_3436;
wire n_4584;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_4759;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_1175;
wire n_2299;
wire n_3751;
wire n_4388;
wire n_3402;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_4477;
wire n_1621;
wire n_4110;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_1221;
wire n_4217;
wire n_4585;
wire n_1785;
wire n_1262;
wire n_4271;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_4687;
wire n_2974;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1183;
wire n_3722;
wire n_3686;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_4605;
wire n_4720;
wire n_3301;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_2503;
wire n_1758;
wire n_3873;
wire n_4649;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_2465;
wire n_1407;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_2428;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_3178;
wire n_2858;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_3100;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_4592;
wire n_1176;
wire n_3721;
wire n_3676;
wire n_3677;
wire n_2010;
wire n_1564;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4644;
wire n_4086;
wire n_4752;
wire n_1482;
wire n_2356;
wire n_1361;
wire n_4746;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_1520;
wire n_2534;
wire n_4656;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_4672;
wire n_3536;
wire n_2564;
wire n_1721;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_1445;
wire n_3034;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_4435;
wire n_4053;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_4750;
wire n_3177;
wire n_4667;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_3091;
wire n_4496;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_4596;
wire n_4673;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_4628;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_2639;
wire n_3855;
wire n_1775;
wire n_1036;
wire n_4738;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_4554;
wire n_2630;
wire n_4105;
wire n_4526;
wire n_2794;
wire n_3663;
wire n_2028;
wire n_3114;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_3225;
wire n_2086;
wire n_1625;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_4578;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_2409;
wire n_1720;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_3360;
wire n_4470;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_2787;
wire n_1809;
wire n_4092;
wire n_3585;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_4659;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_4057;
wire n_2770;
wire n_4550;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4647;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_3042;
wire n_1067;
wire n_4144;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_2012;
wire n_1937;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_4726;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_2212;
wire n_3838;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_4434;
wire n_2835;
wire n_1452;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_4499;
wire n_2569;
wire n_4504;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_4339;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_4497;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_4510;
wire n_3155;
wire n_4300;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4472;
wire n_4253;
wire n_1710;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_1865;
wire n_2463;
wire n_3546;
wire n_2699;
wire n_2355;
wire n_2580;
wire n_1390;
wire n_1344;
wire n_1792;
wire n_4064;
wire n_3351;
wire n_2062;
wire n_4489;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_2153;
wire n_2324;
wire n_1459;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_4519;
wire n_1099;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_3693;
wire n_1575;
wire n_3878;
wire n_4197;
wire n_4564;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_4681;
wire n_3778;
wire n_4654;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_4566;
wire n_3970;
wire n_4371;
wire n_2351;
wire n_1619;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_1902;
wire n_2206;
wire n_2784;
wire n_4414;
wire n_3898;
wire n_2541;
wire n_1643;
wire n_4185;
wire n_3188;
wire n_3232;
wire n_3001;
wire n_1320;
wire n_4448;
wire n_1113;
wire n_4749;
wire n_3218;
wire n_2347;
wire n_4676;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_1733;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_2538;
wire n_1845;
wire n_4295;
wire n_3932;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_4579;
wire n_4507;
wire n_2104;
wire n_4756;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_2552;
wire n_1533;
wire n_1576;
wire n_3445;
wire n_1470;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_4473;
wire n_4619;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_4471;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_4238;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_4691;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_4397;
wire n_4449;
wire n_3285;
wire n_3824;
wire n_4607;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_4753;
wire n_1150;
wire n_4266;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_4373;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_4407;
wire n_2472;
wire n_4695;
wire n_2705;
wire n_2664;
wire n_4165;
wire n_4154;
wire n_4479;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_4668;
wire n_2519;
wire n_3637;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_3941;
wire n_1915;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_2240;
wire n_4168;
wire n_1369;
wire n_4258;
wire n_2846;
wire n_4298;
wire n_4743;
wire n_3371;
wire n_1781;
wire n_4571;
wire n_3137;
wire n_2917;
wire n_4250;
wire n_2544;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_4415;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_2188;
wire n_1777;
wire n_1477;
wire n_1982;
wire n_2097;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_2297;
wire n_3094;
wire n_1410;
wire n_4276;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4700;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_4679;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_4408;
wire n_1983;
wire n_2982;
wire n_1273;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_4767;
wire n_2913;
wire n_4569;
wire n_1862;
wire n_2017;
wire n_3752;
wire n_4483;
wire n_3672;
wire n_3061;
wire n_1810;
wire n_2587;
wire n_3504;
wire n_2839;
wire n_1347;
wire n_4693;
wire n_3237;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_4036;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_4487;
wire n_4548;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_4539;
wire n_4574;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_4698;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_3071;
wire n_3918;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_4501;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_1946;
wire n_2148;
wire n_3244;
wire n_4383;
wire n_3499;
wire n_4391;
wire n_3112;
wire n_2562;
wire n_2051;
wire n_1779;
wire n_1168;
wire n_1821;
wire n_4095;
wire n_4444;
wire n_4663;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_4485;
wire n_4624;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_4678;
wire n_2585;
wire n_3293;
wire n_3361;
wire n_2995;
wire n_1591;
wire n_4533;
wire n_4287;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_2381;
wire n_1732;
wire n_4686;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_3779;
wire n_1705;
wire n_3707;
wire n_3895;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_4627;
wire n_4761;
wire n_3149;
wire n_1063;
wire n_3934;
wire n_4556;
wire n_2205;
wire n_2275;
wire n_2183;
wire n_4338;
wire n_2563;
wire n_3088;
wire n_1724;
wire n_4224;
wire n_4606;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_4573;
wire n_1891;
wire n_4520;
wire n_1328;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_3058;
wire n_2047;
wire n_4072;
wire n_2792;
wire n_1818;
wire n_1146;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_4465;
wire n_4553;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_3557;
wire n_1598;
wire n_3592;
wire n_3725;
wire n_1699;
wire n_3986;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3894;
wire n_4772;
wire n_4612;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1368;
wire n_1211;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_2891;
wire n_1725;
wire n_4335;
wire n_2318;
wire n_3128;
wire n_1827;
wire n_4120;
wire n_4149;
wire n_2361;
wire n_2880;
wire n_2819;
wire n_3030;
wire n_1115;
wire n_2229;
wire n_3075;
wire n_1722;
wire n_1752;
wire n_1313;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_4614;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_4629;
wire n_2551;
wire n_1102;
wire n_4516;
wire n_2255;
wire n_1252;
wire n_2239;
wire n_1129;
wire n_3045;
wire n_4716;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_4730;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_4599;
wire n_2830;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4622;
wire n_4222;
wire n_2514;
wire n_1871;
wire n_4757;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_3201;
wire n_3334;
wire n_1569;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_3162;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_4591;
wire n_4046;
wire n_4467;
wire n_4701;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_4570;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_4696;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_4655;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_2689;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_4493;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_4645;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_2479;
wire n_3204;
wire n_1981;
wire n_1069;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_2345;
wire n_4417;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_339),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_922),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_340),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_208),
.Y(n_1033)
);

CKINVDCx16_ASAP7_75t_R g1034 ( 
.A(n_797),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_793),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_336),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_251),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_698),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_350),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_344),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_455),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_342),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_791),
.Y(n_1043)
);

CKINVDCx16_ASAP7_75t_R g1044 ( 
.A(n_213),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_103),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_1010),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_158),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_433),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_241),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_684),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_844),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_985),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_981),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_915),
.Y(n_1054)
);

CKINVDCx16_ASAP7_75t_R g1055 ( 
.A(n_197),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_290),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_808),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_277),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_938),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_613),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_1026),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_853),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_212),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_954),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_553),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_337),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_646),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_859),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_12),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_354),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_722),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_95),
.Y(n_1072)
);

CKINVDCx16_ASAP7_75t_R g1073 ( 
.A(n_718),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_302),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_507),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_831),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_549),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_489),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_770),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_233),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_900),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_564),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_991),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_327),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_999),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_969),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_427),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_225),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_665),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_359),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1005),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_862),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1024),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_388),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_882),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_833),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1009),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_253),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_392),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_97),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_765),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_509),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_432),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_958),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_766),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_195),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_827),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_932),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_672),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_273),
.Y(n_1110)
);

INVx4_ASAP7_75t_R g1111 ( 
.A(n_304),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_13),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_614),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_732),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_510),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_467),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_933),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_976),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_879),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_734),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_53),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_41),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_41),
.Y(n_1123)
);

CKINVDCx16_ASAP7_75t_R g1124 ( 
.A(n_948),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_799),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1023),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_823),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_774),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_197),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_992),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_712),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_988),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_125),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_826),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_977),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_839),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_982),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_730),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_411),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_646),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_166),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_527),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_485),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_288),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_351),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_898),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_419),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_506),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_929),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_37),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_65),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_943),
.Y(n_1152)
);

BUFx5_ASAP7_75t_L g1153 ( 
.A(n_939),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_858),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_872),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_989),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_794),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_655),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_869),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_239),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_604),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_297),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_867),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_72),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1012),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_499),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_398),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_126),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_195),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_724),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_826),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_886),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_807),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_9),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_711),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_690),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_14),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_399),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_854),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_187),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_125),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_355),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_476),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_191),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_997),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_402),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_617),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_803),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_857),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_462),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_820),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_213),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_553),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_928),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_18),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_547),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_885),
.Y(n_1197)
);

BUFx10_ASAP7_75t_L g1198 ( 
.A(n_840),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_65),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_166),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_892),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_257),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_877),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1002),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_14),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_61),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_142),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_88),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_674),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_245),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_848),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_140),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_792),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_429),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_446),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_192),
.Y(n_1216)
);

BUFx10_ASAP7_75t_L g1217 ( 
.A(n_515),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_722),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_931),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_448),
.Y(n_1220)
);

BUFx5_ASAP7_75t_L g1221 ( 
.A(n_257),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_961),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_494),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_54),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_170),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_794),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_369),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_441),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_864),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_310),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_891),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_720),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_33),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_28),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1020),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_501),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_888),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1014),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_318),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1029),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_818),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_881),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_690),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_73),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_639),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_710),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_613),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_421),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_942),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_754),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_490),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_338),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_436),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_662),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_387),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_371),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_46),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1027),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_786),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_287),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_535),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_893),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_979),
.Y(n_1263)
);

INVxp33_ASAP7_75t_L g1264 ( 
.A(n_901),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1004),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_470),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_845),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_923),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_921),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_885),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_133),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_877),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_372),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_974),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1011),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_855),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_626),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_453),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_864),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_859),
.Y(n_1280)
);

BUFx10_ASAP7_75t_L g1281 ( 
.A(n_940),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_81),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_226),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_809),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_688),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_95),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_685),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_672),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_803),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_880),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_242),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_238),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_181),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_883),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_930),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_50),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_566),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_876),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_874),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_736),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_905),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_827),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_882),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_572),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_536),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_938),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_347),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_831),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1000),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_744),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_705),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_228),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_147),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_711),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_847),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_835),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_78),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_557),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_525),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_786),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_363),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_962),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_543),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_741),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_657),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_92),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_967),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_43),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_763),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_476),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_936),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_81),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_484),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_411),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_901),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_132),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_457),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_895),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_431),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_526),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_922),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_996),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_868),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_32),
.Y(n_1344)
);

CKINVDCx16_ASAP7_75t_R g1345 ( 
.A(n_371),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_968),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_330),
.Y(n_1347)
);

CKINVDCx14_ASAP7_75t_R g1348 ( 
.A(n_998),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_800),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_904),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_925),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_884),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_184),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_448),
.Y(n_1354)
);

CKINVDCx14_ASAP7_75t_R g1355 ( 
.A(n_873),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_240),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_111),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_386),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1018),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_136),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_350),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_828),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_611),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_805),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_579),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_707),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_211),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_978),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_781),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_808),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_790),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_900),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1022),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_401),
.Y(n_1374)
);

BUFx8_ASAP7_75t_SL g1375 ( 
.A(n_801),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_214),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_902),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_217),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_950),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_785),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_915),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_815),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_995),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_490),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_437),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1007),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_511),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_781),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_566),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_481),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_108),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_844),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_679),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_897),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_330),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_72),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1019),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_236),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_562),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_338),
.Y(n_1400)
);

BUFx8_ASAP7_75t_SL g1401 ( 
.A(n_402),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_843),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_675),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_141),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_161),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_409),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_424),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_388),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_382),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_358),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_395),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_871),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_935),
.Y(n_1413)
);

CKINVDCx16_ASAP7_75t_R g1414 ( 
.A(n_986),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_441),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_906),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_138),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_908),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_328),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_209),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_943),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_800),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_194),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_937),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_904),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_463),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_136),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_160),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_817),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_751),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_783),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_634),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_295),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_750),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_290),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_218),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_855),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_229),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_738),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_751),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_923),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_774),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_519),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_940),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1028),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_994),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_101),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_394),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_450),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_682),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_113),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_863),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1008),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_208),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_397),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_806),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1016),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_301),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_799),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_344),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_626),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_360),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_488),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_536),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_615),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_756),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_475),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_795),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_847),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_848),
.Y(n_1470)
);

BUFx5_ASAP7_75t_L g1471 ( 
.A(n_121),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_918),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_910),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_856),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_467),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_686),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_681),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_899),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_277),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_73),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_838),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_498),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_156),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_47),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_39),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_818),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_568),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_308),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_836),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_650),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_983),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_300),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_896),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_458),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_716),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_220),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_133),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_504),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_305),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_750),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_693),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_485),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_813),
.Y(n_1503)
);

INVxp33_ASAP7_75t_R g1504 ( 
.A(n_783),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_840),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_500),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_5),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_917),
.Y(n_1508)
);

BUFx10_ASAP7_75t_L g1509 ( 
.A(n_216),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_765),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_137),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_903),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_163),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_498),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_67),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_375),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_387),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_876),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_934),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_780),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_580),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_89),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1006),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_145),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_364),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_374),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_837),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_155),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_592),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_858),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1021),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_649),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1025),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_647),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_509),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_577),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_911),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_892),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_35),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_302),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_801),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_303),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_273),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_293),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_417),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_706),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_82),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_866),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_452),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_19),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_852),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_821),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_677),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_796),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_917),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_252),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_343),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_810),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_898),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_426),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_311),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_390),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_606),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_230),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_888),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_588),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_354),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_256),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_581),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_554),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_947),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_337),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_883),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_670),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_283),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_942),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_454),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_573),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_916),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_372),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_183),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_61),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_274),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_946),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_532),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_331),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_832),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_540),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_308),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_872),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_473),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_886),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_887),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_40),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_573),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_640),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_769),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_2),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_755),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_834),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_779),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_203),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_17),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_720),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_90),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_325),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_298),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_810),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_667),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_965),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_362),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_91),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_88),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_766),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_217),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_399),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_179),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_343),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_316),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_299),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_561),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_348),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_271),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_890),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_176),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_735),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_990),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_62),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_919),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_912),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_824),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_443),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_805),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_878),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1015),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_703),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_389),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_473),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_369),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_386),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_511),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_279),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_705),
.Y(n_1643)
);

BUFx10_ASAP7_75t_L g1644 ( 
.A(n_907),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_873),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_775),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_183),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_507),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_641),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_204),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_191),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_742),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_278),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1013),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_860),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_993),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_396),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_349),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_655),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_306),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_221),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_718),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_875),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_586),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_286),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_842),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_606),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_804),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_867),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_846),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_172),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_577),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_772),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_924),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_921),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_767),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_912),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_533),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_434),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_216),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_426),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_957),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_819),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_300),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1001),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_305),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_15),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_582),
.Y(n_1688)
);

CKINVDCx16_ASAP7_75t_R g1689 ( 
.A(n_110),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_266),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_933),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_586),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_920),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_320),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_987),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_642),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_784),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_283),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_920),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_22),
.Y(n_1700)
);

CKINVDCx16_ASAP7_75t_R g1701 ( 
.A(n_868),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_865),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_68),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_423),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_214),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_368),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_893),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_841),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_716),
.Y(n_1709)
);

CKINVDCx14_ASAP7_75t_R g1710 ( 
.A(n_228),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_400),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_420),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_857),
.Y(n_1713)
);

INVxp33_ASAP7_75t_SL g1714 ( 
.A(n_687),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_850),
.Y(n_1715)
);

CKINVDCx16_ASAP7_75t_R g1716 ( 
.A(n_812),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_865),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_908),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_698),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_27),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_630),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_29),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_890),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_389),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_555),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_604),
.Y(n_1726)
);

BUFx2_ASAP7_75t_SL g1727 ( 
.A(n_650),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_773),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_250),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_980),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_913),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_944),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_205),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_11),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_436),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_109),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_721),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_176),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1017),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_927),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_836),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_763),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_714),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_796),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_462),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_822),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_771),
.Y(n_1747)
);

BUFx10_ASAP7_75t_L g1748 ( 
.A(n_272),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_319),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1003),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_229),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_335),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_631),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_561),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_849),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_926),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_589),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_902),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_98),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_121),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_656),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_931),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_830),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_878),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_239),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_18),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_636),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_686),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_554),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_692),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_714),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_515),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_379),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_702),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_461),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_984),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_532),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_628),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_687),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_560),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_843),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_723),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_653),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_945),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_547),
.Y(n_1785)
);

BUFx8_ASAP7_75t_SL g1786 ( 
.A(n_681),
.Y(n_1786)
);

CKINVDCx16_ASAP7_75t_R g1787 ( 
.A(n_335),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_334),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_265),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_393),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_113),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_145),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_683),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_816),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_555),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_572),
.Y(n_1796)
);

BUFx10_ASAP7_75t_L g1797 ( 
.A(n_404),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_174),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_298),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_405),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_815),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_519),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_594),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_112),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_292),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_889),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_854),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_220),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_117),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_340),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_99),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_506),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_571),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_633),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_640),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_425),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_590),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_792),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_789),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_8),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_137),
.Y(n_1821)
);

BUFx10_ASAP7_75t_L g1822 ( 
.A(n_331),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_814),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_168),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_752),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_408),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_909),
.Y(n_1827)
);

BUFx10_ASAP7_75t_L g1828 ( 
.A(n_169),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_491),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_84),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_787),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_851),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_753),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_829),
.Y(n_1834)
);

CKINVDCx16_ASAP7_75t_R g1835 ( 
.A(n_504),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_428),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_13),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_93),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_811),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_115),
.Y(n_1840)
);

CKINVDCx16_ASAP7_75t_R g1841 ( 
.A(n_948),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_688),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_590),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_11),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_914),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_323),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_323),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_825),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_541),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_275),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_499),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_918),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_802),
.Y(n_1853)
);

BUFx5_ASAP7_75t_L g1854 ( 
.A(n_746),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_610),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_861),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_101),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_56),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_596),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_679),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_147),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_178),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_824),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_48),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_869),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_788),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_321),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_694),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_804),
.Y(n_1869)
);

BUFx8_ASAP7_75t_SL g1870 ( 
.A(n_552),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_175),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_126),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_941),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_25),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_691),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_7),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_393),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_633),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_360),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_894),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_75),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_505),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_22),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_224),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_63),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_798),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_870),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_361),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_173),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_34),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1441),
.Y(n_1891)
);

INVxp33_ASAP7_75t_L g1892 ( 
.A(n_1270),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1441),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1110),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1441),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1355),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1851),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1851),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1153),
.B(n_0),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1851),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1039),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1039),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1120),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1081),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1081),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1193),
.Y(n_1906)
);

INVxp33_ASAP7_75t_L g1907 ( 
.A(n_1351),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1163),
.Y(n_1908)
);

CKINVDCx20_ASAP7_75t_R g1909 ( 
.A(n_1355),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1417),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1153),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1163),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1053),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1184),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_1710),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1184),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1710),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1205),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1205),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1227),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1227),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1245),
.Y(n_1922)
);

BUFx2_ASAP7_75t_SL g1923 ( 
.A(n_1327),
.Y(n_1923)
);

CKINVDCx14_ASAP7_75t_R g1924 ( 
.A(n_1348),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1375),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1245),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1279),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1375),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1279),
.Y(n_1929)
);

INVxp33_ASAP7_75t_L g1930 ( 
.A(n_1674),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1284),
.Y(n_1931)
);

INVxp67_ASAP7_75t_SL g1932 ( 
.A(n_1284),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1286),
.Y(n_1933)
);

CKINVDCx14_ASAP7_75t_R g1934 ( 
.A(n_1348),
.Y(n_1934)
);

CKINVDCx16_ASAP7_75t_R g1935 ( 
.A(n_1034),
.Y(n_1935)
);

CKINVDCx20_ASAP7_75t_R g1936 ( 
.A(n_1401),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1286),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1053),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1291),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1291),
.Y(n_1940)
);

INVxp33_ASAP7_75t_SL g1941 ( 
.A(n_1818),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1295),
.Y(n_1942)
);

INVxp67_ASAP7_75t_SL g1943 ( 
.A(n_1295),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1304),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1304),
.Y(n_1945)
);

INVxp67_ASAP7_75t_SL g1946 ( 
.A(n_1318),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1318),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1356),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1356),
.Y(n_1949)
);

CKINVDCx16_ASAP7_75t_R g1950 ( 
.A(n_1044),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1369),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1369),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1500),
.Y(n_1953)
);

INVxp67_ASAP7_75t_SL g1954 ( 
.A(n_1500),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1528),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1528),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1530),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1327),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1530),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1268),
.Y(n_1960)
);

INVxp67_ASAP7_75t_SL g1961 ( 
.A(n_1548),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1548),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1565),
.Y(n_1963)
);

CKINVDCx16_ASAP7_75t_R g1964 ( 
.A(n_1055),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1401),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1565),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1299),
.Y(n_1967)
);

INVxp67_ASAP7_75t_SL g1968 ( 
.A(n_1614),
.Y(n_1968)
);

INVxp67_ASAP7_75t_SL g1969 ( 
.A(n_1614),
.Y(n_1969)
);

INVxp67_ASAP7_75t_SL g1970 ( 
.A(n_1642),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1642),
.Y(n_1971)
);

INVxp33_ASAP7_75t_SL g1972 ( 
.A(n_1307),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1786),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1856),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1856),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1053),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1866),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1316),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1866),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1153),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1357),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1153),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1153),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1153),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1153),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1221),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1512),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1221),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1221),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1221),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1221),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1221),
.Y(n_1992)
);

CKINVDCx14_ASAP7_75t_R g1993 ( 
.A(n_1327),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1221),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1471),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1471),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1471),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1786),
.Y(n_1998)
);

INVxp67_ASAP7_75t_SL g1999 ( 
.A(n_1112),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1471),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1471),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1471),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1471),
.Y(n_2003)
);

INVxp33_ASAP7_75t_SL g2004 ( 
.A(n_1590),
.Y(n_2004)
);

CKINVDCx20_ASAP7_75t_R g2005 ( 
.A(n_1870),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1870),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1854),
.Y(n_2007)
);

CKINVDCx20_ASAP7_75t_R g2008 ( 
.A(n_1046),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1073),
.Y(n_2009)
);

INVxp33_ASAP7_75t_SL g2010 ( 
.A(n_1636),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1854),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1854),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1112),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1657),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1854),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1854),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1854),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1854),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1124),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1033),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1036),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1040),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1041),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1063),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1070),
.Y(n_2025)
);

INVxp33_ASAP7_75t_SL g2026 ( 
.A(n_1889),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1164),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1076),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1345),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1087),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1689),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1089),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1090),
.Y(n_2033)
);

CKINVDCx20_ASAP7_75t_R g2034 ( 
.A(n_1046),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1094),
.Y(n_2035)
);

INVxp67_ASAP7_75t_SL g2036 ( 
.A(n_1112),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1727),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1099),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1100),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1101),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1701),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1240),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1108),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1716),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1114),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1119),
.Y(n_2046)
);

INVxp33_ASAP7_75t_SL g2047 ( 
.A(n_1889),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1122),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1123),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1134),
.Y(n_2050)
);

CKINVDCx20_ASAP7_75t_R g2051 ( 
.A(n_1240),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1263),
.Y(n_2052)
);

CKINVDCx14_ASAP7_75t_R g2053 ( 
.A(n_1379),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1138),
.Y(n_2054)
);

INVxp67_ASAP7_75t_SL g2055 ( 
.A(n_1112),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1144),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1145),
.Y(n_2057)
);

CKINVDCx20_ASAP7_75t_R g2058 ( 
.A(n_1263),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1171),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1148),
.Y(n_2060)
);

CKINVDCx20_ASAP7_75t_R g2061 ( 
.A(n_1342),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1149),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1787),
.Y(n_2063)
);

INVxp67_ASAP7_75t_SL g2064 ( 
.A(n_1171),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1835),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1155),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_1342),
.Y(n_2067)
);

INVxp67_ASAP7_75t_SL g2068 ( 
.A(n_1171),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1157),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1158),
.Y(n_2070)
);

INVxp33_ASAP7_75t_SL g2071 ( 
.A(n_1890),
.Y(n_2071)
);

INVxp33_ASAP7_75t_SL g2072 ( 
.A(n_1890),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1160),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1167),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1210),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1213),
.Y(n_2076)
);

CKINVDCx20_ASAP7_75t_R g2077 ( 
.A(n_1386),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_1841),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1030),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1214),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1875),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1215),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1225),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1878),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1229),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1881),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1242),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1251),
.Y(n_2088)
);

OA21x2_ASAP7_75t_L g2089 ( 
.A1(n_1982),
.A2(n_1052),
.B(n_1091),
.Y(n_2089)
);

AOI22x1_ASAP7_75t_SL g2090 ( 
.A1(n_1936),
.A2(n_1071),
.B1(n_1113),
.B2(n_1068),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2013),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1958),
.B(n_1066),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_1908),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_2009),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_2019),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1903),
.B(n_1967),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1924),
.B(n_1104),
.Y(n_2097)
);

BUFx8_ASAP7_75t_L g2098 ( 
.A(n_1894),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2013),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2059),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1913),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1911),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1980),
.Y(n_2103)
);

CKINVDCx6p67_ASAP7_75t_R g2104 ( 
.A(n_2005),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1993),
.B(n_1264),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1997),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1987),
.B(n_1066),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_2014),
.B(n_1092),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1999),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1913),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2036),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_2027),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1913),
.Y(n_2113)
);

BUFx3_ASAP7_75t_L g2114 ( 
.A(n_1908),
.Y(n_2114)
);

INVxp33_ASAP7_75t_SL g2115 ( 
.A(n_1925),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_2008),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1934),
.B(n_1414),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1923),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2055),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1938),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1901),
.B(n_1126),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1931),
.B(n_1137),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1932),
.B(n_1258),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2064),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1938),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1938),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1976),
.Y(n_2127)
);

BUFx3_ASAP7_75t_L g2128 ( 
.A(n_1951),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_1976),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2068),
.Y(n_2130)
);

NOR2x1_ASAP7_75t_L g2131 ( 
.A(n_1951),
.B(n_1118),
.Y(n_2131)
);

BUFx2_ASAP7_75t_L g2132 ( 
.A(n_2029),
.Y(n_2132)
);

CKINVDCx20_ASAP7_75t_R g2133 ( 
.A(n_2034),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2053),
.B(n_1264),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1972),
.A2(n_1071),
.B1(n_1113),
.B2(n_1068),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1976),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1939),
.B(n_1265),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1891),
.Y(n_2138)
);

OA21x2_ASAP7_75t_L g2139 ( 
.A1(n_1983),
.A2(n_1052),
.B(n_1275),
.Y(n_2139)
);

BUFx12f_ASAP7_75t_L g2140 ( 
.A(n_1928),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1897),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1893),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1984),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1943),
.B(n_1322),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_SL g2145 ( 
.A1(n_2042),
.A2(n_2052),
.B1(n_2058),
.B2(n_2051),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1895),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_2031),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_2061),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1946),
.B(n_1368),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1898),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1985),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1986),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_1906),
.B(n_1092),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1954),
.B(n_1523),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1961),
.B(n_1117),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1988),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1900),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1989),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_2079),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1990),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1991),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_1902),
.Y(n_2162)
);

BUFx3_ASAP7_75t_L g2163 ( 
.A(n_1904),
.Y(n_2163)
);

INVxp33_ASAP7_75t_SL g2164 ( 
.A(n_1965),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1992),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1968),
.B(n_1117),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1969),
.B(n_1627),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1994),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1995),
.Y(n_2169)
);

BUFx3_ASAP7_75t_L g2170 ( 
.A(n_1905),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1996),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2000),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_2081),
.B(n_1379),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2026),
.B(n_1739),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_1970),
.B(n_1248),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2001),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_2067),
.Y(n_2177)
);

AOI22x1_ASAP7_75t_SL g2178 ( 
.A1(n_2077),
.A2(n_1121),
.B1(n_1141),
.B2(n_1116),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2002),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_2003),
.Y(n_2180)
);

AND2x6_ASAP7_75t_L g2181 ( 
.A(n_1912),
.B(n_1171),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_2007),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2011),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1914),
.B(n_1635),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_2012),
.Y(n_2185)
);

OAI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_2004),
.A2(n_1116),
.B1(n_1141),
.B2(n_1121),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_2015),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2016),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1916),
.B(n_1656),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2017),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_2084),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2018),
.Y(n_2192)
);

INVx4_ASAP7_75t_L g2193 ( 
.A(n_2086),
.Y(n_2193)
);

AOI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2010),
.A2(n_1445),
.B1(n_1386),
.B2(n_1189),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2020),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2021),
.Y(n_2196)
);

INVx5_ASAP7_75t_L g2197 ( 
.A(n_1935),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1918),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1919),
.B(n_1685),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_1899),
.Y(n_2200)
);

INVx6_ASAP7_75t_L g2201 ( 
.A(n_1950),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1920),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2022),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_1896),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1892),
.B(n_1069),
.Y(n_2205)
);

OA21x2_ASAP7_75t_L g2206 ( 
.A1(n_1921),
.A2(n_1776),
.B(n_1730),
.Y(n_2206)
);

BUFx6f_ASAP7_75t_L g2207 ( 
.A(n_2023),
.Y(n_2207)
);

NOR2x1_ASAP7_75t_L g2208 ( 
.A(n_1922),
.B(n_1446),
.Y(n_2208)
);

CKINVDCx11_ASAP7_75t_R g2209 ( 
.A(n_1964),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2024),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1926),
.Y(n_2211)
);

INVx4_ASAP7_75t_L g2212 ( 
.A(n_2041),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_L g2213 ( 
.A(n_2044),
.B(n_1183),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1927),
.B(n_1739),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1907),
.B(n_1069),
.Y(n_2215)
);

BUFx8_ASAP7_75t_L g2216 ( 
.A(n_1929),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_1973),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_1933),
.A2(n_1453),
.B(n_1043),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1998),
.Y(n_2219)
);

CKINVDCx8_ASAP7_75t_R g2220 ( 
.A(n_2006),
.Y(n_2220)
);

INVx3_ASAP7_75t_L g2221 ( 
.A(n_1937),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2025),
.Y(n_2222)
);

OA21x2_ASAP7_75t_L g2223 ( 
.A1(n_1940),
.A2(n_1064),
.B(n_1061),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2028),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1941),
.A2(n_1189),
.B1(n_1211),
.B2(n_1178),
.Y(n_2225)
);

OAI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_1930),
.A2(n_1211),
.B1(n_1228),
.B2(n_1178),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2030),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_2063),
.Y(n_2228)
);

INVx6_ASAP7_75t_L g2229 ( 
.A(n_1910),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_2032),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_2033),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2035),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1942),
.B(n_1083),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1944),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1945),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2038),
.Y(n_2236)
);

BUFx3_ASAP7_75t_L g2237 ( 
.A(n_1947),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_1960),
.B(n_1252),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2065),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1948),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1949),
.B(n_1085),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1952),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_2039),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_2040),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2043),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_1953),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_SL g2247 ( 
.A1(n_1909),
.A2(n_1243),
.B1(n_1250),
.B2(n_1228),
.Y(n_2247)
);

INVx6_ASAP7_75t_L g2248 ( 
.A(n_1978),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2045),
.Y(n_2249)
);

INVx4_ASAP7_75t_L g2250 ( 
.A(n_2078),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_1955),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1915),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2046),
.Y(n_2253)
);

BUFx3_ASAP7_75t_L g2254 ( 
.A(n_1956),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1957),
.B(n_1086),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_2037),
.B(n_1248),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_2047),
.B(n_1379),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_1981),
.B(n_1276),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2048),
.Y(n_2259)
);

CKINVDCx11_ASAP7_75t_R g2260 ( 
.A(n_1917),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1959),
.B(n_1276),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_2049),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2050),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2054),
.Y(n_2264)
);

INVx4_ASAP7_75t_L g2265 ( 
.A(n_1962),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1963),
.Y(n_2266)
);

INVxp67_ASAP7_75t_L g2267 ( 
.A(n_1966),
.Y(n_2267)
);

OA22x2_ASAP7_75t_SL g2268 ( 
.A1(n_2056),
.A2(n_1504),
.B1(n_1381),
.B2(n_1250),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2057),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2060),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_1971),
.Y(n_2271)
);

INVxp33_ASAP7_75t_SL g2272 ( 
.A(n_1974),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_2062),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2071),
.A2(n_1445),
.B1(n_1260),
.B2(n_1261),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_1975),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2072),
.A2(n_1260),
.B1(n_1261),
.B2(n_1243),
.Y(n_2276)
);

AND2x6_ASAP7_75t_L g2277 ( 
.A(n_1977),
.B(n_1183),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2066),
.Y(n_2278)
);

CKINVDCx6p67_ASAP7_75t_R g2279 ( 
.A(n_1979),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2069),
.Y(n_2280)
);

BUFx8_ASAP7_75t_L g2281 ( 
.A(n_2070),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_2073),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_2074),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2075),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2076),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2080),
.B(n_1069),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2082),
.B(n_1168),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_2083),
.Y(n_2288)
);

INVx4_ASAP7_75t_L g2289 ( 
.A(n_2085),
.Y(n_2289)
);

HB1xp67_ASAP7_75t_L g2290 ( 
.A(n_2087),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2088),
.B(n_1093),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2013),
.Y(n_2292)
);

OA21x2_ASAP7_75t_L g2293 ( 
.A1(n_1982),
.A2(n_1130),
.B(n_1097),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2013),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_1958),
.B(n_1287),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1999),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2013),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1924),
.B(n_1132),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2013),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1913),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2013),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2013),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1999),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_1913),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1993),
.B(n_1168),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_1913),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_1972),
.A2(n_1311),
.B1(n_1387),
.B2(n_1280),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_1993),
.B(n_1168),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_2008),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2013),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2013),
.Y(n_2311)
);

OAI22xp5_ASAP7_75t_SL g2312 ( 
.A1(n_2008),
.A2(n_1311),
.B1(n_1387),
.B2(n_1280),
.Y(n_2312)
);

OAI21x1_ASAP7_75t_L g2313 ( 
.A1(n_1911),
.A2(n_1043),
.B(n_1038),
.Y(n_2313)
);

BUFx8_ASAP7_75t_L g2314 ( 
.A(n_1894),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2013),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2013),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1924),
.B(n_1135),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1958),
.B(n_1714),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1924),
.B(n_1156),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2013),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_1993),
.B(n_1198),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1999),
.Y(n_2322)
);

BUFx8_ASAP7_75t_L g2323 ( 
.A(n_1894),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_1913),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_1958),
.B(n_1714),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1924),
.B(n_1165),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2013),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1999),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1924),
.B(n_1185),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_1913),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_1913),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2013),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_1913),
.Y(n_2333)
);

AOI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_1972),
.A2(n_1469),
.B1(n_1473),
.B2(n_1430),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_1913),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_1924),
.B(n_1204),
.Y(n_2336)
);

CKINVDCx6p67_ASAP7_75t_R g2337 ( 
.A(n_1936),
.Y(n_2337)
);

BUFx3_ASAP7_75t_L g2338 ( 
.A(n_1908),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_1958),
.B(n_1287),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1999),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_1903),
.A2(n_1469),
.B1(n_1473),
.B2(n_1430),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1999),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2013),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1999),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_2008),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2013),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2013),
.Y(n_2347)
);

INVx5_ASAP7_75t_L g2348 ( 
.A(n_1908),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1999),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1999),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_1908),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1924),
.B(n_1222),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2013),
.Y(n_2353)
);

BUFx6f_ASAP7_75t_L g2354 ( 
.A(n_1913),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1999),
.Y(n_2355)
);

INVx5_ASAP7_75t_L g2356 ( 
.A(n_1908),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_1993),
.B(n_1198),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_1993),
.B(n_1198),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_1908),
.Y(n_2359)
);

INVx6_ASAP7_75t_L g2360 ( 
.A(n_1935),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_1958),
.B(n_1323),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_1913),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1999),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_1913),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_2008),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1999),
.Y(n_2366)
);

AND2x6_ASAP7_75t_L g2367 ( 
.A(n_1958),
.B(n_1183),
.Y(n_2367)
);

BUFx3_ASAP7_75t_L g2368 ( 
.A(n_1908),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1999),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1999),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1999),
.Y(n_2371)
);

INVx5_ASAP7_75t_L g2372 ( 
.A(n_1908),
.Y(n_2372)
);

OAI21x1_ASAP7_75t_L g2373 ( 
.A1(n_1911),
.A2(n_1049),
.B(n_1038),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_SL g2374 ( 
.A1(n_2008),
.A2(n_1505),
.B1(n_1513),
.B2(n_1476),
.Y(n_2374)
);

HB1xp67_ASAP7_75t_L g2375 ( 
.A(n_2009),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_1908),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_1958),
.B(n_1323),
.Y(n_2377)
);

BUFx12f_ASAP7_75t_L g2378 ( 
.A(n_1925),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2013),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_1993),
.B(n_1217),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_1908),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2013),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1999),
.Y(n_2383)
);

INVx6_ASAP7_75t_L g2384 ( 
.A(n_1935),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1924),
.B(n_1235),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_1993),
.B(n_1217),
.Y(n_2386)
);

BUFx8_ASAP7_75t_L g2387 ( 
.A(n_1894),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2013),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_1913),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1999),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_1913),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1999),
.Y(n_2392)
);

INVx6_ASAP7_75t_L g2393 ( 
.A(n_1935),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_2008),
.Y(n_2394)
);

BUFx6f_ASAP7_75t_L g2395 ( 
.A(n_1913),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1999),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_1908),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_L g2398 ( 
.A(n_1913),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1999),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2013),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_1993),
.B(n_1217),
.Y(n_2401)
);

OA21x2_ASAP7_75t_L g2402 ( 
.A1(n_1982),
.A2(n_1274),
.B(n_1238),
.Y(n_2402)
);

INVx3_ASAP7_75t_L g2403 ( 
.A(n_1908),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_1913),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_1972),
.A2(n_1505),
.B1(n_1513),
.B2(n_1476),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_1913),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1999),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_1908),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1999),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_SL g2410 ( 
.A1(n_2008),
.A2(n_1522),
.B1(n_1537),
.B2(n_1515),
.Y(n_2410)
);

OAI21x1_ASAP7_75t_L g2411 ( 
.A1(n_1911),
.A2(n_1075),
.B(n_1049),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_1913),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1999),
.Y(n_2413)
);

CKINVDCx6p67_ASAP7_75t_R g2414 ( 
.A(n_1936),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2013),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2013),
.Y(n_2416)
);

AND2x2_ASAP7_75t_SL g2417 ( 
.A(n_1935),
.B(n_1075),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_1958),
.B(n_1333),
.Y(n_2418)
);

INVx3_ASAP7_75t_L g2419 ( 
.A(n_1908),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2013),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_1913),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_1913),
.Y(n_2422)
);

AND2x2_ASAP7_75t_SL g2423 ( 
.A(n_1935),
.B(n_1162),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_1913),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_1913),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_1993),
.B(n_1281),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1999),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2013),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1999),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2013),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_2116),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2091),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2148),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_2177),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2198),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_2309),
.Y(n_2436)
);

INVxp67_ASAP7_75t_L g2437 ( 
.A(n_2105),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2345),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_2101),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_R g2440 ( 
.A(n_2228),
.B(n_1309),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_2201),
.Y(n_2441)
);

BUFx2_ASAP7_75t_L g2442 ( 
.A(n_2248),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2202),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_2365),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2217),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_2219),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_2133),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2394),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2211),
.Y(n_2449)
);

HB1xp67_ASAP7_75t_L g2450 ( 
.A(n_2229),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_2209),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2099),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2140),
.Y(n_2453)
);

CKINVDCx16_ASAP7_75t_R g2454 ( 
.A(n_2204),
.Y(n_2454)
);

AND3x2_ASAP7_75t_L g2455 ( 
.A(n_2095),
.B(n_1159),
.C(n_1103),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_2378),
.Y(n_2456)
);

CKINVDCx20_ASAP7_75t_R g2457 ( 
.A(n_2260),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2292),
.Y(n_2458)
);

CKINVDCx20_ASAP7_75t_R g2459 ( 
.A(n_2252),
.Y(n_2459)
);

CKINVDCx16_ASAP7_75t_R g2460 ( 
.A(n_2132),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2115),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2234),
.Y(n_2462)
);

INVxp67_ASAP7_75t_L g2463 ( 
.A(n_2134),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2164),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2242),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2266),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2280),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2220),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2104),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2337),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2414),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2360),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_2147),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2285),
.Y(n_2474)
);

CKINVDCx20_ASAP7_75t_R g2475 ( 
.A(n_2384),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_L g2476 ( 
.A(n_2118),
.B(n_1333),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2159),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2193),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2138),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2142),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_R g2481 ( 
.A(n_2191),
.B(n_2393),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2348),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2098),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2294),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2314),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_R g2486 ( 
.A(n_2239),
.B(n_1346),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2297),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2146),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2114),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2323),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_2387),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2299),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2197),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_2197),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2094),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2150),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2157),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2112),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2096),
.Y(n_2499)
);

CKINVDCx5p33_ASAP7_75t_R g2500 ( 
.A(n_2375),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2174),
.B(n_1398),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2212),
.Y(n_2502)
);

NOR2xp67_ASAP7_75t_L g2503 ( 
.A(n_2250),
.B(n_2257),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2145),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2195),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2276),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2283),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2226),
.Y(n_2508)
);

BUFx8_ASAP7_75t_L g2509 ( 
.A(n_2205),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_2135),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_2186),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2301),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2225),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_2341),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2302),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2310),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2272),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_2279),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2194),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_R g2520 ( 
.A(n_2093),
.B(n_1359),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2312),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_2410),
.Y(n_2522)
);

NOR2xp67_ASAP7_75t_L g2523 ( 
.A(n_2305),
.B(n_2308),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_R g2524 ( 
.A(n_2351),
.B(n_1373),
.Y(n_2524)
);

BUFx10_ASAP7_75t_L g2525 ( 
.A(n_2318),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2311),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2196),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_2128),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2338),
.Y(n_2529)
);

CKINVDCx20_ASAP7_75t_R g2530 ( 
.A(n_2274),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2315),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2368),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_2163),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_2170),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_2237),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2254),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2203),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2275),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_2281),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2417),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2316),
.Y(n_2541)
);

CKINVDCx6p67_ASAP7_75t_R g2542 ( 
.A(n_2423),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2178),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2101),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_R g2545 ( 
.A(n_2359),
.B(n_1383),
.Y(n_2545)
);

CKINVDCx20_ASAP7_75t_R g2546 ( 
.A(n_2307),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2247),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2374),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_2216),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2200),
.Y(n_2550)
);

CKINVDCx5p33_ASAP7_75t_R g2551 ( 
.A(n_2200),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2215),
.B(n_1281),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_R g2553 ( 
.A(n_2376),
.B(n_1397),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2367),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2287),
.A2(n_1522),
.B1(n_1537),
.B2(n_1515),
.Y(n_2555)
);

BUFx10_ASAP7_75t_L g2556 ( 
.A(n_2325),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2320),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_R g2558 ( 
.A(n_2381),
.B(n_1457),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_R g2559 ( 
.A(n_2397),
.B(n_1491),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_2367),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2321),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2327),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2334),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2405),
.Y(n_2564)
);

NAND2xp33_ASAP7_75t_R g2565 ( 
.A(n_2293),
.B(n_1031),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2403),
.Y(n_2566)
);

CKINVDCx20_ASAP7_75t_R g2567 ( 
.A(n_2357),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_2090),
.Y(n_2568)
);

NAND2xp33_ASAP7_75t_R g2569 ( 
.A(n_2402),
.B(n_1032),
.Y(n_2569)
);

INVxp67_ASAP7_75t_L g2570 ( 
.A(n_2358),
.Y(n_2570)
);

BUFx2_ASAP7_75t_L g2571 ( 
.A(n_2380),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_2408),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2290),
.Y(n_2573)
);

HB1xp67_ASAP7_75t_L g2574 ( 
.A(n_2419),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2386),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2332),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2401),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2426),
.Y(n_2578)
);

INVx2_ASAP7_75t_SL g2579 ( 
.A(n_2097),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_R g2580 ( 
.A(n_2213),
.B(n_1531),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2343),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_R g2582 ( 
.A(n_2162),
.B(n_2221),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2210),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2117),
.B(n_1035),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2207),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2346),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2155),
.A2(n_1559),
.B1(n_1566),
.B2(n_1558),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2207),
.Y(n_2588)
);

CKINVDCx20_ASAP7_75t_R g2589 ( 
.A(n_2173),
.Y(n_2589)
);

CKINVDCx16_ASAP7_75t_R g2590 ( 
.A(n_2153),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2158),
.B(n_1533),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2347),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2230),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2222),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2230),
.Y(n_2595)
);

NAND2xp33_ASAP7_75t_L g2596 ( 
.A(n_2165),
.B(n_1183),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2224),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_2231),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2231),
.Y(n_2599)
);

CKINVDCx20_ASAP7_75t_R g2600 ( 
.A(n_2298),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2227),
.Y(n_2601)
);

CKINVDCx20_ASAP7_75t_R g2602 ( 
.A(n_2317),
.Y(n_2602)
);

XOR2xp5_ASAP7_75t_L g2603 ( 
.A(n_2208),
.B(n_1558),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2232),
.Y(n_2604)
);

BUFx2_ASAP7_75t_L g2605 ( 
.A(n_2238),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2353),
.Y(n_2606)
);

CKINVDCx20_ASAP7_75t_R g2607 ( 
.A(n_2319),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2243),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2243),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2244),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2236),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_2244),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_SL g2613 ( 
.A(n_2258),
.Y(n_2613)
);

NOR2xp33_ASAP7_75t_R g2614 ( 
.A(n_2235),
.B(n_1610),
.Y(n_2614)
);

CKINVDCx20_ASAP7_75t_R g2615 ( 
.A(n_2326),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2379),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2262),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2113),
.Y(n_2618)
);

OR2x2_ASAP7_75t_L g2619 ( 
.A(n_2107),
.B(n_1058),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2108),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2245),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_2262),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2249),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2263),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2263),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2113),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2166),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2121),
.B(n_1060),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2382),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2253),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2388),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2270),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2175),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2270),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2109),
.B(n_1398),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2127),
.Y(n_2636)
);

CKINVDCx5p33_ASAP7_75t_R g2637 ( 
.A(n_2273),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2273),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2282),
.Y(n_2639)
);

NOR2xp67_ASAP7_75t_L g2640 ( 
.A(n_2348),
.B(n_2356),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2400),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2259),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2127),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2264),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2092),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2269),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2282),
.Y(n_2647)
);

AND2x6_ASAP7_75t_L g2648 ( 
.A(n_2131),
.B(n_1053),
.Y(n_2648)
);

NAND2xp33_ASAP7_75t_R g2649 ( 
.A(n_2223),
.B(n_2206),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2278),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_R g2651 ( 
.A(n_2240),
.B(n_1654),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_R g2652 ( 
.A(n_2246),
.B(n_1682),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2284),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2284),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_R g2655 ( 
.A(n_2251),
.B(n_1695),
.Y(n_2655)
);

CKINVDCx20_ASAP7_75t_R g2656 ( 
.A(n_2329),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_2288),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2288),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2415),
.Y(n_2659)
);

NOR2xp67_ASAP7_75t_L g2660 ( 
.A(n_2356),
.B(n_1750),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2129),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2336),
.Y(n_2662)
);

CKINVDCx5p33_ASAP7_75t_R g2663 ( 
.A(n_2352),
.Y(n_2663)
);

BUFx2_ASAP7_75t_L g2664 ( 
.A(n_2295),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_2385),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2256),
.B(n_1281),
.Y(n_2666)
);

XNOR2xp5_ASAP7_75t_L g2667 ( 
.A(n_2286),
.B(n_1559),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2416),
.Y(n_2668)
);

CKINVDCx20_ASAP7_75t_R g2669 ( 
.A(n_2267),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_R g2670 ( 
.A(n_2271),
.B(n_2111),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2265),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_2289),
.Y(n_2672)
);

CKINVDCx20_ASAP7_75t_R g2673 ( 
.A(n_2372),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2119),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2372),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2420),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_2233),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2124),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2241),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2255),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2291),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_2130),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_2296),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_2303),
.Y(n_2684)
);

INVx5_ASAP7_75t_L g2685 ( 
.A(n_2181),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2322),
.Y(n_2686)
);

HB1xp67_ASAP7_75t_L g2687 ( 
.A(n_2339),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2328),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2340),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2342),
.Y(n_2690)
);

CKINVDCx20_ASAP7_75t_R g2691 ( 
.A(n_2122),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2344),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2349),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2361),
.B(n_1037),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2350),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2355),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2363),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2366),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2369),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2370),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2371),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2383),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2390),
.Y(n_2703)
);

BUFx3_ASAP7_75t_L g2704 ( 
.A(n_2392),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2396),
.Y(n_2705)
);

CKINVDCx20_ASAP7_75t_R g2706 ( 
.A(n_2123),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2399),
.Y(n_2707)
);

CKINVDCx20_ASAP7_75t_R g2708 ( 
.A(n_2137),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_2407),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2409),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2413),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_2427),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_R g2713 ( 
.A(n_2429),
.B(n_1042),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2151),
.Y(n_2714)
);

BUFx10_ASAP7_75t_L g2715 ( 
.A(n_2377),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2144),
.Y(n_2716)
);

BUFx3_ASAP7_75t_L g2717 ( 
.A(n_2141),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2149),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_2154),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_2167),
.Y(n_2720)
);

INVxp33_ASAP7_75t_SL g2721 ( 
.A(n_2214),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2152),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2418),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2156),
.Y(n_2724)
);

CKINVDCx20_ASAP7_75t_R g2725 ( 
.A(n_2184),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2161),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2189),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2168),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2129),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2183),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2261),
.B(n_1326),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_R g2732 ( 
.A(n_2169),
.B(n_1045),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_2199),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2143),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2192),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2428),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2102),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2143),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2475),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2716),
.B(n_2172),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2432),
.Y(n_2741)
);

INVx2_ASAP7_75t_SL g2742 ( 
.A(n_2442),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2718),
.B(n_2176),
.Y(n_2743)
);

INVx3_ASAP7_75t_L g2744 ( 
.A(n_2441),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2445),
.Y(n_2745)
);

INVx1_ASAP7_75t_SL g2746 ( 
.A(n_2450),
.Y(n_2746)
);

OR2x2_ASAP7_75t_L g2747 ( 
.A(n_2605),
.B(n_1128),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2674),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2452),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2458),
.Y(n_2750)
);

NAND2xp33_ASAP7_75t_L g2751 ( 
.A(n_2477),
.B(n_2179),
.Y(n_2751)
);

NAND2xp33_ASAP7_75t_L g2752 ( 
.A(n_2478),
.B(n_2188),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2719),
.B(n_2190),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2720),
.B(n_2160),
.Y(n_2754)
);

INVx3_ASAP7_75t_L g2755 ( 
.A(n_2472),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2678),
.Y(n_2756)
);

NAND2xp33_ASAP7_75t_L g2757 ( 
.A(n_2502),
.B(n_2160),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2692),
.Y(n_2758)
);

BUFx10_ASAP7_75t_L g2759 ( 
.A(n_2446),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2721),
.B(n_2171),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2579),
.B(n_2171),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2459),
.Y(n_2762)
);

INVxp67_ASAP7_75t_L g2763 ( 
.A(n_2499),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2484),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2717),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2727),
.B(n_2180),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2489),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2487),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2693),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2698),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2517),
.B(n_2180),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2681),
.B(n_2182),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2677),
.B(n_2182),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2699),
.Y(n_2774)
);

INVx4_ASAP7_75t_L g2775 ( 
.A(n_2468),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2507),
.B(n_1566),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2679),
.B(n_2185),
.Y(n_2777)
);

BUFx6f_ASAP7_75t_L g2778 ( 
.A(n_2544),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_SL g2779 ( 
.A(n_2680),
.B(n_2185),
.Y(n_2779)
);

AND2x4_ASAP7_75t_L g2780 ( 
.A(n_2473),
.B(n_1567),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2705),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2711),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_L g2783 ( 
.A1(n_2514),
.A2(n_2103),
.B1(n_2106),
.B2(n_2089),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2733),
.B(n_2187),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2505),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2501),
.A2(n_2187),
.B1(n_1582),
.B2(n_1586),
.Y(n_2786)
);

NOR2x1p5_ASAP7_75t_L g2787 ( 
.A(n_2461),
.B(n_1047),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2527),
.Y(n_2788)
);

INVx5_ASAP7_75t_L g2789 ( 
.A(n_2460),
.Y(n_2789)
);

NAND2x1p5_ASAP7_75t_L g2790 ( 
.A(n_2561),
.B(n_2430),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_SL g2791 ( 
.A(n_2503),
.B(n_1048),
.Y(n_2791)
);

OR2x6_ASAP7_75t_L g2792 ( 
.A(n_2627),
.B(n_2268),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2492),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2523),
.B(n_1567),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2662),
.B(n_2663),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2633),
.B(n_1582),
.Y(n_2796)
);

INVx3_ASAP7_75t_L g2797 ( 
.A(n_2585),
.Y(n_2797)
);

BUFx2_ASAP7_75t_L g2798 ( 
.A(n_2447),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2665),
.B(n_2218),
.Y(n_2799)
);

NOR2x1p5_ASAP7_75t_L g2800 ( 
.A(n_2464),
.B(n_1050),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2588),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2512),
.Y(n_2802)
);

OAI22xp33_ASAP7_75t_L g2803 ( 
.A1(n_2506),
.A2(n_1586),
.B1(n_1605),
.B2(n_1599),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2537),
.Y(n_2804)
);

INVx4_ASAP7_75t_L g2805 ( 
.A(n_2453),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2431),
.B(n_1599),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2515),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2448),
.Y(n_2808)
);

AND2x4_ASAP7_75t_L g2809 ( 
.A(n_2433),
.B(n_1605),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2440),
.B(n_1051),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2437),
.B(n_1146),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2583),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2594),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_SL g2814 ( 
.A(n_2550),
.B(n_1054),
.Y(n_2814)
);

INVx4_ASAP7_75t_L g2815 ( 
.A(n_2456),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2463),
.B(n_2570),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2597),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2516),
.Y(n_2818)
);

INVxp67_ASAP7_75t_SL g2819 ( 
.A(n_2566),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2551),
.B(n_1056),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2526),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2628),
.B(n_2139),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2531),
.Y(n_2823)
);

OR2x6_ASAP7_75t_L g2824 ( 
.A(n_2620),
.B(n_1416),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2601),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2544),
.Y(n_2826)
);

NAND2xp33_ASAP7_75t_L g2827 ( 
.A(n_2486),
.B(n_1278),
.Y(n_2827)
);

AND2x6_ASAP7_75t_L g2828 ( 
.A(n_2552),
.B(n_1162),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2544),
.Y(n_2829)
);

INVx1_ASAP7_75t_SL g2830 ( 
.A(n_2481),
.Y(n_2830)
);

BUFx6f_ASAP7_75t_L g2831 ( 
.A(n_2636),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2636),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2541),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2604),
.B(n_2100),
.Y(n_2834)
);

NAND2xp33_ASAP7_75t_R g2835 ( 
.A(n_2434),
.B(n_2313),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2573),
.B(n_1057),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2593),
.Y(n_2837)
);

NAND2xp33_ASAP7_75t_L g2838 ( 
.A(n_2672),
.B(n_1278),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2571),
.B(n_1616),
.Y(n_2839)
);

CKINVDCx11_ASAP7_75t_R g2840 ( 
.A(n_2457),
.Y(n_2840)
);

INVx5_ASAP7_75t_L g2841 ( 
.A(n_2715),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2611),
.B(n_2181),
.Y(n_2842)
);

CKINVDCx20_ASAP7_75t_R g2843 ( 
.A(n_2436),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2621),
.Y(n_2844)
);

INVxp67_ASAP7_75t_SL g2845 ( 
.A(n_2574),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2623),
.B(n_2277),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2557),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2630),
.Y(n_2848)
);

AND2x4_ASAP7_75t_L g2849 ( 
.A(n_2438),
.B(n_1616),
.Y(n_2849)
);

AND2x6_ASAP7_75t_L g2850 ( 
.A(n_2666),
.B(n_1226),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2562),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2642),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2636),
.Y(n_2853)
);

NAND2xp33_ASAP7_75t_L g2854 ( 
.A(n_2671),
.B(n_1278),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2644),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2645),
.B(n_1643),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2646),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2650),
.Y(n_2858)
);

INVx1_ASAP7_75t_SL g2859 ( 
.A(n_2669),
.Y(n_2859)
);

OAI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2479),
.A2(n_1421),
.B1(n_1427),
.B2(n_1367),
.Y(n_2860)
);

AOI22xp33_ASAP7_75t_L g2861 ( 
.A1(n_2508),
.A2(n_1709),
.B1(n_1793),
.B2(n_1643),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2480),
.Y(n_2862)
);

BUFx6f_ASAP7_75t_L g2863 ( 
.A(n_2661),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2488),
.B(n_2277),
.Y(n_2864)
);

INVx5_ASAP7_75t_L g2865 ( 
.A(n_2715),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2496),
.B(n_1416),
.Y(n_2866)
);

INVx6_ASAP7_75t_L g2867 ( 
.A(n_2454),
.Y(n_2867)
);

AND2x6_ASAP7_75t_L g2868 ( 
.A(n_2731),
.B(n_1226),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2590),
.B(n_1188),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2525),
.B(n_1200),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2525),
.B(n_1209),
.Y(n_2871)
);

CKINVDCx5p33_ASAP7_75t_R g2872 ( 
.A(n_2444),
.Y(n_2872)
);

INVx3_ASAP7_75t_L g2873 ( 
.A(n_2595),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2497),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2598),
.Y(n_2875)
);

BUFx6f_ASAP7_75t_L g2876 ( 
.A(n_2661),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2435),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2443),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2467),
.B(n_1638),
.Y(n_2879)
);

BUFx3_ASAP7_75t_L g2880 ( 
.A(n_2599),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2556),
.B(n_1246),
.Y(n_2881)
);

OR2x2_ASAP7_75t_L g2882 ( 
.A(n_2619),
.B(n_1329),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2495),
.Y(n_2883)
);

NAND2x1p5_ASAP7_75t_L g2884 ( 
.A(n_2572),
.B(n_1404),
.Y(n_2884)
);

BUFx2_ASAP7_75t_L g2885 ( 
.A(n_2498),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2449),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2474),
.B(n_2682),
.Y(n_2887)
);

AOI22xp33_ASAP7_75t_L g2888 ( 
.A1(n_2513),
.A2(n_2511),
.B1(n_2510),
.B2(n_2714),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2576),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2462),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2465),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2608),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2581),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2683),
.B(n_1638),
.Y(n_2894)
);

INVx3_ASAP7_75t_L g2895 ( 
.A(n_2609),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2610),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2586),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2592),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2556),
.B(n_2723),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_SL g2900 ( 
.A(n_2528),
.B(n_1059),
.Y(n_2900)
);

BUFx4_ASAP7_75t_L g2901 ( 
.A(n_2483),
.Y(n_2901)
);

BUFx3_ASAP7_75t_L g2902 ( 
.A(n_2612),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2617),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2606),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2622),
.Y(n_2905)
);

BUFx2_ASAP7_75t_L g2906 ( 
.A(n_2500),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2575),
.B(n_2577),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2466),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2684),
.B(n_2373),
.Y(n_2909)
);

INVx3_ASAP7_75t_L g2910 ( 
.A(n_2624),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2686),
.B(n_2411),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2722),
.Y(n_2912)
);

BUFx3_ASAP7_75t_L g2913 ( 
.A(n_2625),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2688),
.B(n_1256),
.Y(n_2914)
);

AND3x2_ASAP7_75t_L g2915 ( 
.A(n_2664),
.B(n_2687),
.C(n_2490),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2690),
.B(n_1494),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2578),
.B(n_1709),
.Y(n_2917)
);

AND2x4_ASAP7_75t_L g2918 ( 
.A(n_2518),
.B(n_1793),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_2695),
.B(n_1502),
.Y(n_2919)
);

INVx1_ASAP7_75t_SL g2920 ( 
.A(n_2533),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2696),
.B(n_1543),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2616),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2724),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2726),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2728),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2730),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2735),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2629),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2542),
.B(n_1831),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2534),
.B(n_1831),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2697),
.B(n_1552),
.Y(n_2931)
);

BUFx10_ASAP7_75t_L g2932 ( 
.A(n_2451),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2700),
.B(n_2701),
.Y(n_2933)
);

BUFx10_ASAP7_75t_L g2934 ( 
.A(n_2493),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2737),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2631),
.Y(n_2936)
);

INVx4_ASAP7_75t_L g2937 ( 
.A(n_2632),
.Y(n_2937)
);

INVx4_ASAP7_75t_SL g2938 ( 
.A(n_2613),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2641),
.Y(n_2939)
);

INVxp67_ASAP7_75t_L g2940 ( 
.A(n_2613),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2529),
.B(n_1062),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2689),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2532),
.B(n_1065),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2659),
.Y(n_2944)
);

AND2x6_ASAP7_75t_L g2945 ( 
.A(n_2704),
.B(n_1256),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2668),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2661),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2676),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_2702),
.B(n_1598),
.Y(n_2949)
);

INVx1_ASAP7_75t_SL g2950 ( 
.A(n_2535),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2634),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2591),
.A2(n_1842),
.B1(n_1072),
.B2(n_1074),
.Y(n_2952)
);

NOR2x1p5_ASAP7_75t_L g2953 ( 
.A(n_2539),
.B(n_1067),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_2729),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2736),
.Y(n_2955)
);

BUFx3_ASAP7_75t_L g2956 ( 
.A(n_2637),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2439),
.Y(n_2957)
);

CKINVDCx5p33_ASAP7_75t_R g2958 ( 
.A(n_2469),
.Y(n_2958)
);

OAI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_2587),
.A2(n_1842),
.B1(n_1670),
.B2(n_1671),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2439),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2618),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_SL g2962 ( 
.A1(n_2519),
.A2(n_2563),
.B1(n_2564),
.B2(n_2530),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2618),
.Y(n_2963)
);

INVxp67_ASAP7_75t_SL g2964 ( 
.A(n_2509),
.Y(n_2964)
);

AO22x2_ASAP7_75t_L g2965 ( 
.A1(n_2603),
.A2(n_1683),
.B1(n_1700),
.B2(n_1634),
.Y(n_2965)
);

BUFx4f_ASAP7_75t_L g2966 ( 
.A(n_2648),
.Y(n_2966)
);

A2O1A1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2476),
.A2(n_1290),
.B(n_1336),
.C(n_1271),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2626),
.Y(n_2968)
);

INVx4_ASAP7_75t_L g2969 ( 
.A(n_2638),
.Y(n_2969)
);

AND2x4_ASAP7_75t_L g2970 ( 
.A(n_2470),
.B(n_1713),
.Y(n_2970)
);

INVx5_ASAP7_75t_L g2971 ( 
.A(n_2648),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2626),
.Y(n_2972)
);

INVx4_ASAP7_75t_L g2973 ( 
.A(n_2639),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2643),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2643),
.Y(n_2975)
);

INVx4_ASAP7_75t_L g2976 ( 
.A(n_2647),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2729),
.Y(n_2977)
);

CKINVDCx20_ASAP7_75t_R g2978 ( 
.A(n_2471),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2729),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2653),
.B(n_1731),
.Y(n_2980)
);

BUFx6f_ASAP7_75t_L g2981 ( 
.A(n_2654),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2703),
.Y(n_2982)
);

AO22x2_ASAP7_75t_L g2983 ( 
.A1(n_2546),
.A2(n_2521),
.B1(n_2522),
.B2(n_2547),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2536),
.B(n_1326),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_R g2985 ( 
.A(n_2494),
.B(n_1077),
.Y(n_2985)
);

AOI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2707),
.A2(n_1807),
.B1(n_1853),
.B2(n_1762),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2772),
.B(n_2709),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2741),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2916),
.B(n_2710),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2933),
.B(n_2725),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2919),
.B(n_2921),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2748),
.Y(n_2992)
);

INVx4_ASAP7_75t_L g2993 ( 
.A(n_2745),
.Y(n_2993)
);

NOR2xp33_ASAP7_75t_L g2994 ( 
.A(n_2795),
.B(n_2691),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2749),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_SL g2996 ( 
.A(n_2762),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2750),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2982),
.B(n_2538),
.Y(n_2998)
);

HB1xp67_ASAP7_75t_L g2999 ( 
.A(n_2746),
.Y(n_2999)
);

INVx3_ASAP7_75t_L g3000 ( 
.A(n_2739),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_2742),
.Y(n_3001)
);

NAND2xp33_ASAP7_75t_L g3002 ( 
.A(n_2872),
.B(n_2554),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2920),
.B(n_2582),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2756),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2950),
.B(n_2732),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2981),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2931),
.B(n_2712),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2949),
.B(n_2734),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_2843),
.Y(n_3009)
);

A2O1A1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2816),
.A2(n_2635),
.B(n_2584),
.C(n_2555),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_2840),
.Y(n_3011)
);

NAND2xp33_ASAP7_75t_L g3012 ( 
.A(n_2785),
.B(n_2560),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2760),
.B(n_2738),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2740),
.B(n_2743),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2870),
.B(n_2871),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2881),
.B(n_2706),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2830),
.B(n_2708),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2758),
.Y(n_3018)
);

NOR2xp67_ASAP7_75t_L g3019 ( 
.A(n_2789),
.B(n_2657),
.Y(n_3019)
);

A2O1A1Ixp33_ASAP7_75t_L g3020 ( 
.A1(n_2753),
.A2(n_2660),
.B(n_2694),
.C(n_1255),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2769),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2930),
.B(n_2540),
.Y(n_3022)
);

NAND3xp33_ASAP7_75t_L g3023 ( 
.A(n_2771),
.B(n_2509),
.C(n_2667),
.Y(n_3023)
);

NAND2xp33_ASAP7_75t_L g3024 ( 
.A(n_2788),
.B(n_2520),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2770),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2774),
.Y(n_3026)
);

AND2x6_ASAP7_75t_SL g3027 ( 
.A(n_2806),
.B(n_1253),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2764),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2766),
.B(n_2614),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2761),
.B(n_2658),
.Y(n_3030)
);

BUFx5_ASAP7_75t_L g3031 ( 
.A(n_2946),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2754),
.B(n_2670),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2869),
.B(n_2567),
.Y(n_3033)
);

INVx2_ASAP7_75t_SL g3034 ( 
.A(n_2789),
.Y(n_3034)
);

BUFx8_ASAP7_75t_L g3035 ( 
.A(n_2798),
.Y(n_3035)
);

INVx2_ASAP7_75t_SL g3036 ( 
.A(n_2867),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2781),
.B(n_2648),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2804),
.A2(n_2600),
.B1(n_2607),
.B2(n_2602),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2782),
.B(n_2648),
.Y(n_3039)
);

BUFx6f_ASAP7_75t_SL g3040 ( 
.A(n_2932),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2784),
.B(n_2713),
.Y(n_3041)
);

OR2x2_ASAP7_75t_L g3042 ( 
.A(n_2859),
.B(n_2504),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2883),
.B(n_2651),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2885),
.B(n_2615),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2768),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2812),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_2959),
.A2(n_2656),
.B1(n_2589),
.B2(n_2548),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2856),
.B(n_2549),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2914),
.B(n_2652),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2906),
.B(n_2455),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2776),
.B(n_2485),
.Y(n_3051)
);

AND2x6_ASAP7_75t_SL g3052 ( 
.A(n_2809),
.B(n_2849),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2813),
.B(n_2655),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2917),
.B(n_2899),
.Y(n_3054)
);

OR2x6_ASAP7_75t_L g3055 ( 
.A(n_2981),
.B(n_2482),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2817),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2825),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2793),
.Y(n_3058)
);

INVxp67_ASAP7_75t_SL g3059 ( 
.A(n_2744),
.Y(n_3059)
);

BUFx2_ASAP7_75t_L g3060 ( 
.A(n_2780),
.Y(n_3060)
);

NOR3xp33_ASAP7_75t_L g3061 ( 
.A(n_2907),
.B(n_1259),
.C(n_1257),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2844),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2848),
.B(n_2524),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2852),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2747),
.B(n_2491),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_SL g3066 ( 
.A(n_2887),
.B(n_2545),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2802),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2786),
.B(n_2673),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2807),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2818),
.Y(n_3070)
);

INVx1_ASAP7_75t_SL g3071 ( 
.A(n_2808),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2855),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2857),
.B(n_2553),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2794),
.B(n_2763),
.Y(n_3074)
);

AOI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2751),
.A2(n_2565),
.B1(n_2569),
.B2(n_2649),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2861),
.A2(n_1408),
.B1(n_1450),
.B2(n_1326),
.Y(n_3076)
);

CKINVDCx5p33_ASAP7_75t_R g3077 ( 
.A(n_2958),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_2880),
.B(n_2482),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2937),
.B(n_2675),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2858),
.B(n_2558),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2862),
.B(n_2559),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2874),
.B(n_2811),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2969),
.B(n_1078),
.Y(n_3083)
);

BUFx6f_ASAP7_75t_SL g3084 ( 
.A(n_2759),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2945),
.B(n_2580),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_2973),
.B(n_2685),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2821),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2976),
.B(n_2797),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2945),
.B(n_2640),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_2801),
.B(n_2837),
.Y(n_3090)
);

O2A1O1Ixp33_ASAP7_75t_L g3091 ( 
.A1(n_2952),
.A2(n_1266),
.B(n_1273),
.C(n_1269),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2839),
.B(n_1408),
.Y(n_3092)
);

OAI221xp5_ASAP7_75t_L g3093 ( 
.A1(n_2986),
.A2(n_1294),
.B1(n_1296),
.B2(n_1289),
.C(n_1283),
.Y(n_3093)
);

OAI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_2894),
.A2(n_1080),
.B1(n_1082),
.B2(n_1079),
.Y(n_3094)
);

INVxp33_ASAP7_75t_L g3095 ( 
.A(n_2796),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2834),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_L g3097 ( 
.A(n_2980),
.B(n_1084),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2945),
.B(n_2685),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2828),
.B(n_2685),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_SL g3100 ( 
.A(n_2873),
.B(n_2875),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2984),
.B(n_1408),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2828),
.B(n_1271),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_2896),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2877),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_SL g3105 ( 
.A(n_2978),
.B(n_2543),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2892),
.B(n_1088),
.Y(n_3106)
);

OAI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2819),
.A2(n_1096),
.B1(n_1098),
.B2(n_1095),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2878),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2828),
.B(n_2822),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2886),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_2803),
.A2(n_1509),
.B1(n_1644),
.B2(n_1450),
.Y(n_3111)
);

HB1xp67_ASAP7_75t_L g3112 ( 
.A(n_2902),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2890),
.B(n_2891),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2908),
.B(n_1290),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2912),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2895),
.B(n_1102),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2923),
.B(n_1336),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2924),
.Y(n_3118)
);

NAND2xp33_ASAP7_75t_L g3119 ( 
.A(n_2971),
.B(n_1105),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2823),
.Y(n_3120)
);

AOI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_2888),
.A2(n_1509),
.B1(n_1644),
.B2(n_1450),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2925),
.B(n_1400),
.Y(n_3122)
);

AOI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_2752),
.A2(n_2596),
.B1(n_1107),
.B2(n_1109),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2791),
.A2(n_1437),
.B(n_1400),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2926),
.B(n_1437),
.Y(n_3125)
);

INVx3_ASAP7_75t_L g3126 ( 
.A(n_2755),
.Y(n_3126)
);

INVx2_ASAP7_75t_SL g3127 ( 
.A(n_2913),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_2903),
.B(n_1106),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2833),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2927),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2905),
.B(n_1115),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2935),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2942),
.B(n_1460),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_2910),
.B(n_1125),
.Y(n_3134)
);

A2O1A1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_2909),
.A2(n_1302),
.B(n_1303),
.C(n_1297),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2951),
.B(n_1127),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2841),
.B(n_1129),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2841),
.B(n_1131),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2865),
.B(n_1133),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_2956),
.B(n_2568),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2868),
.B(n_1460),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2865),
.B(n_1136),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_2882),
.B(n_1139),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2847),
.Y(n_3144)
);

NAND3xp33_ASAP7_75t_L g3145 ( 
.A(n_2757),
.B(n_1142),
.C(n_1140),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2868),
.B(n_1481),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2868),
.B(n_1481),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2851),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2850),
.B(n_1482),
.Y(n_3149)
);

BUFx3_ASAP7_75t_L g3150 ( 
.A(n_2765),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_2775),
.B(n_1143),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2850),
.B(n_2845),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2929),
.B(n_1509),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2773),
.B(n_1147),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2948),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2889),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2777),
.B(n_1150),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_2779),
.B(n_1151),
.Y(n_3158)
);

INVx8_ASAP7_75t_L g3159 ( 
.A(n_2850),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2918),
.B(n_1152),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2893),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_2765),
.Y(n_3162)
);

BUFx8_ASAP7_75t_L g3163 ( 
.A(n_2970),
.Y(n_3163)
);

BUFx12f_ASAP7_75t_L g3164 ( 
.A(n_2934),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2897),
.B(n_1482),
.Y(n_3165)
);

OAI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2911),
.A2(n_2799),
.B(n_2967),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2957),
.A2(n_1521),
.B(n_1519),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2898),
.B(n_1519),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2904),
.B(n_1521),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2922),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2778),
.B(n_1154),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2928),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_2778),
.B(n_1161),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2936),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2939),
.B(n_1545),
.Y(n_3175)
);

OR2x6_ASAP7_75t_L g3176 ( 
.A(n_2805),
.B(n_1545),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2944),
.B(n_2955),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2836),
.B(n_1166),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2866),
.B(n_1580),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2838),
.B(n_1580),
.Y(n_3180)
);

A2O1A1Ixp33_ASAP7_75t_L g3181 ( 
.A1(n_2827),
.A2(n_1321),
.B(n_1328),
.C(n_1315),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2854),
.B(n_1589),
.Y(n_3182)
);

AOI22xp5_ASAP7_75t_L g3183 ( 
.A1(n_2835),
.A2(n_1169),
.B1(n_1172),
.B2(n_1170),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2767),
.Y(n_3184)
);

NOR2xp67_ASAP7_75t_SL g3185 ( 
.A(n_2815),
.B(n_1173),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2790),
.B(n_1589),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2826),
.B(n_1607),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2879),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_SL g3189 ( 
.A(n_2826),
.B(n_1174),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_3155),
.Y(n_3190)
);

OAI22xp5_ASAP7_75t_L g3191 ( 
.A1(n_3014),
.A2(n_2900),
.B1(n_2943),
.B2(n_2941),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3113),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_3015),
.B(n_2824),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2988),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2995),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2992),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2997),
.Y(n_3197)
);

AOI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_3053),
.A2(n_2966),
.B(n_2961),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2991),
.B(n_2990),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3004),
.Y(n_3200)
);

A2O1A1Ixp33_ASAP7_75t_L g3201 ( 
.A1(n_3010),
.A2(n_2989),
.B(n_3007),
.C(n_3082),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2987),
.B(n_2962),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_3024),
.A2(n_2963),
.B(n_2960),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_3063),
.A2(n_2974),
.B(n_2968),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_3028),
.Y(n_3205)
);

INVx11_ASAP7_75t_L g3206 ( 
.A(n_3035),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_3054),
.B(n_2884),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3008),
.B(n_2829),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3016),
.B(n_2829),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_2994),
.B(n_2824),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3096),
.B(n_2831),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_3073),
.A2(n_2820),
.B(n_2814),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_3045),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_3013),
.B(n_2831),
.Y(n_3214)
);

INVx2_ASAP7_75t_SL g3215 ( 
.A(n_3009),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3018),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_3033),
.B(n_2810),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_3041),
.B(n_2964),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_3030),
.B(n_2940),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_3036),
.B(n_2938),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_3006),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3022),
.B(n_2983),
.Y(n_3222)
);

AOI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_3080),
.A2(n_2846),
.B(n_2842),
.Y(n_3223)
);

A2O1A1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_3091),
.A2(n_2864),
.B(n_2979),
.C(n_2975),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_3017),
.B(n_2972),
.Y(n_3225)
);

AOI21x1_ASAP7_75t_L g3226 ( 
.A1(n_3166),
.A2(n_2977),
.B(n_2120),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_3127),
.B(n_2915),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3068),
.A2(n_2792),
.B1(n_2965),
.B2(n_2800),
.Y(n_3228)
);

AOI22xp5_ASAP7_75t_L g3229 ( 
.A1(n_3044),
.A2(n_2787),
.B1(n_2792),
.B2(n_2860),
.Y(n_3229)
);

INVx3_ASAP7_75t_L g3230 ( 
.A(n_3006),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3021),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_3025),
.A2(n_2783),
.B1(n_2971),
.B2(n_2853),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_SL g3233 ( 
.A(n_3049),
.B(n_2832),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_3081),
.A2(n_2853),
.B(n_2832),
.Y(n_3234)
);

CKINVDCx20_ASAP7_75t_R g3235 ( 
.A(n_3011),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_3058),
.Y(n_3236)
);

INVx3_ASAP7_75t_L g3237 ( 
.A(n_3164),
.Y(n_3237)
);

O2A1O1Ixp33_ASAP7_75t_L g3238 ( 
.A1(n_3066),
.A2(n_1330),
.B(n_1337),
.C(n_1335),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_L g3239 ( 
.A(n_3032),
.B(n_2863),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3067),
.Y(n_3240)
);

AO21x1_ASAP7_75t_L g3241 ( 
.A1(n_3109),
.A2(n_1349),
.B(n_1340),
.Y(n_3241)
);

OAI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3188),
.A2(n_1358),
.B(n_1353),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3026),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3029),
.A2(n_2876),
.B(n_2863),
.Y(n_3244)
);

OAI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_3135),
.A2(n_3108),
.B(n_3104),
.Y(n_3245)
);

OAI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_3110),
.A2(n_1361),
.B(n_1360),
.Y(n_3246)
);

INVx3_ASAP7_75t_L g3247 ( 
.A(n_3162),
.Y(n_3247)
);

OAI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3115),
.A2(n_1365),
.B(n_1362),
.Y(n_3248)
);

AO21x1_ASAP7_75t_L g3249 ( 
.A1(n_3075),
.A2(n_1376),
.B(n_1371),
.Y(n_3249)
);

O2A1O1Ixp33_ASAP7_75t_L g3250 ( 
.A1(n_3061),
.A2(n_1377),
.B(n_1385),
.C(n_1382),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_3065),
.B(n_3074),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3143),
.B(n_2876),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3046),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3037),
.A2(n_2954),
.B(n_2947),
.Y(n_3254)
);

OAI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3118),
.A2(n_1391),
.B(n_1390),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_3038),
.B(n_2947),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3056),
.B(n_2954),
.Y(n_3257)
);

CKINVDCx10_ASAP7_75t_R g3258 ( 
.A(n_2996),
.Y(n_3258)
);

AO21x1_ASAP7_75t_L g3259 ( 
.A1(n_3039),
.A2(n_1402),
.B(n_1394),
.Y(n_3259)
);

OAI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3130),
.A2(n_1409),
.B(n_1403),
.Y(n_3260)
);

INVx2_ASAP7_75t_SL g3261 ( 
.A(n_3077),
.Y(n_3261)
);

BUFx6f_ASAP7_75t_L g3262 ( 
.A(n_3162),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3020),
.A2(n_1647),
.B(n_1607),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3057),
.Y(n_3264)
);

O2A1O1Ixp5_ASAP7_75t_L g3265 ( 
.A1(n_3171),
.A2(n_1766),
.B(n_1649),
.C(n_1664),
.Y(n_3265)
);

NAND2xp33_ASAP7_75t_L g3266 ( 
.A(n_3031),
.B(n_2985),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_3062),
.A2(n_1649),
.B(n_1647),
.Y(n_3267)
);

INVxp67_ASAP7_75t_L g3268 ( 
.A(n_2999),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3064),
.B(n_1175),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3092),
.B(n_2953),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3072),
.B(n_1176),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_3095),
.B(n_1177),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3101),
.B(n_1179),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3132),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_3071),
.B(n_1180),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3083),
.B(n_1181),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3153),
.B(n_1644),
.Y(n_3277)
);

AND2x4_ASAP7_75t_L g3278 ( 
.A(n_3150),
.B(n_2901),
.Y(n_3278)
);

AOI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_3152),
.A2(n_1692),
.B(n_1664),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3069),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3106),
.B(n_1182),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3001),
.Y(n_3282)
);

O2A1O1Ixp33_ASAP7_75t_L g3283 ( 
.A1(n_3094),
.A2(n_1412),
.B(n_1418),
.C(n_1415),
.Y(n_3283)
);

OAI22xp5_ASAP7_75t_L g3284 ( 
.A1(n_3059),
.A2(n_1186),
.B1(n_1190),
.B2(n_1187),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_3055),
.Y(n_3285)
);

A2O1A1Ixp33_ASAP7_75t_L g3286 ( 
.A1(n_3178),
.A2(n_1702),
.B(n_1766),
.C(n_1692),
.Y(n_3286)
);

NAND2x1p5_ASAP7_75t_L g3287 ( 
.A(n_3000),
.B(n_2110),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_3070),
.Y(n_3288)
);

NOR3xp33_ASAP7_75t_L g3289 ( 
.A(n_3005),
.B(n_1424),
.C(n_1422),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_3085),
.A2(n_1814),
.B(n_1702),
.Y(n_3290)
);

CKINVDCx11_ASAP7_75t_R g3291 ( 
.A(n_3052),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_3055),
.Y(n_3292)
);

AOI21x1_ASAP7_75t_L g3293 ( 
.A1(n_3114),
.A2(n_2126),
.B(n_2125),
.Y(n_3293)
);

AND2x4_ASAP7_75t_L g3294 ( 
.A(n_3078),
.B(n_1429),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3043),
.A2(n_1859),
.B(n_1814),
.Y(n_3295)
);

OAI22xp5_ASAP7_75t_L g3296 ( 
.A1(n_3183),
.A2(n_1191),
.B1(n_1194),
.B2(n_1192),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3177),
.A2(n_1859),
.B(n_1433),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3186),
.B(n_1195),
.Y(n_3298)
);

BUFx6f_ASAP7_75t_L g3299 ( 
.A(n_3034),
.Y(n_3299)
);

AOI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_3012),
.A2(n_1434),
.B(n_1431),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3116),
.A2(n_1442),
.B(n_1440),
.Y(n_3301)
);

BUFx6f_ASAP7_75t_L g3302 ( 
.A(n_2993),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_3019),
.B(n_1196),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3159),
.B(n_1197),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3159),
.B(n_3097),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3128),
.A2(n_1448),
.B(n_1444),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3154),
.B(n_1199),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3157),
.B(n_1201),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3158),
.B(n_1202),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_3048),
.B(n_1203),
.Y(n_3310)
);

AOI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_3131),
.A2(n_3136),
.B(n_3134),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3126),
.A2(n_1206),
.B1(n_1208),
.B2(n_1207),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3117),
.B(n_1212),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_L g3314 ( 
.A(n_3060),
.B(n_1216),
.Y(n_3314)
);

INVx11_ASAP7_75t_L g3315 ( 
.A(n_3163),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3165),
.Y(n_3316)
);

OAI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_3179),
.A2(n_1461),
.B(n_1452),
.Y(n_3317)
);

INVx2_ASAP7_75t_SL g3318 ( 
.A(n_3103),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3003),
.A2(n_2998),
.B(n_3151),
.Y(n_3319)
);

NOR2xp33_ASAP7_75t_L g3320 ( 
.A(n_3042),
.B(n_1218),
.Y(n_3320)
);

OAI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3124),
.A2(n_1465),
.B(n_1464),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3184),
.A2(n_1219),
.B1(n_1223),
.B2(n_1220),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3122),
.B(n_1224),
.Y(n_3323)
);

HB1xp67_ASAP7_75t_L g3324 ( 
.A(n_3112),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3090),
.A2(n_1479),
.B(n_1475),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_SL g3326 ( 
.A(n_3079),
.B(n_1230),
.Y(n_3326)
);

OAI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3167),
.A2(n_1484),
.B(n_1483),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3125),
.B(n_1231),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3161),
.B(n_1232),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3051),
.B(n_3160),
.Y(n_3330)
);

O2A1O1Ixp33_ASAP7_75t_L g3331 ( 
.A1(n_3107),
.A2(n_1486),
.B(n_1495),
.C(n_1492),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_SL g3332 ( 
.A(n_3050),
.B(n_1233),
.Y(n_3332)
);

INVx4_ASAP7_75t_L g3333 ( 
.A(n_3040),
.Y(n_3333)
);

HB1xp67_ASAP7_75t_L g3334 ( 
.A(n_3176),
.Y(n_3334)
);

INVxp67_ASAP7_75t_L g3335 ( 
.A(n_3187),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3002),
.B(n_1234),
.Y(n_3336)
);

AOI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_3111),
.A2(n_1236),
.B1(n_1239),
.B2(n_1237),
.Y(n_3337)
);

AOI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_3100),
.A2(n_1514),
.B(n_1507),
.Y(n_3338)
);

O2A1O1Ixp33_ASAP7_75t_L g3339 ( 
.A1(n_3173),
.A2(n_1518),
.B(n_1527),
.C(n_1524),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3168),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3087),
.B(n_1241),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3190),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3196),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3200),
.Y(n_3344)
);

OAI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_3201),
.A2(n_3121),
.B1(n_3076),
.B2(n_3145),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3281),
.A2(n_3176),
.B1(n_3088),
.B2(n_3023),
.Y(n_3346)
);

BUFx2_ASAP7_75t_L g3347 ( 
.A(n_3324),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3216),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3231),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3243),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3266),
.A2(n_3198),
.B(n_3223),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3199),
.B(n_3047),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_R g3353 ( 
.A(n_3235),
.B(n_3084),
.Y(n_3353)
);

INVx5_ASAP7_75t_L g3354 ( 
.A(n_3221),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_3276),
.A2(n_3123),
.B1(n_3189),
.B2(n_3181),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_L g3356 ( 
.A(n_3202),
.B(n_3027),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3222),
.A2(n_3093),
.B1(n_3129),
.B2(n_3120),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3253),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_3193),
.B(n_3140),
.Y(n_3359)
);

INVxp67_ASAP7_75t_L g3360 ( 
.A(n_3282),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_R g3361 ( 
.A(n_3258),
.B(n_3105),
.Y(n_3361)
);

A2O1A1Ixp33_ASAP7_75t_L g3362 ( 
.A1(n_3217),
.A2(n_3141),
.B(n_3147),
.C(n_3146),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_3283),
.A2(n_3149),
.B(n_3102),
.C(n_3089),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_3251),
.B(n_3330),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3192),
.B(n_3144),
.Y(n_3365)
);

CKINVDCx5p33_ASAP7_75t_R g3366 ( 
.A(n_3206),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3194),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_3221),
.Y(n_3368)
);

NOR3xp33_ASAP7_75t_SL g3369 ( 
.A(n_3326),
.B(n_3138),
.C(n_3137),
.Y(n_3369)
);

OAI21xp33_ASAP7_75t_L g3370 ( 
.A1(n_3307),
.A2(n_3185),
.B(n_1292),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_SL g3371 ( 
.A(n_3218),
.B(n_3209),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3225),
.B(n_3148),
.Y(n_3372)
);

NOR2x1p5_ASAP7_75t_L g3373 ( 
.A(n_3237),
.B(n_3099),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3228),
.A2(n_3156),
.B1(n_3172),
.B2(n_3170),
.Y(n_3374)
);

NOR3xp33_ASAP7_75t_SL g3375 ( 
.A(n_3311),
.B(n_3142),
.C(n_3139),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3308),
.A2(n_3133),
.B1(n_3182),
.B2(n_3180),
.Y(n_3376)
);

AOI21xp5_ASAP7_75t_L g3377 ( 
.A1(n_3204),
.A2(n_3119),
.B(n_3098),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_SL g3378 ( 
.A(n_3333),
.B(n_3174),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_3210),
.B(n_3086),
.Y(n_3379)
);

NAND3xp33_ASAP7_75t_L g3380 ( 
.A(n_3309),
.B(n_1247),
.C(n_1244),
.Y(n_3380)
);

INVx4_ASAP7_75t_L g3381 ( 
.A(n_3315),
.Y(n_3381)
);

BUFx2_ASAP7_75t_L g3382 ( 
.A(n_3247),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3195),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3197),
.Y(n_3384)
);

BUFx2_ASAP7_75t_L g3385 ( 
.A(n_3285),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_3203),
.A2(n_3175),
.B(n_3169),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3205),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3264),
.Y(n_3388)
);

O2A1O1Ixp33_ASAP7_75t_SL g3389 ( 
.A1(n_3191),
.A2(n_1534),
.B(n_1536),
.C(n_1529),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3310),
.B(n_3031),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3212),
.A2(n_3031),
.B(n_1540),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_3213),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_3291),
.Y(n_3393)
);

INVx3_ASAP7_75t_L g3394 ( 
.A(n_3262),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3277),
.B(n_3031),
.Y(n_3395)
);

CKINVDCx14_ASAP7_75t_R g3396 ( 
.A(n_3278),
.Y(n_3396)
);

BUFx6f_ASAP7_75t_L g3397 ( 
.A(n_3285),
.Y(n_3397)
);

NAND3xp33_ASAP7_75t_L g3398 ( 
.A(n_3320),
.B(n_1254),
.C(n_1249),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_SL g3399 ( 
.A(n_3252),
.B(n_1748),
.Y(n_3399)
);

BUFx6f_ASAP7_75t_L g3400 ( 
.A(n_3292),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3274),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3245),
.A2(n_1541),
.B(n_1539),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3233),
.A2(n_1554),
.B(n_1544),
.Y(n_3403)
);

BUFx6f_ASAP7_75t_L g3404 ( 
.A(n_3292),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_3242),
.A2(n_1557),
.B(n_1561),
.C(n_1555),
.Y(n_3405)
);

O2A1O1Ixp33_ASAP7_75t_L g3406 ( 
.A1(n_3331),
.A2(n_1573),
.B(n_1578),
.C(n_1576),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3236),
.Y(n_3407)
);

HB1xp67_ASAP7_75t_L g3408 ( 
.A(n_3268),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3234),
.A2(n_1596),
.B(n_1588),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3256),
.B(n_1262),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3270),
.B(n_1748),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3240),
.Y(n_3412)
);

OAI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_3246),
.A2(n_1601),
.B(n_1597),
.Y(n_3413)
);

BUFx8_ASAP7_75t_L g3414 ( 
.A(n_3220),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3280),
.Y(n_3415)
);

AND2x2_ASAP7_75t_L g3416 ( 
.A(n_3314),
.B(n_1748),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_3239),
.B(n_1797),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3288),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3257),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3219),
.B(n_1267),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3211),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3248),
.B(n_1272),
.Y(n_3422)
);

O2A1O1Ixp33_ASAP7_75t_L g3423 ( 
.A1(n_3250),
.A2(n_1602),
.B(n_1608),
.C(n_1606),
.Y(n_3423)
);

A2O1A1Ixp33_ASAP7_75t_L g3424 ( 
.A1(n_3255),
.A2(n_1617),
.B(n_1618),
.C(n_1615),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_3208),
.B(n_1797),
.Y(n_3425)
);

HB1xp67_ASAP7_75t_L g3426 ( 
.A(n_3318),
.Y(n_3426)
);

OAI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3229),
.A2(n_1277),
.B1(n_1285),
.B2(n_1282),
.Y(n_3427)
);

INVx2_ASAP7_75t_SL g3428 ( 
.A(n_3262),
.Y(n_3428)
);

O2A1O1Ixp33_ASAP7_75t_L g3429 ( 
.A1(n_3296),
.A2(n_1619),
.B(n_1631),
.C(n_1626),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3260),
.B(n_1288),
.Y(n_3430)
);

BUFx6f_ASAP7_75t_L g3431 ( 
.A(n_3302),
.Y(n_3431)
);

INVx3_ASAP7_75t_L g3432 ( 
.A(n_3302),
.Y(n_3432)
);

OA21x2_ASAP7_75t_L g3433 ( 
.A1(n_3226),
.A2(n_2136),
.B(n_1641),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_3207),
.B(n_1797),
.Y(n_3434)
);

INVx3_ASAP7_75t_L g3435 ( 
.A(n_3299),
.Y(n_3435)
);

CKINVDCx14_ASAP7_75t_R g3436 ( 
.A(n_3227),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3254),
.A2(n_3214),
.B(n_3244),
.Y(n_3437)
);

O2A1O1Ixp33_ASAP7_75t_L g3438 ( 
.A1(n_3273),
.A2(n_1640),
.B(n_1655),
.C(n_1651),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3215),
.B(n_1822),
.Y(n_3439)
);

O2A1O1Ixp33_ASAP7_75t_L g3440 ( 
.A1(n_3286),
.A2(n_1658),
.B(n_1662),
.C(n_1661),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3335),
.B(n_1293),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_3230),
.Y(n_3442)
);

O2A1O1Ixp33_ASAP7_75t_L g3443 ( 
.A1(n_3238),
.A2(n_1663),
.B(n_1669),
.C(n_1665),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3224),
.A2(n_1676),
.B(n_1673),
.Y(n_3444)
);

OAI21x1_ASAP7_75t_L g3445 ( 
.A1(n_3293),
.A2(n_1679),
.B(n_1677),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3232),
.A2(n_1690),
.B(n_1688),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_3261),
.B(n_1822),
.Y(n_3447)
);

A2O1A1Ixp33_ASAP7_75t_SL g3448 ( 
.A1(n_3319),
.A2(n_1708),
.B(n_1719),
.C(n_1706),
.Y(n_3448)
);

AND2x4_ASAP7_75t_L g3449 ( 
.A(n_3299),
.B(n_1722),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3316),
.A2(n_1725),
.B(n_1724),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3305),
.B(n_1298),
.Y(n_3451)
);

INVx4_ASAP7_75t_L g3452 ( 
.A(n_3294),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_L g3453 ( 
.A(n_3332),
.B(n_1300),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3269),
.A2(n_1305),
.B1(n_1306),
.B2(n_1301),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3340),
.Y(n_3455)
);

AOI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3313),
.A2(n_1728),
.B(n_1726),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3334),
.B(n_1822),
.Y(n_3457)
);

O2A1O1Ixp33_ASAP7_75t_L g3458 ( 
.A1(n_3323),
.A2(n_1729),
.B(n_1745),
.C(n_1740),
.Y(n_3458)
);

HB1xp67_ASAP7_75t_L g3459 ( 
.A(n_3272),
.Y(n_3459)
);

CKINVDCx20_ASAP7_75t_R g3460 ( 
.A(n_3275),
.Y(n_3460)
);

BUFx4f_ASAP7_75t_SL g3461 ( 
.A(n_3303),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3328),
.A2(n_1752),
.B(n_1747),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3317),
.B(n_1308),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_R g3464 ( 
.A(n_3304),
.B(n_1828),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3336),
.A2(n_1757),
.B(n_1754),
.Y(n_3465)
);

OAI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_3271),
.A2(n_1312),
.B1(n_1313),
.B2(n_1310),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_SL g3467 ( 
.A1(n_3300),
.A2(n_1828),
.B1(n_1764),
.B2(n_1765),
.Y(n_3467)
);

O2A1O1Ixp33_ASAP7_75t_L g3468 ( 
.A1(n_3289),
.A2(n_1758),
.B(n_1770),
.C(n_1769),
.Y(n_3468)
);

AOI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3290),
.A2(n_1773),
.B(n_1771),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3341),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3279),
.Y(n_3471)
);

A2O1A1Ixp33_ASAP7_75t_L g3472 ( 
.A1(n_3263),
.A2(n_1780),
.B(n_1781),
.C(n_1777),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3329),
.Y(n_3473)
);

A2O1A1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3327),
.A2(n_1784),
.B(n_1789),
.C(n_1783),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3298),
.B(n_1314),
.Y(n_3475)
);

O2A1O1Ixp33_ASAP7_75t_L g3476 ( 
.A1(n_3339),
.A2(n_3284),
.B(n_3322),
.C(n_3312),
.Y(n_3476)
);

AOI22xp33_ASAP7_75t_L g3477 ( 
.A1(n_3249),
.A2(n_1828),
.B1(n_1319),
.B2(n_1324),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3265),
.Y(n_3478)
);

NOR2x1_ASAP7_75t_L g3479 ( 
.A(n_3321),
.B(n_3295),
.Y(n_3479)
);

OR2x2_ASAP7_75t_L g3480 ( 
.A(n_3287),
.B(n_1791),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3241),
.B(n_1317),
.Y(n_3481)
);

O2A1O1Ixp33_ASAP7_75t_SL g3482 ( 
.A1(n_3390),
.A2(n_1803),
.B(n_1804),
.C(n_1800),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3351),
.A2(n_3259),
.B(n_3297),
.Y(n_3483)
);

NAND2x1p5_ASAP7_75t_L g3484 ( 
.A(n_3354),
.B(n_3325),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3343),
.Y(n_3485)
);

BUFx6f_ASAP7_75t_L g3486 ( 
.A(n_3397),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3342),
.Y(n_3487)
);

CKINVDCx20_ASAP7_75t_R g3488 ( 
.A(n_3361),
.Y(n_3488)
);

OAI21x1_ASAP7_75t_L g3489 ( 
.A1(n_3445),
.A2(n_3386),
.B(n_3437),
.Y(n_3489)
);

OAI21x1_ASAP7_75t_L g3490 ( 
.A1(n_3471),
.A2(n_3267),
.B(n_3301),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3364),
.B(n_3352),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3371),
.B(n_3338),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3459),
.B(n_3306),
.Y(n_3493)
);

OAI21x1_ASAP7_75t_L g3494 ( 
.A1(n_3377),
.A2(n_1811),
.B(n_1809),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3344),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3391),
.A2(n_3395),
.B(n_3389),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3448),
.A2(n_1816),
.B(n_1813),
.Y(n_3497)
);

NAND2x1p5_ASAP7_75t_L g3498 ( 
.A(n_3354),
.B(n_3368),
.Y(n_3498)
);

AND2x4_ASAP7_75t_L g3499 ( 
.A(n_3452),
.B(n_3337),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3367),
.Y(n_3500)
);

OAI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3420),
.A2(n_3398),
.B(n_3422),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3379),
.B(n_3362),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_3356),
.B(n_1325),
.Y(n_3503)
);

INVxp67_ASAP7_75t_L g3504 ( 
.A(n_3426),
.Y(n_3504)
);

OAI21x1_ASAP7_75t_L g3505 ( 
.A1(n_3433),
.A2(n_1821),
.B(n_1819),
.Y(n_3505)
);

AO21x1_ASAP7_75t_L g3506 ( 
.A1(n_3402),
.A2(n_1837),
.B(n_1824),
.Y(n_3506)
);

INVx1_ASAP7_75t_SL g3507 ( 
.A(n_3359),
.Y(n_3507)
);

INVxp67_ASAP7_75t_SL g3508 ( 
.A(n_3360),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3354),
.B(n_1838),
.Y(n_3509)
);

OAI21x1_ASAP7_75t_L g3510 ( 
.A1(n_3433),
.A2(n_1844),
.B(n_1839),
.Y(n_3510)
);

AOI211x1_ASAP7_75t_L g3511 ( 
.A1(n_3427),
.A2(n_1852),
.B(n_1857),
.C(n_1855),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_SL g3512 ( 
.A1(n_3363),
.A2(n_1320),
.B(n_1278),
.Y(n_3512)
);

OAI21x1_ASAP7_75t_SL g3513 ( 
.A1(n_3476),
.A2(n_1862),
.B(n_1858),
.Y(n_3513)
);

AO31x2_ASAP7_75t_L g3514 ( 
.A1(n_3478),
.A2(n_1863),
.A3(n_1880),
.B(n_1876),
.Y(n_3514)
);

OAI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3430),
.A2(n_1882),
.B(n_1354),
.Y(n_3515)
);

NAND2x1p5_ASAP7_75t_L g3516 ( 
.A(n_3368),
.B(n_2300),
.Y(n_3516)
);

BUFx6f_ASAP7_75t_L g3517 ( 
.A(n_3397),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3479),
.A2(n_1347),
.B(n_1320),
.Y(n_3518)
);

OAI21x1_ASAP7_75t_SL g3519 ( 
.A1(n_3413),
.A2(n_1111),
.B(n_0),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3348),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3473),
.B(n_1331),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3372),
.B(n_3408),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3349),
.Y(n_3523)
);

NAND2x1p5_ASAP7_75t_L g3524 ( 
.A(n_3400),
.B(n_2300),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3346),
.B(n_1332),
.Y(n_3525)
);

OAI21x1_ASAP7_75t_L g3526 ( 
.A1(n_3444),
.A2(n_951),
.B(n_949),
.Y(n_3526)
);

NOR3xp33_ASAP7_75t_L g3527 ( 
.A(n_3345),
.B(n_1338),
.C(n_1334),
.Y(n_3527)
);

HB1xp67_ASAP7_75t_L g3528 ( 
.A(n_3347),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3376),
.A2(n_3370),
.B(n_3355),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3470),
.B(n_1339),
.Y(n_3530)
);

AO31x2_ASAP7_75t_L g3531 ( 
.A1(n_3455),
.A2(n_3384),
.A3(n_3387),
.B(n_3383),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3350),
.Y(n_3532)
);

CKINVDCx16_ASAP7_75t_R g3533 ( 
.A(n_3353),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3421),
.B(n_1341),
.Y(n_3534)
);

CKINVDCx20_ASAP7_75t_R g3535 ( 
.A(n_3366),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3481),
.A2(n_1347),
.B(n_1320),
.Y(n_3536)
);

BUFx4f_ASAP7_75t_SL g3537 ( 
.A(n_3381),
.Y(n_3537)
);

AOI21x1_ASAP7_75t_L g3538 ( 
.A1(n_3446),
.A2(n_2306),
.B(n_2304),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3358),
.Y(n_3539)
);

CKINVDCx6p67_ASAP7_75t_R g3540 ( 
.A(n_3442),
.Y(n_3540)
);

OA21x2_ASAP7_75t_L g3541 ( 
.A1(n_3409),
.A2(n_1344),
.B(n_1343),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3392),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3419),
.B(n_1350),
.Y(n_3543)
);

AOI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3365),
.A2(n_1347),
.B(n_1320),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3407),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3378),
.B(n_1352),
.Y(n_3546)
);

NOR2xp67_ASAP7_75t_L g3547 ( 
.A(n_3435),
.B(n_3428),
.Y(n_3547)
);

OAI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_3463),
.A2(n_3410),
.B(n_3429),
.Y(n_3548)
);

NAND3xp33_ASAP7_75t_L g3549 ( 
.A(n_3458),
.B(n_1364),
.C(n_1363),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3380),
.A2(n_1410),
.B(n_1347),
.Y(n_3550)
);

BUFx8_ASAP7_75t_L g3551 ( 
.A(n_3431),
.Y(n_3551)
);

OAI21x1_ASAP7_75t_L g3552 ( 
.A1(n_3388),
.A2(n_953),
.B(n_952),
.Y(n_3552)
);

NOR2xp67_ASAP7_75t_L g3553 ( 
.A(n_3394),
.B(n_955),
.Y(n_3553)
);

OAI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3475),
.A2(n_1395),
.B(n_1374),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3401),
.B(n_1366),
.Y(n_3555)
);

OAI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3406),
.A2(n_1405),
.B(n_1380),
.Y(n_3556)
);

INVx3_ASAP7_75t_SL g3557 ( 
.A(n_3393),
.Y(n_3557)
);

AOI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3417),
.A2(n_3399),
.B(n_3425),
.Y(n_3558)
);

A2O1A1Ixp33_ASAP7_75t_L g3559 ( 
.A1(n_3438),
.A2(n_1372),
.B(n_1378),
.C(n_1370),
.Y(n_3559)
);

INVxp33_ASAP7_75t_SL g3560 ( 
.A(n_3464),
.Y(n_3560)
);

OAI21x1_ASAP7_75t_L g3561 ( 
.A1(n_3469),
.A2(n_959),
.B(n_956),
.Y(n_3561)
);

AO31x2_ASAP7_75t_L g3562 ( 
.A1(n_3412),
.A2(n_963),
.A3(n_964),
.B(n_960),
.Y(n_3562)
);

OAI21x1_ASAP7_75t_L g3563 ( 
.A1(n_3403),
.A2(n_970),
.B(n_966),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3415),
.Y(n_3564)
);

OR2x2_ASAP7_75t_L g3565 ( 
.A(n_3385),
.B(n_1410),
.Y(n_3565)
);

AOI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3434),
.A2(n_1435),
.B(n_1410),
.Y(n_3566)
);

A2O1A1Ixp33_ASAP7_75t_L g3567 ( 
.A1(n_3443),
.A2(n_1388),
.B(n_1389),
.C(n_1384),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_3369),
.B(n_1392),
.Y(n_3568)
);

AOI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3465),
.A2(n_2306),
.B(n_2304),
.Y(n_3569)
);

OAI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3405),
.A2(n_1423),
.B(n_1399),
.Y(n_3570)
);

INVx2_ASAP7_75t_SL g3571 ( 
.A(n_3414),
.Y(n_3571)
);

AOI221x1_ASAP7_75t_L g3572 ( 
.A1(n_3474),
.A2(n_1560),
.B1(n_1646),
.B2(n_1435),
.C(n_1410),
.Y(n_3572)
);

OR2x2_ASAP7_75t_L g3573 ( 
.A(n_3418),
.B(n_1435),
.Y(n_3573)
);

INVx2_ASAP7_75t_SL g3574 ( 
.A(n_3431),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3440),
.A2(n_1560),
.B(n_1435),
.Y(n_3575)
);

OAI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3451),
.A2(n_1428),
.B(n_1406),
.Y(n_3576)
);

OAI22x1_ASAP7_75t_L g3577 ( 
.A1(n_3416),
.A2(n_1396),
.B1(n_1407),
.B2(n_1393),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3375),
.B(n_1411),
.Y(n_3578)
);

OAI21x1_ASAP7_75t_L g3579 ( 
.A1(n_3373),
.A2(n_972),
.B(n_971),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3411),
.B(n_1413),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3382),
.B(n_3400),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3480),
.Y(n_3582)
);

AND2x4_ASAP7_75t_L g3583 ( 
.A(n_3404),
.B(n_3432),
.Y(n_3583)
);

INVxp67_ASAP7_75t_SL g3584 ( 
.A(n_3357),
.Y(n_3584)
);

BUFx6f_ASAP7_75t_L g3585 ( 
.A(n_3404),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3374),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3449),
.B(n_1419),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3424),
.B(n_1420),
.Y(n_3588)
);

OAI21x1_ASAP7_75t_L g3589 ( 
.A1(n_3450),
.A2(n_975),
.B(n_973),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3477),
.B(n_1425),
.Y(n_3590)
);

INVx3_ASAP7_75t_L g3591 ( 
.A(n_3461),
.Y(n_3591)
);

BUFx2_ASAP7_75t_L g3592 ( 
.A(n_3460),
.Y(n_3592)
);

AO31x2_ASAP7_75t_L g3593 ( 
.A1(n_3529),
.A2(n_3472),
.A3(n_3456),
.B(n_3462),
.Y(n_3593)
);

OAI21x1_ASAP7_75t_L g3594 ( 
.A1(n_3489),
.A2(n_3483),
.B(n_3518),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3491),
.B(n_3396),
.Y(n_3595)
);

AOI22xp33_ASAP7_75t_L g3596 ( 
.A1(n_3584),
.A2(n_3436),
.B1(n_3453),
.B2(n_3457),
.Y(n_3596)
);

INVx1_ASAP7_75t_SL g3597 ( 
.A(n_3507),
.Y(n_3597)
);

HB1xp67_ASAP7_75t_L g3598 ( 
.A(n_3528),
.Y(n_3598)
);

OA21x2_ASAP7_75t_L g3599 ( 
.A1(n_3544),
.A2(n_3502),
.B(n_3494),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3545),
.Y(n_3600)
);

O2A1O1Ixp33_ASAP7_75t_L g3601 ( 
.A1(n_3548),
.A2(n_3423),
.B(n_3468),
.C(n_3466),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3485),
.Y(n_3602)
);

NOR2xp33_ASAP7_75t_SL g3603 ( 
.A(n_3533),
.B(n_3441),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3495),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3487),
.Y(n_3605)
);

BUFx10_ASAP7_75t_L g3606 ( 
.A(n_3571),
.Y(n_3606)
);

OA21x2_ASAP7_75t_L g3607 ( 
.A1(n_3490),
.A2(n_3439),
.B(n_3447),
.Y(n_3607)
);

CKINVDCx11_ASAP7_75t_R g3608 ( 
.A(n_3488),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3522),
.B(n_1426),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3520),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3531),
.Y(n_3611)
);

BUFx3_ASAP7_75t_L g3612 ( 
.A(n_3551),
.Y(n_3612)
);

AOI221xp5_ASAP7_75t_L g3613 ( 
.A1(n_3515),
.A2(n_3454),
.B1(n_1438),
.B2(n_1439),
.C(n_1436),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3503),
.A2(n_3467),
.B1(n_1468),
.B2(n_1487),
.Y(n_3614)
);

O2A1O1Ixp33_ASAP7_75t_L g3615 ( 
.A1(n_3527),
.A2(n_1443),
.B(n_1447),
.C(n_1432),
.Y(n_3615)
);

AO21x2_ASAP7_75t_L g3616 ( 
.A1(n_3512),
.A2(n_2330),
.B(n_2324),
.Y(n_3616)
);

AOI22xp5_ASAP7_75t_L g3617 ( 
.A1(n_3525),
.A2(n_3499),
.B1(n_3577),
.B2(n_3560),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3586),
.A2(n_1646),
.B1(n_1659),
.B2(n_1560),
.Y(n_3618)
);

AO21x2_ASAP7_75t_L g3619 ( 
.A1(n_3505),
.A2(n_2330),
.B(n_2324),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3587),
.A2(n_1646),
.B1(n_1659),
.B2(n_1560),
.Y(n_3620)
);

O2A1O1Ixp33_ASAP7_75t_L g3621 ( 
.A1(n_3559),
.A2(n_1451),
.B(n_1454),
.C(n_1449),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3523),
.B(n_1),
.Y(n_3622)
);

NOR2x1_ASAP7_75t_R g3623 ( 
.A(n_3591),
.B(n_3592),
.Y(n_3623)
);

AOI22xp33_ASAP7_75t_L g3624 ( 
.A1(n_3582),
.A2(n_1659),
.B1(n_1733),
.B2(n_1646),
.Y(n_3624)
);

HB1xp67_ASAP7_75t_L g3625 ( 
.A(n_3508),
.Y(n_3625)
);

INVx6_ASAP7_75t_L g3626 ( 
.A(n_3486),
.Y(n_3626)
);

OAI21x1_ASAP7_75t_SL g3627 ( 
.A1(n_3513),
.A2(n_1),
.B(n_2),
.Y(n_3627)
);

OAI21x1_ASAP7_75t_L g3628 ( 
.A1(n_3496),
.A2(n_2333),
.B(n_2331),
.Y(n_3628)
);

AND2x4_ASAP7_75t_L g3629 ( 
.A(n_3504),
.B(n_2331),
.Y(n_3629)
);

OA21x2_ASAP7_75t_L g3630 ( 
.A1(n_3510),
.A2(n_1456),
.B(n_1455),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3532),
.Y(n_3631)
);

BUFx10_ASAP7_75t_L g3632 ( 
.A(n_3486),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_L g3633 ( 
.A1(n_3506),
.A2(n_1733),
.B1(n_1755),
.B2(n_1659),
.Y(n_3633)
);

AO21x2_ASAP7_75t_L g3634 ( 
.A1(n_3497),
.A2(n_2335),
.B(n_2333),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3531),
.Y(n_3635)
);

CKINVDCx20_ASAP7_75t_R g3636 ( 
.A(n_3535),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3492),
.A2(n_1755),
.B(n_1733),
.Y(n_3637)
);

AND2x6_ASAP7_75t_SL g3638 ( 
.A(n_3557),
.B(n_3),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3539),
.Y(n_3639)
);

BUFx6f_ASAP7_75t_L g3640 ( 
.A(n_3517),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3579),
.A2(n_2354),
.B(n_2335),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_L g3642 ( 
.A1(n_3519),
.A2(n_1755),
.B1(n_1756),
.B2(n_1733),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_3500),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3564),
.Y(n_3644)
);

OAI21x1_ASAP7_75t_L g3645 ( 
.A1(n_3552),
.A2(n_2362),
.B(n_2354),
.Y(n_3645)
);

AND2x4_ASAP7_75t_L g3646 ( 
.A(n_3581),
.B(n_2362),
.Y(n_3646)
);

OA21x2_ASAP7_75t_L g3647 ( 
.A1(n_3572),
.A2(n_1459),
.B(n_1458),
.Y(n_3647)
);

OAI21x1_ASAP7_75t_L g3648 ( 
.A1(n_3526),
.A2(n_2389),
.B(n_2364),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3542),
.Y(n_3649)
);

AND2x4_ASAP7_75t_L g3650 ( 
.A(n_3547),
.B(n_2364),
.Y(n_3650)
);

A2O1A1Ixp33_ASAP7_75t_L g3651 ( 
.A1(n_3501),
.A2(n_1463),
.B(n_1467),
.C(n_1466),
.Y(n_3651)
);

OA21x2_ASAP7_75t_L g3652 ( 
.A1(n_3550),
.A2(n_1470),
.B(n_1462),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3493),
.B(n_1472),
.Y(n_3653)
);

AND2x4_ASAP7_75t_L g3654 ( 
.A(n_3583),
.B(n_2389),
.Y(n_3654)
);

OAI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_3576),
.A2(n_1493),
.B(n_1474),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3514),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3514),
.Y(n_3657)
);

BUFx3_ASAP7_75t_L g3658 ( 
.A(n_3537),
.Y(n_3658)
);

INVx1_ASAP7_75t_SL g3659 ( 
.A(n_3540),
.Y(n_3659)
);

AND2x4_ASAP7_75t_L g3660 ( 
.A(n_3574),
.B(n_3585),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3573),
.Y(n_3661)
);

INVx6_ASAP7_75t_L g3662 ( 
.A(n_3517),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3509),
.B(n_3),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3565),
.Y(n_3664)
);

INVx6_ASAP7_75t_L g3665 ( 
.A(n_3585),
.Y(n_3665)
);

INVx3_ASAP7_75t_L g3666 ( 
.A(n_3498),
.Y(n_3666)
);

OAI21x1_ASAP7_75t_L g3667 ( 
.A1(n_3569),
.A2(n_3538),
.B(n_3561),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3555),
.B(n_3534),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3602),
.Y(n_3669)
);

INVx2_ASAP7_75t_SL g3670 ( 
.A(n_3626),
.Y(n_3670)
);

NAND2x1p5_ASAP7_75t_L g3671 ( 
.A(n_3666),
.B(n_3546),
.Y(n_3671)
);

BUFx12f_ASAP7_75t_L g3672 ( 
.A(n_3608),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3604),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3603),
.B(n_3558),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3625),
.B(n_3543),
.Y(n_3675)
);

HB1xp67_ASAP7_75t_L g3676 ( 
.A(n_3598),
.Y(n_3676)
);

BUFx2_ASAP7_75t_R g3677 ( 
.A(n_3612),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3610),
.Y(n_3678)
);

AO21x2_ASAP7_75t_L g3679 ( 
.A1(n_3657),
.A2(n_3578),
.B(n_3536),
.Y(n_3679)
);

AO21x1_ASAP7_75t_L g3680 ( 
.A1(n_3653),
.A2(n_3568),
.B(n_3530),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3637),
.A2(n_3482),
.B(n_3575),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3631),
.B(n_3521),
.Y(n_3682)
);

INVx3_ASAP7_75t_L g3683 ( 
.A(n_3640),
.Y(n_3683)
);

OAI21x1_ASAP7_75t_L g3684 ( 
.A1(n_3628),
.A2(n_3589),
.B(n_3563),
.Y(n_3684)
);

OAI21x1_ASAP7_75t_L g3685 ( 
.A1(n_3594),
.A2(n_3566),
.B(n_3484),
.Y(n_3685)
);

NAND2x1p5_ASAP7_75t_L g3686 ( 
.A(n_3640),
.B(n_3553),
.Y(n_3686)
);

OA21x2_ASAP7_75t_L g3687 ( 
.A1(n_3656),
.A2(n_3588),
.B(n_3570),
.Y(n_3687)
);

AOI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3601),
.A2(n_3567),
.B(n_3554),
.Y(n_3688)
);

HB1xp67_ASAP7_75t_L g3689 ( 
.A(n_3639),
.Y(n_3689)
);

OA21x2_ASAP7_75t_L g3690 ( 
.A1(n_3667),
.A2(n_3556),
.B(n_3549),
.Y(n_3690)
);

HB1xp67_ASAP7_75t_L g3691 ( 
.A(n_3644),
.Y(n_3691)
);

OAI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3648),
.A2(n_3524),
.B(n_3516),
.Y(n_3692)
);

AND2x4_ASAP7_75t_L g3693 ( 
.A(n_3597),
.B(n_3562),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3600),
.Y(n_3694)
);

OR2x2_ASAP7_75t_L g3695 ( 
.A(n_3664),
.B(n_3580),
.Y(n_3695)
);

OR2x2_ASAP7_75t_L g3696 ( 
.A(n_3661),
.B(n_1755),
.Y(n_3696)
);

AO31x2_ASAP7_75t_L g3697 ( 
.A1(n_3611),
.A2(n_3590),
.A3(n_3562),
.B(n_3511),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3605),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3643),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3622),
.B(n_1756),
.Y(n_3700)
);

AOI221xp5_ASAP7_75t_L g3701 ( 
.A1(n_3614),
.A2(n_1480),
.B1(n_1485),
.B2(n_1478),
.C(n_1477),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3622),
.B(n_1756),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3649),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3635),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3599),
.A2(n_3541),
.B(n_1767),
.Y(n_3705)
);

AOI21x1_ASAP7_75t_L g3706 ( 
.A1(n_3607),
.A2(n_3645),
.B(n_3641),
.Y(n_3706)
);

NOR2x1_ASAP7_75t_L g3707 ( 
.A(n_3660),
.B(n_1756),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3668),
.B(n_1767),
.Y(n_3708)
);

INVx3_ASAP7_75t_L g3709 ( 
.A(n_3626),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3646),
.Y(n_3710)
);

OAI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_3651),
.A2(n_3655),
.B(n_3615),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3616),
.A2(n_3634),
.B(n_3647),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3629),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3627),
.A2(n_1808),
.B(n_1767),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3668),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3650),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3593),
.Y(n_3717)
);

INVx2_ASAP7_75t_SL g3718 ( 
.A(n_3662),
.Y(n_3718)
);

BUFx8_ASAP7_75t_L g3719 ( 
.A(n_3658),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3609),
.B(n_1767),
.Y(n_3720)
);

BUFx2_ASAP7_75t_L g3721 ( 
.A(n_3623),
.Y(n_3721)
);

BUFx3_ASAP7_75t_L g3722 ( 
.A(n_3636),
.Y(n_3722)
);

BUFx3_ASAP7_75t_L g3723 ( 
.A(n_3606),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3662),
.Y(n_3724)
);

BUFx3_ASAP7_75t_L g3725 ( 
.A(n_3665),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3689),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3676),
.B(n_3659),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3691),
.B(n_3595),
.Y(n_3728)
);

OAI211xp5_ASAP7_75t_L g3729 ( 
.A1(n_3688),
.A2(n_3613),
.B(n_3617),
.C(n_3621),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3694),
.Y(n_3730)
);

BUFx3_ASAP7_75t_L g3731 ( 
.A(n_3719),
.Y(n_3731)
);

OAI21x1_ASAP7_75t_L g3732 ( 
.A1(n_3706),
.A2(n_3630),
.B(n_3642),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3669),
.Y(n_3733)
);

OA21x2_ASAP7_75t_L g3734 ( 
.A1(n_3705),
.A2(n_3596),
.B(n_3624),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3673),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_3721),
.B(n_3674),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3698),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3678),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3715),
.Y(n_3739)
);

HB1xp67_ASAP7_75t_L g3740 ( 
.A(n_3675),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3721),
.B(n_3663),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3682),
.B(n_3663),
.Y(n_3742)
);

AOI21x1_ASAP7_75t_L g3743 ( 
.A1(n_3706),
.A2(n_3654),
.B(n_3652),
.Y(n_3743)
);

AO21x1_ASAP7_75t_SL g3744 ( 
.A1(n_3717),
.A2(n_3620),
.B(n_3618),
.Y(n_3744)
);

INVx3_ASAP7_75t_L g3745 ( 
.A(n_3725),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3699),
.Y(n_3746)
);

OAI21x1_ASAP7_75t_L g3747 ( 
.A1(n_3712),
.A2(n_3633),
.B(n_3619),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3703),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3696),
.Y(n_3749)
);

HB1xp67_ASAP7_75t_L g3750 ( 
.A(n_3700),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3724),
.B(n_3632),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3693),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3683),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3685),
.A2(n_3593),
.B(n_3665),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3704),
.Y(n_3755)
);

BUFx2_ASAP7_75t_L g3756 ( 
.A(n_3672),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3708),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3695),
.Y(n_3758)
);

HB1xp67_ASAP7_75t_L g3759 ( 
.A(n_3702),
.Y(n_3759)
);

OA21x2_ASAP7_75t_L g3760 ( 
.A1(n_3684),
.A2(n_1489),
.B(n_1488),
.Y(n_3760)
);

OR2x6_ASAP7_75t_L g3761 ( 
.A(n_3670),
.B(n_3638),
.Y(n_3761)
);

CKINVDCx20_ASAP7_75t_R g3762 ( 
.A(n_3722),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3710),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3720),
.B(n_1808),
.Y(n_3764)
);

OA21x2_ASAP7_75t_L g3765 ( 
.A1(n_3713),
.A2(n_1496),
.B(n_1490),
.Y(n_3765)
);

HB1xp67_ASAP7_75t_L g3766 ( 
.A(n_3687),
.Y(n_3766)
);

AO21x2_ASAP7_75t_L g3767 ( 
.A1(n_3680),
.A2(n_1885),
.B(n_1808),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3723),
.B(n_1808),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3677),
.B(n_1885),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3697),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3697),
.Y(n_3771)
);

HB1xp67_ASAP7_75t_L g3772 ( 
.A(n_3687),
.Y(n_3772)
);

OA21x2_ASAP7_75t_L g3773 ( 
.A1(n_3714),
.A2(n_1498),
.B(n_1497),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3716),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3679),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_L g3776 ( 
.A(n_3709),
.B(n_1885),
.Y(n_3776)
);

OA21x2_ASAP7_75t_L g3777 ( 
.A1(n_3692),
.A2(n_3681),
.B(n_3711),
.Y(n_3777)
);

BUFx2_ASAP7_75t_L g3778 ( 
.A(n_3718),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3707),
.A2(n_3690),
.B(n_3686),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3690),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3671),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3701),
.B(n_1885),
.Y(n_3782)
);

BUFx2_ASAP7_75t_L g3783 ( 
.A(n_3676),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3694),
.Y(n_3784)
);

AND2x4_ASAP7_75t_L g3785 ( 
.A(n_3783),
.B(n_4),
.Y(n_3785)
);

OAI22xp5_ASAP7_75t_SL g3786 ( 
.A1(n_3761),
.A2(n_1501),
.B1(n_1503),
.B2(n_1499),
.Y(n_3786)
);

INVx1_ASAP7_75t_SL g3787 ( 
.A(n_3762),
.Y(n_3787)
);

OAI22xp5_ASAP7_75t_L g3788 ( 
.A1(n_3736),
.A2(n_1508),
.B1(n_1510),
.B2(n_1506),
.Y(n_3788)
);

OAI22xp33_ASAP7_75t_L g3789 ( 
.A1(n_3777),
.A2(n_1517),
.B1(n_1520),
.B2(n_1511),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3740),
.B(n_1516),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3734),
.A2(n_1888),
.B1(n_1526),
.B2(n_1532),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3755),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3755),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3777),
.A2(n_1535),
.B(n_1525),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3779),
.A2(n_4),
.B(n_5),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3752),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3726),
.B(n_3750),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3759),
.B(n_1538),
.Y(n_3798)
);

OAI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_3729),
.A2(n_3768),
.B(n_3760),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3733),
.Y(n_3800)
);

AOI22xp33_ASAP7_75t_L g3801 ( 
.A1(n_3734),
.A2(n_1546),
.B1(n_1547),
.B2(n_1542),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3760),
.A2(n_1550),
.B1(n_1551),
.B2(n_1549),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3727),
.B(n_6),
.Y(n_3803)
);

AOI22xp33_ASAP7_75t_L g3804 ( 
.A1(n_3765),
.A2(n_1884),
.B1(n_1556),
.B2(n_1562),
.Y(n_3804)
);

AOI211xp5_ASAP7_75t_L g3805 ( 
.A1(n_3769),
.A2(n_1563),
.B(n_1564),
.C(n_1553),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3765),
.A2(n_1569),
.B1(n_1570),
.B2(n_1568),
.Y(n_3806)
);

AOI22xp33_ASAP7_75t_SL g3807 ( 
.A1(n_3767),
.A2(n_1591),
.B1(n_1609),
.B2(n_1575),
.Y(n_3807)
);

BUFx6f_ASAP7_75t_L g3808 ( 
.A(n_3731),
.Y(n_3808)
);

BUFx2_ASAP7_75t_L g3809 ( 
.A(n_3745),
.Y(n_3809)
);

AOI22xp5_ASAP7_75t_L g3810 ( 
.A1(n_3761),
.A2(n_1572),
.B1(n_1574),
.B2(n_1571),
.Y(n_3810)
);

OAI22xp5_ASAP7_75t_L g3811 ( 
.A1(n_3745),
.A2(n_1579),
.B1(n_1581),
.B2(n_1577),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3778),
.B(n_6),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3735),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3738),
.Y(n_3814)
);

NAND4xp25_ASAP7_75t_L g3815 ( 
.A(n_3728),
.B(n_3780),
.C(n_3756),
.D(n_3742),
.Y(n_3815)
);

BUFx6f_ASAP7_75t_L g3816 ( 
.A(n_3751),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_L g3817 ( 
.A1(n_3744),
.A2(n_1584),
.B1(n_1585),
.B2(n_1583),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3781),
.A2(n_1592),
.B1(n_1593),
.B2(n_1587),
.Y(n_3818)
);

INVxp67_ASAP7_75t_L g3819 ( 
.A(n_3809),
.Y(n_3819)
);

BUFx3_ASAP7_75t_L g3820 ( 
.A(n_3808),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3792),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3800),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3813),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3793),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3814),
.Y(n_3825)
);

INVx1_ASAP7_75t_SL g3826 ( 
.A(n_3787),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3797),
.B(n_3739),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3796),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3790),
.B(n_3757),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3785),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3785),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3815),
.B(n_3757),
.Y(n_3832)
);

INVxp67_ASAP7_75t_SL g3833 ( 
.A(n_3789),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3816),
.B(n_3741),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3798),
.B(n_3812),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3816),
.B(n_3753),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3795),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3803),
.Y(n_3838)
);

OR2x2_ASAP7_75t_L g3839 ( 
.A(n_3799),
.B(n_3758),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3794),
.B(n_3746),
.Y(n_3840)
);

OAI221xp5_ASAP7_75t_SL g3841 ( 
.A1(n_3804),
.A2(n_3782),
.B1(n_3776),
.B2(n_3764),
.C(n_3766),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3791),
.Y(n_3842)
);

AND2x4_ASAP7_75t_L g3843 ( 
.A(n_3808),
.B(n_3753),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3810),
.B(n_3763),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3788),
.B(n_3749),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3801),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3802),
.B(n_3748),
.Y(n_3847)
);

OR2x2_ASAP7_75t_L g3848 ( 
.A(n_3818),
.B(n_3737),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3786),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3806),
.B(n_3772),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3817),
.B(n_3774),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3822),
.Y(n_3852)
);

INVx2_ASAP7_75t_SL g3853 ( 
.A(n_3820),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3836),
.B(n_3754),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3834),
.B(n_3775),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3837),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_L g3857 ( 
.A1(n_3832),
.A2(n_3807),
.B1(n_3805),
.B2(n_3811),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3824),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3829),
.B(n_3732),
.Y(n_3859)
);

OR2x6_ASAP7_75t_SL g3860 ( 
.A(n_3835),
.B(n_3770),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3823),
.B(n_3743),
.Y(n_3861)
);

BUFx2_ASAP7_75t_L g3862 ( 
.A(n_3843),
.Y(n_3862)
);

NOR2xp33_ASAP7_75t_L g3863 ( 
.A(n_3849),
.B(n_7),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3825),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3828),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3827),
.B(n_3773),
.Y(n_3866)
);

BUFx2_ASAP7_75t_L g3867 ( 
.A(n_3843),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3819),
.B(n_3730),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3838),
.B(n_3784),
.Y(n_3869)
);

OA21x2_ASAP7_75t_L g3870 ( 
.A1(n_3821),
.A2(n_3771),
.B(n_3747),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3838),
.B(n_3773),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3830),
.B(n_8),
.Y(n_3872)
);

HB1xp67_ASAP7_75t_L g3873 ( 
.A(n_3821),
.Y(n_3873)
);

OR2x2_ASAP7_75t_L g3874 ( 
.A(n_3839),
.B(n_9),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3840),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3831),
.B(n_10),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3826),
.B(n_10),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3845),
.B(n_12),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3833),
.B(n_1594),
.Y(n_3879)
);

INVx2_ASAP7_75t_SL g3880 ( 
.A(n_3848),
.Y(n_3880)
);

INVxp67_ASAP7_75t_SL g3881 ( 
.A(n_3850),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3844),
.B(n_15),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3841),
.A2(n_1600),
.B(n_1595),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3851),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3847),
.B(n_16),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3846),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3852),
.Y(n_3887)
);

AND2x4_ASAP7_75t_L g3888 ( 
.A(n_3862),
.B(n_3842),
.Y(n_3888)
);

BUFx2_ASAP7_75t_L g3889 ( 
.A(n_3867),
.Y(n_3889)
);

OR2x2_ASAP7_75t_L g3890 ( 
.A(n_3875),
.B(n_3842),
.Y(n_3890)
);

AOI22xp33_ASAP7_75t_L g3891 ( 
.A1(n_3881),
.A2(n_1604),
.B1(n_1611),
.B2(n_1603),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3875),
.B(n_1612),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3880),
.Y(n_3893)
);

OAI221xp5_ASAP7_75t_L g3894 ( 
.A1(n_3874),
.A2(n_1621),
.B1(n_1622),
.B2(n_1620),
.C(n_1613),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3871),
.B(n_1623),
.Y(n_3895)
);

NAND3xp33_ASAP7_75t_L g3896 ( 
.A(n_3866),
.B(n_3856),
.C(n_3857),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3853),
.B(n_16),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3852),
.Y(n_3898)
);

NOR2x1_ASAP7_75t_L g3899 ( 
.A(n_3877),
.B(n_17),
.Y(n_3899)
);

OAI221xp5_ASAP7_75t_L g3900 ( 
.A1(n_3879),
.A2(n_1628),
.B1(n_1629),
.B2(n_1625),
.C(n_1624),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3855),
.Y(n_3901)
);

AOI21xp33_ASAP7_75t_L g3902 ( 
.A1(n_3859),
.A2(n_1632),
.B(n_1630),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3864),
.Y(n_3903)
);

AOI22xp33_ASAP7_75t_L g3904 ( 
.A1(n_3886),
.A2(n_1637),
.B1(n_1639),
.B2(n_1633),
.Y(n_3904)
);

NOR3xp33_ASAP7_75t_L g3905 ( 
.A(n_3863),
.B(n_1648),
.C(n_1645),
.Y(n_3905)
);

HB1xp67_ASAP7_75t_L g3906 ( 
.A(n_3864),
.Y(n_3906)
);

AOI221xp5_ASAP7_75t_L g3907 ( 
.A1(n_3883),
.A2(n_1653),
.B1(n_1660),
.B2(n_1652),
.C(n_1650),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3868),
.B(n_19),
.Y(n_3908)
);

INVxp67_ASAP7_75t_L g3909 ( 
.A(n_3878),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3885),
.B(n_1666),
.Y(n_3910)
);

NOR2xp33_ASAP7_75t_L g3911 ( 
.A(n_3882),
.B(n_1877),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3873),
.Y(n_3912)
);

NOR2xp33_ASAP7_75t_L g3913 ( 
.A(n_3872),
.B(n_1879),
.Y(n_3913)
);

OAI221xp5_ASAP7_75t_L g3914 ( 
.A1(n_3886),
.A2(n_1672),
.B1(n_1675),
.B2(n_1668),
.C(n_1667),
.Y(n_3914)
);

NAND4xp25_ASAP7_75t_L g3915 ( 
.A(n_3861),
.B(n_23),
.C(n_20),
.D(n_21),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3854),
.B(n_20),
.Y(n_3916)
);

INVx2_ASAP7_75t_SL g3917 ( 
.A(n_3876),
.Y(n_3917)
);

HB1xp67_ASAP7_75t_L g3918 ( 
.A(n_3865),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3869),
.B(n_21),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3906),
.Y(n_3920)
);

OAI31xp33_ASAP7_75t_L g3921 ( 
.A1(n_3896),
.A2(n_3860),
.A3(n_3884),
.B(n_3858),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3887),
.Y(n_3922)
);

NAND2xp33_ASAP7_75t_L g3923 ( 
.A(n_3899),
.B(n_1678),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3889),
.B(n_3870),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3909),
.B(n_3870),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3898),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3888),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3903),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3897),
.B(n_23),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3916),
.B(n_24),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3888),
.B(n_1680),
.Y(n_3931)
);

BUFx2_ASAP7_75t_L g3932 ( 
.A(n_3893),
.Y(n_3932)
);

AOI21xp5_ASAP7_75t_SL g3933 ( 
.A1(n_3908),
.A2(n_1684),
.B(n_1681),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3918),
.Y(n_3934)
);

HB1xp67_ASAP7_75t_L g3935 ( 
.A(n_3912),
.Y(n_3935)
);

NAND4xp25_ASAP7_75t_L g3936 ( 
.A(n_3915),
.B(n_3891),
.C(n_3902),
.D(n_3907),
.Y(n_3936)
);

AND2x2_ASAP7_75t_L g3937 ( 
.A(n_3901),
.B(n_24),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3917),
.B(n_25),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3919),
.Y(n_3939)
);

NAND3xp33_ASAP7_75t_L g3940 ( 
.A(n_3905),
.B(n_1687),
.C(n_1686),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3895),
.B(n_3892),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3911),
.B(n_1691),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3890),
.Y(n_3943)
);

INVxp33_ASAP7_75t_L g3944 ( 
.A(n_3913),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3894),
.Y(n_3945)
);

AND2x4_ASAP7_75t_L g3946 ( 
.A(n_3910),
.B(n_26),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3904),
.B(n_3914),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3900),
.B(n_26),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3909),
.B(n_1693),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3906),
.Y(n_3950)
);

AND2x2_ASAP7_75t_L g3951 ( 
.A(n_3889),
.B(n_27),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3909),
.B(n_28),
.Y(n_3952)
);

OR2x2_ASAP7_75t_L g3953 ( 
.A(n_3909),
.B(n_29),
.Y(n_3953)
);

NAND4xp75_ASAP7_75t_L g3954 ( 
.A(n_3899),
.B(n_32),
.C(n_30),
.D(n_31),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3909),
.B(n_1694),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_SL g3956 ( 
.A(n_3888),
.B(n_1696),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3889),
.B(n_30),
.Y(n_3957)
);

OAI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3915),
.A2(n_1712),
.B(n_1697),
.Y(n_3958)
);

HB1xp67_ASAP7_75t_L g3959 ( 
.A(n_3889),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3889),
.B(n_31),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3894),
.B(n_1698),
.Y(n_3961)
);

OR2x2_ASAP7_75t_L g3962 ( 
.A(n_3909),
.B(n_33),
.Y(n_3962)
);

OR2x6_ASAP7_75t_L g3963 ( 
.A(n_3899),
.B(n_34),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3889),
.B(n_35),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3932),
.B(n_36),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3927),
.B(n_36),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3939),
.B(n_1699),
.Y(n_3967)
);

OR2x2_ASAP7_75t_L g3968 ( 
.A(n_3959),
.B(n_37),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3951),
.B(n_3957),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_3960),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3964),
.B(n_3941),
.Y(n_3971)
);

AND2x4_ASAP7_75t_L g3972 ( 
.A(n_3934),
.B(n_38),
.Y(n_3972)
);

BUFx2_ASAP7_75t_L g3973 ( 
.A(n_3935),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3938),
.B(n_38),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3933),
.B(n_1703),
.Y(n_3975)
);

OR2x2_ASAP7_75t_L g3976 ( 
.A(n_3943),
.B(n_3952),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3937),
.B(n_1704),
.Y(n_3977)
);

NAND2xp33_ASAP7_75t_SL g3978 ( 
.A(n_3956),
.B(n_1705),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3953),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3962),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3947),
.B(n_39),
.Y(n_3981)
);

OR2x2_ASAP7_75t_L g3982 ( 
.A(n_3950),
.B(n_40),
.Y(n_3982)
);

AND2x2_ASAP7_75t_L g3983 ( 
.A(n_3929),
.B(n_42),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3930),
.B(n_42),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3920),
.B(n_43),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3946),
.B(n_3931),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3920),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3949),
.B(n_3955),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3946),
.B(n_3945),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3922),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3925),
.B(n_1707),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3926),
.Y(n_3992)
);

OR2x2_ASAP7_75t_L g3993 ( 
.A(n_3928),
.B(n_44),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3944),
.B(n_1711),
.Y(n_3994)
);

OAI21xp33_ASAP7_75t_L g3995 ( 
.A1(n_3936),
.A2(n_1717),
.B(n_1715),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3963),
.B(n_1718),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3963),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3948),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3954),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3924),
.B(n_44),
.Y(n_4000)
);

OAI22xp5_ASAP7_75t_L g4001 ( 
.A1(n_3921),
.A2(n_1721),
.B1(n_1723),
.B2(n_1720),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3942),
.B(n_45),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3958),
.B(n_3923),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3940),
.Y(n_4004)
);

OAI32xp33_ASAP7_75t_L g4005 ( 
.A1(n_3961),
.A2(n_1735),
.A3(n_1736),
.B1(n_1734),
.B2(n_1732),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3959),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3932),
.B(n_45),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3963),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3959),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3959),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3959),
.Y(n_4011)
);

INVxp67_ASAP7_75t_L g4012 ( 
.A(n_3963),
.Y(n_4012)
);

NOR2xp67_ASAP7_75t_L g4013 ( 
.A(n_3959),
.B(n_46),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3939),
.B(n_1737),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3939),
.B(n_1738),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3959),
.B(n_47),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3932),
.B(n_48),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3959),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3939),
.B(n_1741),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3932),
.B(n_49),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3939),
.B(n_1742),
.Y(n_4021)
);

BUFx2_ASAP7_75t_L g4022 ( 
.A(n_3927),
.Y(n_4022)
);

INVxp67_ASAP7_75t_SL g4023 ( 
.A(n_3959),
.Y(n_4023)
);

OR2x2_ASAP7_75t_L g4024 ( 
.A(n_3959),
.B(n_49),
.Y(n_4024)
);

AND2x2_ASAP7_75t_SL g4025 ( 
.A(n_3932),
.B(n_50),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_3939),
.B(n_1743),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3932),
.B(n_51),
.Y(n_4027)
);

NAND2x1_ASAP7_75t_L g4028 ( 
.A(n_3927),
.B(n_51),
.Y(n_4028)
);

OR2x2_ASAP7_75t_L g4029 ( 
.A(n_3959),
.B(n_52),
.Y(n_4029)
);

HB1xp67_ASAP7_75t_L g4030 ( 
.A(n_3970),
.Y(n_4030)
);

NOR3xp33_ASAP7_75t_L g4031 ( 
.A(n_4001),
.B(n_1746),
.C(n_1744),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_4023),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3973),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3965),
.B(n_1749),
.Y(n_4034)
);

INVx1_ASAP7_75t_SL g4035 ( 
.A(n_3969),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_4025),
.Y(n_4036)
);

AOI32xp33_ASAP7_75t_L g4037 ( 
.A1(n_4000),
.A2(n_1759),
.A3(n_1760),
.B1(n_1753),
.B2(n_1751),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_SL g4038 ( 
.A(n_3971),
.B(n_1761),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3968),
.Y(n_4039)
);

AOI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_4013),
.A2(n_1768),
.B(n_1763),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_4007),
.B(n_4017),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_4016),
.Y(n_4042)
);

INVxp67_ASAP7_75t_L g4043 ( 
.A(n_3975),
.Y(n_4043)
);

OR2x2_ASAP7_75t_L g4044 ( 
.A(n_3976),
.B(n_4006),
.Y(n_4044)
);

INVx2_ASAP7_75t_SL g4045 ( 
.A(n_4020),
.Y(n_4045)
);

AOI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_3998),
.A2(n_1774),
.B1(n_1775),
.B2(n_1772),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3985),
.B(n_1778),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_4024),
.Y(n_4048)
);

OAI31xp33_ASAP7_75t_L g4049 ( 
.A1(n_3997),
.A2(n_54),
.A3(n_52),
.B(n_53),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_4029),
.Y(n_4050)
);

BUFx2_ASAP7_75t_L g4051 ( 
.A(n_4022),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_4027),
.B(n_1779),
.Y(n_4052)
);

INVx2_ASAP7_75t_L g4053 ( 
.A(n_4028),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3972),
.B(n_1782),
.Y(n_4054)
);

INVx2_ASAP7_75t_SL g4055 ( 
.A(n_3972),
.Y(n_4055)
);

OAI21xp5_ASAP7_75t_SL g4056 ( 
.A1(n_4009),
.A2(n_55),
.B(n_56),
.Y(n_4056)
);

AND2x4_ASAP7_75t_L g4057 ( 
.A(n_3966),
.B(n_55),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_4010),
.Y(n_4058)
);

OAI321xp33_ASAP7_75t_L g4059 ( 
.A1(n_3987),
.A2(n_2404),
.A3(n_2395),
.B1(n_2406),
.B2(n_2398),
.C(n_2391),
.Y(n_4059)
);

AND2x4_ASAP7_75t_L g4060 ( 
.A(n_4012),
.B(n_57),
.Y(n_4060)
);

AOI21xp33_ASAP7_75t_L g4061 ( 
.A1(n_3989),
.A2(n_1788),
.B(n_1785),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_4011),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_4018),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3984),
.B(n_1790),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3983),
.B(n_1792),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3974),
.B(n_1794),
.Y(n_4066)
);

XOR2x2_ASAP7_75t_L g4067 ( 
.A(n_3981),
.B(n_57),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3994),
.Y(n_4068)
);

INVx2_ASAP7_75t_L g4069 ( 
.A(n_3993),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3988),
.B(n_1795),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3967),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_4014),
.Y(n_4072)
);

NAND3xp33_ASAP7_75t_L g4073 ( 
.A(n_4008),
.B(n_1798),
.C(n_1796),
.Y(n_4073)
);

INVxp67_ASAP7_75t_SL g4074 ( 
.A(n_3977),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3982),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3979),
.B(n_1799),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_4015),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4019),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_4021),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_4026),
.Y(n_4080)
);

AOI31xp33_ASAP7_75t_L g4081 ( 
.A1(n_3980),
.A2(n_1802),
.A3(n_1805),
.B(n_1801),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3990),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3992),
.Y(n_4083)
);

AOI32xp33_ASAP7_75t_L g4084 ( 
.A1(n_3999),
.A2(n_1812),
.A3(n_1815),
.B1(n_1810),
.B2(n_1806),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4004),
.B(n_1817),
.Y(n_4085)
);

NAND3xp33_ASAP7_75t_L g4086 ( 
.A(n_3991),
.B(n_1823),
.C(n_1820),
.Y(n_4086)
);

INVx2_ASAP7_75t_SL g4087 ( 
.A(n_4002),
.Y(n_4087)
);

OAI221xp5_ASAP7_75t_L g4088 ( 
.A1(n_3986),
.A2(n_1827),
.B1(n_1829),
.B2(n_1826),
.C(n_1825),
.Y(n_4088)
);

AOI22xp5_ASAP7_75t_L g4089 ( 
.A1(n_4003),
.A2(n_1832),
.B1(n_1833),
.B2(n_1830),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3996),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3995),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4005),
.Y(n_4092)
);

NAND3xp33_ASAP7_75t_L g4093 ( 
.A(n_3978),
.B(n_1836),
.C(n_1834),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4005),
.Y(n_4094)
);

NOR3xp33_ASAP7_75t_L g4095 ( 
.A(n_4001),
.B(n_1843),
.C(n_1840),
.Y(n_4095)
);

AOI21xp33_ASAP7_75t_SL g4096 ( 
.A1(n_4001),
.A2(n_68),
.B(n_58),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3970),
.B(n_1845),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_3969),
.B(n_1846),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4023),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4023),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_4023),
.Y(n_4101)
);

OAI221xp5_ASAP7_75t_L g4102 ( 
.A1(n_4001),
.A2(n_1849),
.B1(n_1850),
.B2(n_1848),
.C(n_1847),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4023),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4023),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4023),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_4023),
.Y(n_4106)
);

OAI32xp33_ASAP7_75t_L g4107 ( 
.A1(n_4001),
.A2(n_1864),
.A3(n_1865),
.B1(n_1861),
.B2(n_1860),
.Y(n_4107)
);

NOR2xp33_ASAP7_75t_SL g4108 ( 
.A(n_3970),
.B(n_1869),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4023),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_4025),
.Y(n_4110)
);

INVx1_ASAP7_75t_SL g4111 ( 
.A(n_3969),
.Y(n_4111)
);

AND2x2_ASAP7_75t_L g4112 ( 
.A(n_3969),
.B(n_1867),
.Y(n_4112)
);

NOR2xp33_ASAP7_75t_L g4113 ( 
.A(n_3971),
.B(n_1868),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4023),
.Y(n_4114)
);

OAI22xp33_ASAP7_75t_L g4115 ( 
.A1(n_4001),
.A2(n_1872),
.B1(n_1873),
.B2(n_1871),
.Y(n_4115)
);

OR2x2_ASAP7_75t_L g4116 ( 
.A(n_3971),
.B(n_58),
.Y(n_4116)
);

INVxp67_ASAP7_75t_L g4117 ( 
.A(n_4051),
.Y(n_4117)
);

HB1xp67_ASAP7_75t_L g4118 ( 
.A(n_4030),
.Y(n_4118)
);

OR2x2_ASAP7_75t_L g4119 ( 
.A(n_4035),
.B(n_59),
.Y(n_4119)
);

NOR2xp33_ASAP7_75t_L g4120 ( 
.A(n_4108),
.B(n_1874),
.Y(n_4120)
);

INVx2_ASAP7_75t_SL g4121 ( 
.A(n_4055),
.Y(n_4121)
);

INVxp67_ASAP7_75t_L g4122 ( 
.A(n_4070),
.Y(n_4122)
);

AOI322xp5_ASAP7_75t_L g4123 ( 
.A1(n_4036),
.A2(n_1886),
.A3(n_1887),
.B1(n_1883),
.B2(n_62),
.C1(n_66),
.C2(n_64),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4111),
.B(n_4098),
.Y(n_4124)
);

OAI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_4045),
.A2(n_63),
.B1(n_59),
.B2(n_60),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4116),
.Y(n_4126)
);

NOR2xp33_ASAP7_75t_L g4127 ( 
.A(n_4081),
.B(n_60),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_4087),
.B(n_64),
.Y(n_4128)
);

AOI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_4110),
.A2(n_2395),
.B1(n_2398),
.B2(n_2391),
.Y(n_4129)
);

OAI211xp5_ASAP7_75t_L g4130 ( 
.A1(n_4032),
.A2(n_69),
.B(n_66),
.C(n_67),
.Y(n_4130)
);

INVxp67_ASAP7_75t_L g4131 ( 
.A(n_4041),
.Y(n_4131)
);

OR2x2_ASAP7_75t_L g4132 ( 
.A(n_4044),
.B(n_69),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4076),
.Y(n_4133)
);

OAI22xp33_ASAP7_75t_L g4134 ( 
.A1(n_4053),
.A2(n_4075),
.B1(n_4039),
.B2(n_4048),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_4099),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_4112),
.B(n_70),
.Y(n_4136)
);

OAI31xp33_ASAP7_75t_L g4137 ( 
.A1(n_4092),
.A2(n_4094),
.A3(n_4056),
.B(n_4042),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_4047),
.B(n_70),
.Y(n_4138)
);

OAI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_4100),
.A2(n_71),
.B(n_74),
.Y(n_4139)
);

INVx2_ASAP7_75t_SL g4140 ( 
.A(n_4033),
.Y(n_4140)
);

INVxp67_ASAP7_75t_L g4141 ( 
.A(n_4057),
.Y(n_4141)
);

OAI32xp33_ASAP7_75t_L g4142 ( 
.A1(n_4101),
.A2(n_75),
.A3(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4103),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4104),
.Y(n_4144)
);

NAND4xp25_ASAP7_75t_L g4145 ( 
.A(n_4105),
.B(n_78),
.C(n_76),
.D(n_77),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_4057),
.Y(n_4146)
);

OAI21xp33_ASAP7_75t_SL g4147 ( 
.A1(n_4106),
.A2(n_77),
.B(n_79),
.Y(n_4147)
);

OAI32xp33_ASAP7_75t_L g4148 ( 
.A1(n_4109),
.A2(n_82),
.A3(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_SL g4149 ( 
.A(n_4037),
.B(n_4114),
.Y(n_4149)
);

AOI21xp33_ASAP7_75t_SL g4150 ( 
.A1(n_4050),
.A2(n_80),
.B(n_83),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4085),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4074),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_4060),
.B(n_4113),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4060),
.B(n_84),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4069),
.B(n_85),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4097),
.Y(n_4156)
);

NOR3xp33_ASAP7_75t_L g4157 ( 
.A(n_4043),
.B(n_85),
.C(n_86),
.Y(n_4157)
);

AOI221xp5_ASAP7_75t_L g4158 ( 
.A1(n_4090),
.A2(n_4068),
.B1(n_4071),
.B2(n_4077),
.C(n_4072),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4064),
.Y(n_4159)
);

AND2x4_ASAP7_75t_L g4160 ( 
.A(n_4058),
.B(n_86),
.Y(n_4160)
);

AOI21xp33_ASAP7_75t_L g4161 ( 
.A1(n_4082),
.A2(n_87),
.B(n_89),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4065),
.Y(n_4162)
);

OAI21xp33_ASAP7_75t_SL g4163 ( 
.A1(n_4083),
.A2(n_87),
.B(n_90),
.Y(n_4163)
);

AOI32xp33_ASAP7_75t_L g4164 ( 
.A1(n_4062),
.A2(n_109),
.A3(n_118),
.B1(n_100),
.B2(n_91),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4066),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_4063),
.B(n_92),
.Y(n_4166)
);

AOI22xp33_ASAP7_75t_L g4167 ( 
.A1(n_4078),
.A2(n_2406),
.B1(n_2412),
.B2(n_2404),
.Y(n_4167)
);

AOI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_4079),
.A2(n_2421),
.B1(n_2422),
.B2(n_2412),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4067),
.Y(n_4169)
);

O2A1O1Ixp33_ASAP7_75t_L g4170 ( 
.A1(n_4096),
.A2(n_96),
.B(n_93),
.C(n_94),
.Y(n_4170)
);

NOR2xp33_ASAP7_75t_L g4171 ( 
.A(n_4034),
.B(n_94),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4049),
.B(n_96),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4054),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4080),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4084),
.B(n_97),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_4038),
.B(n_98),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4046),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_4052),
.B(n_99),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4091),
.Y(n_4179)
);

OAI321xp33_ASAP7_75t_L g4180 ( 
.A1(n_4073),
.A2(n_103),
.A3(n_105),
.B1(n_106),
.B2(n_102),
.C(n_104),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_4086),
.A2(n_104),
.B1(n_100),
.B2(n_102),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4089),
.B(n_105),
.Y(n_4182)
);

OR2x2_ASAP7_75t_L g4183 ( 
.A(n_4088),
.B(n_4061),
.Y(n_4183)
);

OAI221xp5_ASAP7_75t_SL g4184 ( 
.A1(n_4031),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.C(n_110),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4093),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_R g4186 ( 
.A(n_4107),
.B(n_107),
.Y(n_4186)
);

INVx1_ASAP7_75t_SL g4187 ( 
.A(n_4040),
.Y(n_4187)
);

INVx1_ASAP7_75t_SL g4188 ( 
.A(n_4095),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4115),
.B(n_111),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4102),
.B(n_112),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4059),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_4051),
.Y(n_4192)
);

OAI22x1_ASAP7_75t_L g4193 ( 
.A1(n_4051),
.A2(n_116),
.B1(n_117),
.B2(n_115),
.Y(n_4193)
);

AOI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_4036),
.A2(n_2422),
.B1(n_2424),
.B2(n_2421),
.Y(n_4194)
);

INVx2_ASAP7_75t_SL g4195 ( 
.A(n_4051),
.Y(n_4195)
);

AOI22xp33_ASAP7_75t_L g4196 ( 
.A1(n_4036),
.A2(n_2425),
.B1(n_2424),
.B2(n_118),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4051),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4051),
.Y(n_4198)
);

OAI221xp5_ASAP7_75t_SL g4199 ( 
.A1(n_4035),
.A2(n_119),
.B1(n_114),
.B2(n_116),
.C(n_120),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4051),
.B(n_114),
.Y(n_4200)
);

OAI221xp5_ASAP7_75t_L g4201 ( 
.A1(n_4036),
.A2(n_122),
.B1(n_119),
.B2(n_120),
.C(n_123),
.Y(n_4201)
);

O2A1O1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_4056),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_4202)
);

OAI32xp33_ASAP7_75t_L g4203 ( 
.A1(n_4032),
.A2(n_128),
.A3(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4051),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4087),
.B(n_127),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_4036),
.A2(n_2425),
.B1(n_130),
.B2(n_128),
.Y(n_4206)
);

NAND2x1_ASAP7_75t_L g4207 ( 
.A(n_4051),
.B(n_129),
.Y(n_4207)
);

AOI21xp33_ASAP7_75t_SL g4208 ( 
.A1(n_4055),
.A2(n_130),
.B(n_131),
.Y(n_4208)
);

NAND3xp33_ASAP7_75t_L g4209 ( 
.A(n_4051),
.B(n_131),
.C(n_132),
.Y(n_4209)
);

AND2x4_ASAP7_75t_L g4210 ( 
.A(n_4055),
.B(n_134),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4051),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4051),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4051),
.Y(n_4213)
);

OR2x2_ASAP7_75t_L g4214 ( 
.A(n_4035),
.B(n_134),
.Y(n_4214)
);

NOR3xp33_ASAP7_75t_L g4215 ( 
.A(n_4092),
.B(n_135),
.C(n_138),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_4051),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4087),
.B(n_135),
.Y(n_4217)
);

NAND2xp33_ASAP7_75t_R g4218 ( 
.A(n_4051),
.B(n_139),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_4051),
.B(n_139),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4051),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4051),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4051),
.Y(n_4222)
);

OAI22xp5_ASAP7_75t_L g4223 ( 
.A1(n_4035),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_4051),
.B(n_143),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4051),
.B(n_143),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4051),
.B(n_144),
.Y(n_4226)
);

AOI222xp33_ASAP7_75t_L g4227 ( 
.A1(n_4092),
.A2(n_148),
.B1(n_150),
.B2(n_144),
.C1(n_146),
.C2(n_149),
.Y(n_4227)
);

NOR3xp33_ASAP7_75t_L g4228 ( 
.A(n_4092),
.B(n_146),
.C(n_148),
.Y(n_4228)
);

INVx2_ASAP7_75t_SL g4229 ( 
.A(n_4051),
.Y(n_4229)
);

AOI222xp33_ASAP7_75t_L g4230 ( 
.A1(n_4092),
.A2(n_151),
.B1(n_153),
.B2(n_149),
.C1(n_150),
.C2(n_152),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4087),
.B(n_151),
.Y(n_4231)
);

INVx3_ASAP7_75t_L g4232 ( 
.A(n_4051),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4051),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4087),
.B(n_152),
.Y(n_4234)
);

O2A1O1Ixp33_ASAP7_75t_L g4235 ( 
.A1(n_4056),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_4235)
);

AOI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4036),
.A2(n_157),
.B1(n_154),
.B2(n_156),
.Y(n_4236)
);

NAND3xp33_ASAP7_75t_L g4237 ( 
.A(n_4051),
.B(n_157),
.C(n_158),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4087),
.B(n_159),
.Y(n_4238)
);

AOI322xp5_ASAP7_75t_L g4239 ( 
.A1(n_4036),
.A2(n_164),
.A3(n_163),
.B1(n_161),
.B2(n_159),
.C1(n_160),
.C2(n_162),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_SL g4240 ( 
.A(n_4051),
.B(n_162),
.Y(n_4240)
);

NAND2xp33_ASAP7_75t_SL g4241 ( 
.A(n_4051),
.B(n_164),
.Y(n_4241)
);

AOI22xp5_ASAP7_75t_L g4242 ( 
.A1(n_4036),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4051),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4051),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_4108),
.B(n_165),
.Y(n_4245)
);

AOI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_4056),
.A2(n_167),
.B(n_169),
.Y(n_4246)
);

NAND3xp33_ASAP7_75t_L g4247 ( 
.A(n_4051),
.B(n_170),
.C(n_171),
.Y(n_4247)
);

AOI22xp33_ASAP7_75t_L g4248 ( 
.A1(n_4036),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4051),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4087),
.B(n_174),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4087),
.B(n_175),
.Y(n_4251)
);

OAI21xp5_ASAP7_75t_L g4252 ( 
.A1(n_4056),
.A2(n_177),
.B(n_178),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4051),
.B(n_177),
.Y(n_4253)
);

OAI21xp5_ASAP7_75t_L g4254 ( 
.A1(n_4056),
.A2(n_179),
.B(n_180),
.Y(n_4254)
);

AOI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_4036),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_4255)
);

OAI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_4041),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_SL g4257 ( 
.A(n_4051),
.B(n_185),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4051),
.Y(n_4258)
);

NOR3xp33_ASAP7_75t_L g4259 ( 
.A(n_4092),
.B(n_186),
.C(n_187),
.Y(n_4259)
);

INVxp67_ASAP7_75t_SL g4260 ( 
.A(n_4051),
.Y(n_4260)
);

OAI22x1_ASAP7_75t_L g4261 ( 
.A1(n_4051),
.A2(n_189),
.B1(n_190),
.B2(n_188),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4051),
.Y(n_4262)
);

NOR2xp33_ASAP7_75t_L g4263 ( 
.A(n_4108),
.B(n_186),
.Y(n_4263)
);

AOI221xp5_ASAP7_75t_L g4264 ( 
.A1(n_4092),
.A2(n_190),
.B1(n_193),
.B2(n_189),
.C(n_192),
.Y(n_4264)
);

BUFx2_ASAP7_75t_L g4265 ( 
.A(n_4051),
.Y(n_4265)
);

AOI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_4036),
.A2(n_194),
.B1(n_188),
.B2(n_193),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4265),
.Y(n_4267)
);

OAI221xp5_ASAP7_75t_L g4268 ( 
.A1(n_4137),
.A2(n_4147),
.B1(n_4163),
.B2(n_4218),
.C(n_4241),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4210),
.B(n_196),
.Y(n_4269)
);

OAI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_4131),
.A2(n_4260),
.B1(n_4192),
.B2(n_4216),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4232),
.Y(n_4271)
);

AOI211xp5_ASAP7_75t_L g4272 ( 
.A1(n_4134),
.A2(n_199),
.B(n_196),
.C(n_198),
.Y(n_4272)
);

AOI21xp33_ASAP7_75t_SL g4273 ( 
.A1(n_4195),
.A2(n_200),
.B(n_199),
.Y(n_4273)
);

AOI21xp33_ASAP7_75t_L g4274 ( 
.A1(n_4187),
.A2(n_198),
.B(n_200),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4210),
.B(n_201),
.Y(n_4275)
);

INVxp67_ASAP7_75t_L g4276 ( 
.A(n_4118),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4232),
.Y(n_4277)
);

INVx1_ASAP7_75t_SL g4278 ( 
.A(n_4124),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4207),
.Y(n_4279)
);

INVxp67_ASAP7_75t_SL g4280 ( 
.A(n_4117),
.Y(n_4280)
);

NAND4xp25_ASAP7_75t_L g4281 ( 
.A(n_4197),
.B(n_203),
.C(n_201),
.D(n_202),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4208),
.B(n_202),
.Y(n_4282)
);

AOI21xp33_ASAP7_75t_SL g4283 ( 
.A1(n_4229),
.A2(n_206),
.B(n_205),
.Y(n_4283)
);

INVx3_ASAP7_75t_L g4284 ( 
.A(n_4160),
.Y(n_4284)
);

A2O1A1Ixp33_ASAP7_75t_L g4285 ( 
.A1(n_4202),
.A2(n_207),
.B(n_204),
.C(n_206),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4200),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4224),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4225),
.Y(n_4288)
);

INVx1_ASAP7_75t_SL g4289 ( 
.A(n_4226),
.Y(n_4289)
);

INVxp67_ASAP7_75t_L g4290 ( 
.A(n_4127),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4253),
.B(n_207),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4119),
.B(n_4214),
.Y(n_4292)
);

OAI32xp33_ASAP7_75t_L g4293 ( 
.A1(n_4198),
.A2(n_211),
.A3(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_4160),
.B(n_210),
.Y(n_4294)
);

OAI22xp33_ASAP7_75t_L g4295 ( 
.A1(n_4153),
.A2(n_219),
.B1(n_215),
.B2(n_218),
.Y(n_4295)
);

OR2x2_ASAP7_75t_L g4296 ( 
.A(n_4121),
.B(n_215),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4150),
.B(n_219),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4132),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4166),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4154),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4204),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_4211),
.B(n_4212),
.Y(n_4302)
);

OAI21xp5_ASAP7_75t_SL g4303 ( 
.A1(n_4213),
.A2(n_221),
.B(n_222),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4146),
.Y(n_4304)
);

OAI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_4246),
.A2(n_222),
.B(n_223),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_4141),
.B(n_223),
.Y(n_4306)
);

AO22x1_ASAP7_75t_L g4307 ( 
.A1(n_4252),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4220),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4221),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4222),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4233),
.B(n_227),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4243),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4193),
.Y(n_4313)
);

AOI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_4159),
.A2(n_231),
.B1(n_227),
.B2(n_230),
.Y(n_4314)
);

AOI22xp33_ASAP7_75t_L g4315 ( 
.A1(n_4215),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_4261),
.Y(n_4316)
);

OAI21xp33_ASAP7_75t_L g4317 ( 
.A1(n_4244),
.A2(n_232),
.B(n_234),
.Y(n_4317)
);

NOR2x1_ASAP7_75t_L g4318 ( 
.A(n_4209),
.B(n_234),
.Y(n_4318)
);

OAI22xp5_ASAP7_75t_L g4319 ( 
.A1(n_4152),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4249),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4258),
.B(n_235),
.Y(n_4321)
);

AOI21xp33_ASAP7_75t_L g4322 ( 
.A1(n_4169),
.A2(n_237),
.B(n_238),
.Y(n_4322)
);

NAND4xp25_ASAP7_75t_SL g4323 ( 
.A(n_4262),
.B(n_242),
.C(n_243),
.D(n_241),
.Y(n_4323)
);

AOI222xp33_ASAP7_75t_L g4324 ( 
.A1(n_4179),
.A2(n_244),
.B1(n_246),
.B2(n_240),
.C1(n_243),
.C2(n_245),
.Y(n_4324)
);

INVxp67_ASAP7_75t_L g4325 ( 
.A(n_4120),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4126),
.Y(n_4326)
);

OAI22xp33_ASAP7_75t_SL g4327 ( 
.A1(n_4122),
.A2(n_247),
.B1(n_244),
.B2(n_246),
.Y(n_4327)
);

AO32x1_ASAP7_75t_L g4328 ( 
.A1(n_4140),
.A2(n_249),
.A3(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_4328)
);

NOR2xp33_ASAP7_75t_L g4329 ( 
.A(n_4145),
.B(n_248),
.Y(n_4329)
);

INVxp67_ASAP7_75t_L g4330 ( 
.A(n_4245),
.Y(n_4330)
);

OAI22xp33_ASAP7_75t_L g4331 ( 
.A1(n_4151),
.A2(n_252),
.B1(n_249),
.B2(n_251),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4219),
.B(n_253),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4128),
.Y(n_4333)
);

OAI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_4133),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4227),
.B(n_254),
.Y(n_4335)
);

OAI22xp5_ASAP7_75t_L g4336 ( 
.A1(n_4237),
.A2(n_259),
.B1(n_255),
.B2(n_258),
.Y(n_4336)
);

OAI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4236),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4205),
.Y(n_4338)
);

AOI21xp33_ASAP7_75t_L g4339 ( 
.A1(n_4191),
.A2(n_260),
.B(n_261),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4217),
.Y(n_4340)
);

AOI32xp33_ASAP7_75t_L g4341 ( 
.A1(n_4228),
.A2(n_263),
.A3(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_4341)
);

OAI31xp33_ASAP7_75t_L g4342 ( 
.A1(n_4130),
.A2(n_264),
.A3(n_262),
.B(n_263),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4231),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4240),
.B(n_265),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_4247),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_4345)
);

AOI22xp33_ASAP7_75t_SL g4346 ( 
.A1(n_4162),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_4346)
);

OR2x2_ASAP7_75t_L g4347 ( 
.A(n_4234),
.B(n_269),
.Y(n_4347)
);

OAI21xp33_ASAP7_75t_L g4348 ( 
.A1(n_4156),
.A2(n_4149),
.B(n_4183),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4230),
.B(n_270),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_4123),
.B(n_270),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4257),
.B(n_271),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4139),
.B(n_4135),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_SL g4353 ( 
.A(n_4254),
.B(n_272),
.Y(n_4353)
);

NAND2xp33_ASAP7_75t_SL g4354 ( 
.A(n_4143),
.B(n_274),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4176),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4238),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4164),
.B(n_275),
.Y(n_4357)
);

OAI221xp5_ASAP7_75t_SL g4358 ( 
.A1(n_4158),
.A2(n_279),
.B1(n_276),
.B2(n_278),
.C(n_280),
.Y(n_4358)
);

INVx1_ASAP7_75t_SL g4359 ( 
.A(n_4186),
.Y(n_4359)
);

AND2x2_ASAP7_75t_SL g4360 ( 
.A(n_4259),
.B(n_276),
.Y(n_4360)
);

OAI221xp5_ASAP7_75t_SL g4361 ( 
.A1(n_4174),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.C(n_284),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_4157),
.B(n_281),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_4171),
.B(n_282),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4144),
.B(n_284),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4250),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4256),
.B(n_285),
.Y(n_4366)
);

OAI32xp33_ASAP7_75t_L g4367 ( 
.A1(n_4172),
.A2(n_287),
.A3(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_4367)
);

OAI21xp33_ASAP7_75t_L g4368 ( 
.A1(n_4185),
.A2(n_289),
.B(n_291),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4251),
.Y(n_4369)
);

AOI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_4165),
.A2(n_292),
.B1(n_289),
.B2(n_291),
.Y(n_4370)
);

OAI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_4242),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4371)
);

OAI222xp33_ASAP7_75t_L g4372 ( 
.A1(n_4173),
.A2(n_297),
.B1(n_301),
.B2(n_294),
.C1(n_296),
.C2(n_299),
.Y(n_4372)
);

NOR2xp67_ASAP7_75t_L g4373 ( 
.A(n_4223),
.B(n_296),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4239),
.B(n_303),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4138),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4178),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4177),
.B(n_304),
.Y(n_4377)
);

OAI21xp33_ASAP7_75t_L g4378 ( 
.A1(n_4188),
.A2(n_306),
.B(n_307),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_4199),
.B(n_307),
.Y(n_4379)
);

AOI21x1_ASAP7_75t_L g4380 ( 
.A1(n_4155),
.A2(n_4175),
.B(n_4136),
.Y(n_4380)
);

AOI22xp33_ASAP7_75t_SL g4381 ( 
.A1(n_4201),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4248),
.B(n_4235),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4190),
.Y(n_4383)
);

OAI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4266),
.A2(n_313),
.B1(n_309),
.B2(n_312),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4189),
.Y(n_4385)
);

AOI21xp33_ASAP7_75t_L g4386 ( 
.A1(n_4268),
.A2(n_4194),
.B(n_4129),
.Y(n_4386)
);

OAI221xp5_ASAP7_75t_L g4387 ( 
.A1(n_4289),
.A2(n_4354),
.B1(n_4313),
.B2(n_4316),
.C(n_4290),
.Y(n_4387)
);

NOR3xp33_ASAP7_75t_L g4388 ( 
.A(n_4348),
.B(n_4180),
.C(n_4264),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_SL g4389 ( 
.A(n_4278),
.B(n_4170),
.Y(n_4389)
);

AOI221xp5_ASAP7_75t_L g4390 ( 
.A1(n_4382),
.A2(n_4161),
.B1(n_4148),
.B2(n_4203),
.C(n_4142),
.Y(n_4390)
);

AOI22xp5_ASAP7_75t_L g4391 ( 
.A1(n_4383),
.A2(n_4255),
.B1(n_4263),
.B2(n_4206),
.Y(n_4391)
);

AOI211xp5_ASAP7_75t_SL g4392 ( 
.A1(n_4270),
.A2(n_4125),
.B(n_4184),
.C(n_4181),
.Y(n_4392)
);

AOI21xp33_ASAP7_75t_L g4393 ( 
.A1(n_4292),
.A2(n_4168),
.B(n_4167),
.Y(n_4393)
);

OAI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4279),
.A2(n_4182),
.B1(n_4196),
.B2(n_314),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4328),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_4328),
.A2(n_314),
.B(n_313),
.Y(n_4396)
);

NAND3xp33_ASAP7_75t_L g4397 ( 
.A(n_4272),
.B(n_312),
.C(n_315),
.Y(n_4397)
);

AOI21xp5_ASAP7_75t_L g4398 ( 
.A1(n_4328),
.A2(n_317),
.B(n_316),
.Y(n_4398)
);

AOI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_4385),
.A2(n_325),
.B1(n_336),
.B2(n_315),
.Y(n_4399)
);

NOR3xp33_ASAP7_75t_L g4400 ( 
.A(n_4359),
.B(n_4284),
.C(n_4330),
.Y(n_4400)
);

AOI322xp5_ASAP7_75t_L g4401 ( 
.A1(n_4376),
.A2(n_4318),
.A3(n_4375),
.B1(n_4352),
.B2(n_4335),
.C1(n_4349),
.C2(n_4360),
.Y(n_4401)
);

OAI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4276),
.A2(n_4280),
.B(n_4373),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4284),
.B(n_317),
.Y(n_4403)
);

OR4x1_ASAP7_75t_L g4404 ( 
.A(n_4271),
.B(n_320),
.C(n_318),
.D(n_319),
.Y(n_4404)
);

OAI31xp33_ASAP7_75t_L g4405 ( 
.A1(n_4285),
.A2(n_324),
.A3(n_321),
.B(n_322),
.Y(n_4405)
);

AOI211x1_ASAP7_75t_L g4406 ( 
.A1(n_4277),
.A2(n_326),
.B(n_322),
.C(n_324),
.Y(n_4406)
);

AOI221xp5_ASAP7_75t_L g4407 ( 
.A1(n_4333),
.A2(n_4343),
.B1(n_4356),
.B2(n_4340),
.C(n_4338),
.Y(n_4407)
);

OAI221xp5_ASAP7_75t_SL g4408 ( 
.A1(n_4286),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4307),
.B(n_329),
.Y(n_4409)
);

OAI21xp33_ASAP7_75t_L g4410 ( 
.A1(n_4267),
.A2(n_332),
.B(n_333),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4298),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_4411)
);

AOI221xp5_ASAP7_75t_L g4412 ( 
.A1(n_4365),
.A2(n_361),
.B1(n_370),
.B2(n_351),
.C(n_339),
.Y(n_4412)
);

NAND4xp25_ASAP7_75t_L g4413 ( 
.A(n_4302),
.B(n_345),
.C(n_341),
.D(n_342),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_SL g4414 ( 
.A(n_4273),
.B(n_341),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4326),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_4415)
);

OAI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4296),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_4323),
.A2(n_355),
.B(n_353),
.Y(n_4417)
);

INVxp67_ASAP7_75t_L g4418 ( 
.A(n_4269),
.Y(n_4418)
);

AOI211xp5_ASAP7_75t_SL g4419 ( 
.A1(n_4301),
.A2(n_4308),
.B(n_4310),
.C(n_4309),
.Y(n_4419)
);

NOR3xp33_ASAP7_75t_L g4420 ( 
.A(n_4339),
.B(n_352),
.C(n_353),
.Y(n_4420)
);

HB1xp67_ASAP7_75t_L g4421 ( 
.A(n_4287),
.Y(n_4421)
);

OAI21xp33_ASAP7_75t_L g4422 ( 
.A1(n_4288),
.A2(n_4302),
.B(n_4312),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_4283),
.B(n_352),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4275),
.Y(n_4424)
);

NOR2xp33_ASAP7_75t_L g4425 ( 
.A(n_4281),
.B(n_4327),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4346),
.B(n_4299),
.Y(n_4426)
);

OAI311xp33_ASAP7_75t_L g4427 ( 
.A1(n_4320),
.A2(n_358),
.A3(n_356),
.B1(n_357),
.C1(n_359),
.Y(n_4427)
);

NOR3xp33_ASAP7_75t_L g4428 ( 
.A(n_4325),
.B(n_356),
.C(n_357),
.Y(n_4428)
);

OAI21xp33_ASAP7_75t_L g4429 ( 
.A1(n_4369),
.A2(n_362),
.B(n_363),
.Y(n_4429)
);

AOI211xp5_ASAP7_75t_SL g4430 ( 
.A1(n_4358),
.A2(n_4317),
.B(n_4303),
.C(n_4361),
.Y(n_4430)
);

NOR3xp33_ASAP7_75t_L g4431 ( 
.A(n_4322),
.B(n_364),
.C(n_365),
.Y(n_4431)
);

NAND3xp33_ASAP7_75t_L g4432 ( 
.A(n_4304),
.B(n_365),
.C(n_366),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4291),
.Y(n_4433)
);

AOI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_4353),
.A2(n_4355),
.B1(n_4300),
.B2(n_4379),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4364),
.Y(n_4435)
);

OAI22xp5_ASAP7_75t_L g4436 ( 
.A1(n_4350),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_4436)
);

NAND3xp33_ASAP7_75t_SL g4437 ( 
.A(n_4342),
.B(n_367),
.C(n_370),
.Y(n_4437)
);

AOI221xp5_ASAP7_75t_L g4438 ( 
.A1(n_4305),
.A2(n_4367),
.B1(n_4374),
.B2(n_4384),
.C(n_4337),
.Y(n_4438)
);

A2O1A1Ixp33_ASAP7_75t_L g4439 ( 
.A1(n_4341),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_4311),
.B(n_4321),
.Y(n_4440)
);

OAI21xp5_ASAP7_75t_SL g4441 ( 
.A1(n_4329),
.A2(n_373),
.B(n_376),
.Y(n_4441)
);

A2O1A1Ixp33_ASAP7_75t_L g4442 ( 
.A1(n_4297),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_4442)
);

NOR4xp75_ASAP7_75t_SL g4443 ( 
.A(n_4336),
.B(n_379),
.C(n_377),
.D(n_378),
.Y(n_4443)
);

OAI221xp5_ASAP7_75t_L g4444 ( 
.A1(n_4381),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.C(n_383),
.Y(n_4444)
);

AOI22xp5_ASAP7_75t_L g4445 ( 
.A1(n_4378),
.A2(n_394),
.B1(n_404),
.B2(n_380),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4324),
.B(n_381),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4294),
.Y(n_4447)
);

AOI211xp5_ASAP7_75t_L g4448 ( 
.A1(n_4345),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_4448)
);

AOI221xp5_ASAP7_75t_L g4449 ( 
.A1(n_4371),
.A2(n_409),
.B1(n_418),
.B2(n_398),
.C(n_384),
.Y(n_4449)
);

OAI211xp5_ASAP7_75t_SL g4450 ( 
.A1(n_4368),
.A2(n_4357),
.B(n_4315),
.C(n_4366),
.Y(n_4450)
);

NOR2xp33_ASAP7_75t_L g4451 ( 
.A(n_4293),
.B(n_385),
.Y(n_4451)
);

NOR2xp33_ASAP7_75t_L g4452 ( 
.A(n_4282),
.B(n_390),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4332),
.B(n_391),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4344),
.B(n_391),
.Y(n_4454)
);

NAND3xp33_ASAP7_75t_SL g4455 ( 
.A(n_4306),
.B(n_392),
.C(n_395),
.Y(n_4455)
);

OAI22x1_ASAP7_75t_L g4456 ( 
.A1(n_4314),
.A2(n_400),
.B1(n_396),
.B2(n_397),
.Y(n_4456)
);

XOR2xp5_ASAP7_75t_L g4457 ( 
.A(n_4380),
.B(n_401),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4363),
.Y(n_4458)
);

AOI221xp5_ASAP7_75t_L g4459 ( 
.A1(n_4274),
.A2(n_422),
.B1(n_431),
.B2(n_414),
.C(n_403),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4377),
.Y(n_4460)
);

OAI21xp5_ASAP7_75t_SL g4461 ( 
.A1(n_4372),
.A2(n_4351),
.B(n_4370),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4347),
.Y(n_4462)
);

AOI221xp5_ASAP7_75t_L g4463 ( 
.A1(n_4362),
.A2(n_422),
.B1(n_432),
.B2(n_414),
.C(n_403),
.Y(n_4463)
);

O2A1O1Ixp33_ASAP7_75t_SL g4464 ( 
.A1(n_4295),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_4464)
);

AOI222xp33_ASAP7_75t_L g4465 ( 
.A1(n_4319),
.A2(n_408),
.B1(n_412),
.B2(n_406),
.C1(n_407),
.C2(n_410),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4331),
.B(n_410),
.Y(n_4466)
);

AOI211xp5_ASAP7_75t_L g4467 ( 
.A1(n_4334),
.A2(n_415),
.B(n_412),
.C(n_413),
.Y(n_4467)
);

OR3x1_ASAP7_75t_L g4468 ( 
.A(n_4267),
.B(n_413),
.C(n_415),
.Y(n_4468)
);

AOI322xp5_ASAP7_75t_L g4469 ( 
.A1(n_4359),
.A2(n_421),
.A3(n_420),
.B1(n_418),
.B2(n_416),
.C1(n_417),
.C2(n_419),
.Y(n_4469)
);

OAI32xp33_ASAP7_75t_L g4470 ( 
.A1(n_4278),
.A2(n_424),
.A3(n_416),
.B1(n_423),
.B2(n_425),
.Y(n_4470)
);

NAND3xp33_ASAP7_75t_SL g4471 ( 
.A(n_4278),
.B(n_427),
.C(n_428),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4278),
.B(n_429),
.Y(n_4472)
);

OAI322xp33_ASAP7_75t_L g4473 ( 
.A1(n_4268),
.A2(n_438),
.A3(n_437),
.B1(n_434),
.B2(n_430),
.C1(n_433),
.C2(n_435),
.Y(n_4473)
);

AOI211xp5_ASAP7_75t_L g4474 ( 
.A1(n_4268),
.A2(n_438),
.B(n_430),
.C(n_435),
.Y(n_4474)
);

NAND2x1_ASAP7_75t_L g4475 ( 
.A(n_4279),
.B(n_439),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4284),
.Y(n_4476)
);

A2O1A1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_4268),
.A2(n_442),
.B(n_439),
.C(n_440),
.Y(n_4477)
);

OAI21x1_ASAP7_75t_L g4478 ( 
.A1(n_4284),
.A2(n_440),
.B(n_442),
.Y(n_4478)
);

OAI321xp33_ASAP7_75t_L g4479 ( 
.A1(n_4268),
.A2(n_445),
.A3(n_447),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_4479)
);

AOI211xp5_ASAP7_75t_L g4480 ( 
.A1(n_4268),
.A2(n_447),
.B(n_444),
.C(n_445),
.Y(n_4480)
);

A2O1A1Ixp33_ASAP7_75t_L g4481 ( 
.A1(n_4268),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4284),
.B(n_449),
.Y(n_4482)
);

INVx1_ASAP7_75t_SL g4483 ( 
.A(n_4278),
.Y(n_4483)
);

AOI221xp5_ASAP7_75t_L g4484 ( 
.A1(n_4268),
.A2(n_469),
.B1(n_479),
.B2(n_459),
.C(n_451),
.Y(n_4484)
);

NAND4xp25_ASAP7_75t_L g4485 ( 
.A(n_4278),
.B(n_454),
.C(n_452),
.D(n_453),
.Y(n_4485)
);

OAI22xp5_ASAP7_75t_L g4486 ( 
.A1(n_4278),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_4486)
);

INVxp67_ASAP7_75t_L g4487 ( 
.A(n_4268),
.Y(n_4487)
);

AOI21xp5_ASAP7_75t_L g4488 ( 
.A1(n_4268),
.A2(n_459),
.B(n_458),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4328),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_SL g4490 ( 
.A(n_4278),
.B(n_456),
.Y(n_4490)
);

OAI21xp33_ASAP7_75t_L g4491 ( 
.A1(n_4278),
.A2(n_460),
.B(n_461),
.Y(n_4491)
);

AOI21xp5_ASAP7_75t_L g4492 ( 
.A1(n_4268),
.A2(n_464),
.B(n_463),
.Y(n_4492)
);

AOI211xp5_ASAP7_75t_L g4493 ( 
.A1(n_4268),
.A2(n_465),
.B(n_460),
.C(n_464),
.Y(n_4493)
);

AOI32xp33_ASAP7_75t_L g4494 ( 
.A1(n_4268),
.A2(n_468),
.A3(n_465),
.B1(n_466),
.B2(n_469),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4284),
.B(n_466),
.Y(n_4495)
);

NOR2x1_ASAP7_75t_L g4496 ( 
.A(n_4278),
.B(n_468),
.Y(n_4496)
);

OAI321xp33_ASAP7_75t_L g4497 ( 
.A1(n_4268),
.A2(n_472),
.A3(n_475),
.B1(n_470),
.B2(n_471),
.C(n_474),
.Y(n_4497)
);

AOI211xp5_ASAP7_75t_L g4498 ( 
.A1(n_4268),
.A2(n_474),
.B(n_471),
.C(n_472),
.Y(n_4498)
);

NOR3x1_ASAP7_75t_L g4499 ( 
.A(n_4280),
.B(n_477),
.C(n_478),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4383),
.A2(n_486),
.B1(n_495),
.B2(n_477),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4278),
.B(n_478),
.Y(n_4501)
);

NOR4xp75_ASAP7_75t_SL g4502 ( 
.A(n_4270),
.B(n_481),
.C(n_479),
.D(n_480),
.Y(n_4502)
);

OAI211xp5_ASAP7_75t_L g4503 ( 
.A1(n_4280),
.A2(n_483),
.B(n_480),
.C(n_482),
.Y(n_4503)
);

AOI221xp5_ASAP7_75t_L g4504 ( 
.A1(n_4268),
.A2(n_502),
.B1(n_516),
.B2(n_492),
.C(n_482),
.Y(n_4504)
);

OAI21xp5_ASAP7_75t_L g4505 ( 
.A1(n_4278),
.A2(n_483),
.B(n_484),
.Y(n_4505)
);

NOR2xp33_ASAP7_75t_L g4506 ( 
.A(n_4278),
.B(n_486),
.Y(n_4506)
);

NAND4xp75_ASAP7_75t_L g4507 ( 
.A(n_4267),
.B(n_489),
.C(n_487),
.D(n_488),
.Y(n_4507)
);

NAND3xp33_ASAP7_75t_L g4508 ( 
.A(n_4272),
.B(n_487),
.C(n_491),
.Y(n_4508)
);

AOI221xp5_ASAP7_75t_L g4509 ( 
.A1(n_4268),
.A2(n_516),
.B1(n_525),
.B2(n_502),
.C(n_492),
.Y(n_4509)
);

OA21x2_ASAP7_75t_L g4510 ( 
.A1(n_4348),
.A2(n_493),
.B(n_494),
.Y(n_4510)
);

AOI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_4383),
.A2(n_496),
.B1(n_493),
.B2(n_495),
.Y(n_4511)
);

OAI22xp33_ASAP7_75t_L g4512 ( 
.A1(n_4268),
.A2(n_500),
.B1(n_496),
.B2(n_497),
.Y(n_4512)
);

AOI221xp5_ASAP7_75t_L g4513 ( 
.A1(n_4268),
.A2(n_503),
.B1(n_497),
.B2(n_501),
.C(n_505),
.Y(n_4513)
);

AOI211xp5_ASAP7_75t_L g4514 ( 
.A1(n_4268),
.A2(n_510),
.B(n_503),
.C(n_508),
.Y(n_4514)
);

AO21x1_ASAP7_75t_L g4515 ( 
.A1(n_4354),
.A2(n_508),
.B(n_512),
.Y(n_4515)
);

AOI21xp33_ASAP7_75t_L g4516 ( 
.A1(n_4268),
.A2(n_512),
.B(n_513),
.Y(n_4516)
);

AOI22xp5_ASAP7_75t_L g4517 ( 
.A1(n_4383),
.A2(n_517),
.B1(n_513),
.B2(n_514),
.Y(n_4517)
);

AOI221xp5_ASAP7_75t_L g4518 ( 
.A1(n_4268),
.A2(n_518),
.B1(n_514),
.B2(n_517),
.C(n_520),
.Y(n_4518)
);

OAI221xp5_ASAP7_75t_SL g4519 ( 
.A1(n_4268),
.A2(n_521),
.B1(n_518),
.B2(n_520),
.C(n_522),
.Y(n_4519)
);

OAI21xp5_ASAP7_75t_SL g4520 ( 
.A1(n_4278),
.A2(n_521),
.B(n_522),
.Y(n_4520)
);

AOI22xp33_ASAP7_75t_L g4521 ( 
.A1(n_4383),
.A2(n_526),
.B1(n_523),
.B2(n_524),
.Y(n_4521)
);

NAND3xp33_ASAP7_75t_SL g4522 ( 
.A(n_4278),
.B(n_523),
.C(n_524),
.Y(n_4522)
);

NAND4xp75_ASAP7_75t_L g4523 ( 
.A(n_4267),
.B(n_529),
.C(n_527),
.D(n_528),
.Y(n_4523)
);

AOI21xp5_ASAP7_75t_L g4524 ( 
.A1(n_4268),
.A2(n_528),
.B(n_529),
.Y(n_4524)
);

OAI21xp5_ASAP7_75t_SL g4525 ( 
.A1(n_4278),
.A2(n_530),
.B(n_531),
.Y(n_4525)
);

AOI221x1_ASAP7_75t_L g4526 ( 
.A1(n_4270),
.A2(n_533),
.B1(n_530),
.B2(n_531),
.C(n_534),
.Y(n_4526)
);

AOI221xp5_ASAP7_75t_L g4527 ( 
.A1(n_4268),
.A2(n_537),
.B1(n_534),
.B2(n_535),
.C(n_538),
.Y(n_4527)
);

NOR2x1_ASAP7_75t_L g4528 ( 
.A(n_4278),
.B(n_537),
.Y(n_4528)
);

OAI221xp5_ASAP7_75t_L g4529 ( 
.A1(n_4268),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.C(n_541),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4328),
.Y(n_4530)
);

AOI221xp5_ASAP7_75t_L g4531 ( 
.A1(n_4268),
.A2(n_543),
.B1(n_539),
.B2(n_542),
.C(n_544),
.Y(n_4531)
);

AOI221xp5_ASAP7_75t_L g4532 ( 
.A1(n_4268),
.A2(n_545),
.B1(n_542),
.B2(n_544),
.C(n_546),
.Y(n_4532)
);

AO221x1_ASAP7_75t_L g4533 ( 
.A1(n_4284),
.A2(n_548),
.B1(n_545),
.B2(n_546),
.C(n_549),
.Y(n_4533)
);

OAI211xp5_ASAP7_75t_L g4534 ( 
.A1(n_4280),
.A2(n_551),
.B(n_548),
.C(n_550),
.Y(n_4534)
);

OAI221xp5_ASAP7_75t_L g4535 ( 
.A1(n_4487),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.C(n_556),
.Y(n_4535)
);

INVxp67_ASAP7_75t_SL g4536 ( 
.A(n_4496),
.Y(n_4536)
);

OAI22xp5_ASAP7_75t_L g4537 ( 
.A1(n_4483),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_4537)
);

OAI32xp33_ASAP7_75t_L g4538 ( 
.A1(n_4388),
.A2(n_560),
.A3(n_558),
.B1(n_559),
.B2(n_562),
.Y(n_4538)
);

AOI31xp33_ASAP7_75t_L g4539 ( 
.A1(n_4419),
.A2(n_4402),
.A3(n_4421),
.B(n_4422),
.Y(n_4539)
);

INVx1_ASAP7_75t_SL g4540 ( 
.A(n_4468),
.Y(n_4540)
);

O2A1O1Ixp33_ASAP7_75t_L g4541 ( 
.A1(n_4427),
.A2(n_564),
.B(n_559),
.C(n_563),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4533),
.B(n_563),
.Y(n_4542)
);

INVxp67_ASAP7_75t_L g4543 ( 
.A(n_4528),
.Y(n_4543)
);

AOI21xp33_ASAP7_75t_L g4544 ( 
.A1(n_4395),
.A2(n_565),
.B(n_567),
.Y(n_4544)
);

AOI22xp5_ASAP7_75t_SL g4545 ( 
.A1(n_4489),
.A2(n_568),
.B1(n_565),
.B2(n_567),
.Y(n_4545)
);

A2O1A1Ixp33_ASAP7_75t_L g4546 ( 
.A1(n_4530),
.A2(n_571),
.B(n_569),
.C(n_570),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_L g4547 ( 
.A(n_4406),
.B(n_4454),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4499),
.B(n_569),
.Y(n_4548)
);

OAI22xp5_ASAP7_75t_L g4549 ( 
.A1(n_4476),
.A2(n_575),
.B1(n_570),
.B2(n_574),
.Y(n_4549)
);

OAI21xp5_ASAP7_75t_L g4550 ( 
.A1(n_4488),
.A2(n_4524),
.B(n_4492),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4520),
.B(n_4525),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4472),
.B(n_4501),
.Y(n_4552)
);

AOI22xp5_ASAP7_75t_L g4553 ( 
.A1(n_4440),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_4553)
);

OAI22xp5_ASAP7_75t_L g4554 ( 
.A1(n_4506),
.A2(n_4389),
.B1(n_4387),
.B2(n_4519),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4404),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4510),
.Y(n_4556)
);

AND2x4_ASAP7_75t_L g4557 ( 
.A(n_4400),
.B(n_576),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4515),
.B(n_578),
.Y(n_4558)
);

AOI22xp5_ASAP7_75t_L g4559 ( 
.A1(n_4436),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_SL g4560 ( 
.A(n_4502),
.B(n_581),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4526),
.B(n_582),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_SL g4562 ( 
.A(n_4443),
.B(n_4390),
.Y(n_4562)
);

NAND3xp33_ASAP7_75t_SL g4563 ( 
.A(n_4474),
.B(n_583),
.C(n_584),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4457),
.Y(n_4564)
);

OAI21xp33_ASAP7_75t_L g4565 ( 
.A1(n_4425),
.A2(n_583),
.B(n_584),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4510),
.B(n_585),
.Y(n_4566)
);

INVx1_ASAP7_75t_SL g4567 ( 
.A(n_4475),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4423),
.Y(n_4568)
);

AOI22xp5_ASAP7_75t_L g4569 ( 
.A1(n_4471),
.A2(n_588),
.B1(n_585),
.B2(n_587),
.Y(n_4569)
);

OAI21xp33_ASAP7_75t_L g4570 ( 
.A1(n_4494),
.A2(n_587),
.B(n_589),
.Y(n_4570)
);

AOI21xp5_ASAP7_75t_L g4571 ( 
.A1(n_4490),
.A2(n_591),
.B(n_592),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_4464),
.A2(n_591),
.B(n_593),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4414),
.A2(n_593),
.B(n_594),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4435),
.B(n_595),
.Y(n_4574)
);

OAI21xp5_ASAP7_75t_SL g4575 ( 
.A1(n_4392),
.A2(n_595),
.B(n_596),
.Y(n_4575)
);

OAI221xp5_ASAP7_75t_L g4576 ( 
.A1(n_4461),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.C(n_600),
.Y(n_4576)
);

BUFx6f_ASAP7_75t_L g4577 ( 
.A(n_4403),
.Y(n_4577)
);

AOI322xp5_ASAP7_75t_L g4578 ( 
.A1(n_4512),
.A2(n_4516),
.A3(n_4438),
.B1(n_4437),
.B2(n_4391),
.C1(n_4513),
.C2(n_4509),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4482),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4529),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_4580)
);

NOR4xp25_ASAP7_75t_L g4581 ( 
.A(n_4477),
.B(n_602),
.C(n_600),
.D(n_601),
.Y(n_4581)
);

OAI221xp5_ASAP7_75t_L g4582 ( 
.A1(n_4505),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.C(n_605),
.Y(n_4582)
);

AOI221xp5_ASAP7_75t_L g4583 ( 
.A1(n_4479),
.A2(n_607),
.B1(n_603),
.B2(n_605),
.C(n_608),
.Y(n_4583)
);

XNOR2x1_ASAP7_75t_L g4584 ( 
.A(n_4456),
.B(n_607),
.Y(n_4584)
);

CKINVDCx20_ASAP7_75t_R g4585 ( 
.A(n_4434),
.Y(n_4585)
);

OAI221xp5_ASAP7_75t_L g4586 ( 
.A1(n_4441),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.C(n_611),
.Y(n_4586)
);

AOI22xp5_ASAP7_75t_L g4587 ( 
.A1(n_4522),
.A2(n_614),
.B1(n_609),
.B2(n_612),
.Y(n_4587)
);

INVx1_ASAP7_75t_SL g4588 ( 
.A(n_4507),
.Y(n_4588)
);

NAND4xp25_ASAP7_75t_L g4589 ( 
.A(n_4430),
.B(n_616),
.C(n_612),
.D(n_615),
.Y(n_4589)
);

AOI31xp33_ASAP7_75t_L g4590 ( 
.A1(n_4480),
.A2(n_618),
.A3(n_616),
.B(n_617),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4495),
.Y(n_4591)
);

OAI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_4481),
.A2(n_4417),
.B(n_4497),
.Y(n_4592)
);

INVx2_ASAP7_75t_SL g4593 ( 
.A(n_4478),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4453),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4460),
.Y(n_4595)
);

A2O1A1Ixp33_ASAP7_75t_L g4596 ( 
.A1(n_4452),
.A2(n_620),
.B(n_618),
.C(n_619),
.Y(n_4596)
);

AOI22xp33_ASAP7_75t_SL g4597 ( 
.A1(n_4458),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_4597)
);

AOI221x1_ASAP7_75t_L g4598 ( 
.A1(n_4386),
.A2(n_623),
.B1(n_621),
.B2(n_622),
.C(n_624),
.Y(n_4598)
);

OAI322xp33_ASAP7_75t_L g4599 ( 
.A1(n_4426),
.A2(n_628),
.A3(n_627),
.B1(n_624),
.B2(n_622),
.C1(n_623),
.C2(n_625),
.Y(n_4599)
);

INVx3_ASAP7_75t_L g4600 ( 
.A(n_4523),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4462),
.B(n_625),
.Y(n_4601)
);

AOI22xp33_ASAP7_75t_L g4602 ( 
.A1(n_4433),
.A2(n_630),
.B1(n_627),
.B2(n_629),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4410),
.B(n_629),
.Y(n_4603)
);

NOR2x1_ASAP7_75t_L g4604 ( 
.A(n_4413),
.B(n_631),
.Y(n_4604)
);

OAI21xp33_ASAP7_75t_SL g4605 ( 
.A1(n_4401),
.A2(n_632),
.B(n_634),
.Y(n_4605)
);

INVxp67_ASAP7_75t_L g4606 ( 
.A(n_4451),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4469),
.B(n_632),
.Y(n_4607)
);

AOI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_4396),
.A2(n_635),
.B(n_636),
.Y(n_4608)
);

AOI21xp33_ASAP7_75t_L g4609 ( 
.A1(n_4418),
.A2(n_635),
.B(n_637),
.Y(n_4609)
);

O2A1O1Ixp33_ASAP7_75t_L g4610 ( 
.A1(n_4473),
.A2(n_639),
.B(n_637),
.C(n_638),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4465),
.B(n_638),
.Y(n_4611)
);

AOI21xp33_ASAP7_75t_L g4612 ( 
.A1(n_4394),
.A2(n_641),
.B(n_642),
.Y(n_4612)
);

AOI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4424),
.A2(n_645),
.B1(n_643),
.B2(n_644),
.Y(n_4613)
);

NAND4xp25_ASAP7_75t_L g4614 ( 
.A(n_4493),
.B(n_645),
.C(n_643),
.D(n_644),
.Y(n_4614)
);

AOI21xp5_ASAP7_75t_L g4615 ( 
.A1(n_4398),
.A2(n_647),
.B(n_648),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4446),
.Y(n_4616)
);

OAI21xp5_ASAP7_75t_SL g4617 ( 
.A1(n_4484),
.A2(n_648),
.B(n_649),
.Y(n_4617)
);

AOI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4485),
.A2(n_653),
.B1(n_651),
.B2(n_652),
.Y(n_4618)
);

AOI221xp5_ASAP7_75t_L g4619 ( 
.A1(n_4450),
.A2(n_654),
.B1(n_651),
.B2(n_652),
.C(n_656),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_4409),
.Y(n_4620)
);

INVxp67_ASAP7_75t_L g4621 ( 
.A(n_4455),
.Y(n_4621)
);

AOI322xp5_ASAP7_75t_L g4622 ( 
.A1(n_4504),
.A2(n_654),
.A3(n_657),
.B1(n_658),
.B2(n_659),
.C1(n_660),
.C2(n_661),
.Y(n_4622)
);

NAND3xp33_ASAP7_75t_SL g4623 ( 
.A(n_4585),
.B(n_4514),
.C(n_4498),
.Y(n_4623)
);

OAI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4605),
.A2(n_4508),
.B(n_4397),
.Y(n_4624)
);

NOR2xp67_ASAP7_75t_L g4625 ( 
.A(n_4555),
.B(n_4486),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4577),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4556),
.Y(n_4627)
);

AOI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4616),
.A2(n_4447),
.B1(n_4420),
.B2(n_4431),
.Y(n_4628)
);

INVx1_ASAP7_75t_SL g4629 ( 
.A(n_4540),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4577),
.Y(n_4630)
);

INVx1_ASAP7_75t_SL g4631 ( 
.A(n_4547),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4620),
.A2(n_4491),
.B1(n_4527),
.B2(n_4518),
.Y(n_4632)
);

NAND5xp2_ASAP7_75t_L g4633 ( 
.A(n_4575),
.B(n_4407),
.C(n_4532),
.D(n_4531),
.E(n_4405),
.Y(n_4633)
);

OAI31xp33_ASAP7_75t_L g4634 ( 
.A1(n_4567),
.A2(n_4503),
.A3(n_4534),
.B(n_4442),
.Y(n_4634)
);

O2A1O1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4539),
.A2(n_4439),
.B(n_4428),
.C(n_4470),
.Y(n_4635)
);

AOI322xp5_ASAP7_75t_L g4636 ( 
.A1(n_4536),
.A2(n_4429),
.A3(n_4393),
.B1(n_4459),
.B2(n_4466),
.C1(n_4463),
.C2(n_4511),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4543),
.Y(n_4637)
);

AOI21xp5_ASAP7_75t_L g4638 ( 
.A1(n_4562),
.A2(n_4444),
.B(n_4416),
.Y(n_4638)
);

AOI221xp5_ASAP7_75t_L g4639 ( 
.A1(n_4541),
.A2(n_4544),
.B1(n_4564),
.B2(n_4554),
.C(n_4572),
.Y(n_4639)
);

OAI221xp5_ASAP7_75t_L g4640 ( 
.A1(n_4551),
.A2(n_4615),
.B1(n_4608),
.B2(n_4592),
.C(n_4606),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4566),
.Y(n_4641)
);

A2O1A1Ixp33_ASAP7_75t_L g4642 ( 
.A1(n_4545),
.A2(n_4432),
.B(n_4445),
.C(n_4500),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4558),
.Y(n_4643)
);

OAI21xp5_ASAP7_75t_SL g4644 ( 
.A1(n_4557),
.A2(n_4517),
.B(n_4399),
.Y(n_4644)
);

OAI321xp33_ASAP7_75t_L g4645 ( 
.A1(n_4593),
.A2(n_4408),
.A3(n_4448),
.B1(n_4467),
.B2(n_4521),
.C(n_4411),
.Y(n_4645)
);

OAI321xp33_ASAP7_75t_L g4646 ( 
.A1(n_4621),
.A2(n_4550),
.A3(n_4552),
.B1(n_4568),
.B2(n_4595),
.C(n_4594),
.Y(n_4646)
);

AOI221x1_ASAP7_75t_L g4647 ( 
.A1(n_4612),
.A2(n_4557),
.B1(n_4589),
.B2(n_4546),
.C(n_4565),
.Y(n_4647)
);

OAI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4604),
.A2(n_4415),
.B(n_4449),
.Y(n_4648)
);

BUFx2_ASAP7_75t_L g4649 ( 
.A(n_4600),
.Y(n_4649)
);

AOI322xp5_ASAP7_75t_L g4650 ( 
.A1(n_4588),
.A2(n_4412),
.A3(n_659),
.B1(n_660),
.B2(n_661),
.C1(n_662),
.C2(n_663),
.Y(n_4650)
);

INVx1_ASAP7_75t_SL g4651 ( 
.A(n_4584),
.Y(n_4651)
);

AOI221xp5_ASAP7_75t_SL g4652 ( 
.A1(n_4570),
.A2(n_664),
.B1(n_658),
.B2(n_663),
.C(n_665),
.Y(n_4652)
);

AOI221xp5_ASAP7_75t_L g4653 ( 
.A1(n_4610),
.A2(n_667),
.B1(n_664),
.B2(n_666),
.C(n_668),
.Y(n_4653)
);

CKINVDCx20_ASAP7_75t_R g4654 ( 
.A(n_4600),
.Y(n_4654)
);

INVxp67_ASAP7_75t_SL g4655 ( 
.A(n_4560),
.Y(n_4655)
);

OAI22xp5_ASAP7_75t_L g4656 ( 
.A1(n_4542),
.A2(n_669),
.B1(n_666),
.B2(n_668),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4561),
.Y(n_4657)
);

INVxp67_ASAP7_75t_L g4658 ( 
.A(n_4548),
.Y(n_4658)
);

OAI22xp33_ASAP7_75t_L g4659 ( 
.A1(n_4569),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.Y(n_4659)
);

XNOR2x1_ASAP7_75t_L g4660 ( 
.A(n_4618),
.B(n_671),
.Y(n_4660)
);

AOI221xp5_ASAP7_75t_L g4661 ( 
.A1(n_4581),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.C(n_676),
.Y(n_4661)
);

AND2x4_ASAP7_75t_L g4662 ( 
.A(n_4574),
.B(n_673),
.Y(n_4662)
);

AOI32xp33_ASAP7_75t_L g4663 ( 
.A1(n_4579),
.A2(n_678),
.A3(n_676),
.B1(n_677),
.B2(n_680),
.Y(n_4663)
);

XNOR2x1_ASAP7_75t_L g4664 ( 
.A(n_4587),
.B(n_678),
.Y(n_4664)
);

AOI21xp33_ASAP7_75t_L g4665 ( 
.A1(n_4591),
.A2(n_680),
.B(n_682),
.Y(n_4665)
);

OAI21xp33_ASAP7_75t_L g4666 ( 
.A1(n_4578),
.A2(n_683),
.B(n_684),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4603),
.B(n_685),
.Y(n_4667)
);

AOI322xp5_ASAP7_75t_L g4668 ( 
.A1(n_4563),
.A2(n_4611),
.A3(n_4607),
.B1(n_4577),
.B2(n_4601),
.C1(n_4583),
.C2(n_4619),
.Y(n_4668)
);

AOI21xp33_ASAP7_75t_L g4669 ( 
.A1(n_4590),
.A2(n_689),
.B(n_691),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4598),
.B(n_689),
.Y(n_4670)
);

OAI21xp5_ASAP7_75t_SL g4671 ( 
.A1(n_4617),
.A2(n_692),
.B(n_693),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4599),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4614),
.Y(n_4673)
);

O2A1O1Ixp5_ASAP7_75t_L g4674 ( 
.A1(n_4538),
.A2(n_696),
.B(n_694),
.C(n_695),
.Y(n_4674)
);

AOI221xp5_ASAP7_75t_L g4675 ( 
.A1(n_4573),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.C(n_699),
.Y(n_4675)
);

XNOR2xp5_ASAP7_75t_L g4676 ( 
.A(n_4537),
.B(n_697),
.Y(n_4676)
);

AOI22xp33_ASAP7_75t_SL g4677 ( 
.A1(n_4580),
.A2(n_701),
.B1(n_699),
.B2(n_700),
.Y(n_4677)
);

INVx1_ASAP7_75t_SL g4678 ( 
.A(n_4597),
.Y(n_4678)
);

AOI221xp5_ASAP7_75t_L g4679 ( 
.A1(n_4571),
.A2(n_702),
.B1(n_700),
.B2(n_701),
.C(n_703),
.Y(n_4679)
);

OAI22xp5_ASAP7_75t_L g4680 ( 
.A1(n_4576),
.A2(n_707),
.B1(n_704),
.B2(n_706),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4655),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4627),
.Y(n_4682)
);

INVx1_ASAP7_75t_SL g4683 ( 
.A(n_4654),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4662),
.B(n_4596),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4662),
.B(n_4622),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4649),
.B(n_4626),
.Y(n_4686)
);

AOI22xp5_ASAP7_75t_L g4687 ( 
.A1(n_4631),
.A2(n_4582),
.B1(n_4559),
.B2(n_4586),
.Y(n_4687)
);

XNOR2xp5_ASAP7_75t_L g4688 ( 
.A(n_4623),
.B(n_4553),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4674),
.Y(n_4689)
);

AOI211x1_ASAP7_75t_SL g4690 ( 
.A1(n_4625),
.A2(n_4549),
.B(n_4609),
.C(n_4535),
.Y(n_4690)
);

AOI322xp5_ASAP7_75t_L g4691 ( 
.A1(n_4629),
.A2(n_4602),
.A3(n_4613),
.B1(n_709),
.B2(n_710),
.C1(n_712),
.C2(n_713),
.Y(n_4691)
);

AOI22xp33_ASAP7_75t_L g4692 ( 
.A1(n_4657),
.A2(n_709),
.B1(n_704),
.B2(n_708),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4652),
.B(n_708),
.Y(n_4693)
);

AOI31xp33_ASAP7_75t_L g4694 ( 
.A1(n_4630),
.A2(n_717),
.A3(n_713),
.B(n_715),
.Y(n_4694)
);

AOI222xp33_ASAP7_75t_L g4695 ( 
.A1(n_4651),
.A2(n_4658),
.B1(n_4643),
.B2(n_4624),
.C1(n_4641),
.C2(n_4637),
.Y(n_4695)
);

OAI221xp5_ASAP7_75t_L g4696 ( 
.A1(n_4639),
.A2(n_719),
.B1(n_715),
.B2(n_717),
.C(n_721),
.Y(n_4696)
);

AOI221xp5_ASAP7_75t_L g4697 ( 
.A1(n_4640),
.A2(n_724),
.B1(n_719),
.B2(n_723),
.C(n_725),
.Y(n_4697)
);

AOI221xp5_ASAP7_75t_L g4698 ( 
.A1(n_4646),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.C(n_728),
.Y(n_4698)
);

INVxp33_ASAP7_75t_SL g4699 ( 
.A(n_4656),
.Y(n_4699)
);

INVx1_ASAP7_75t_SL g4700 ( 
.A(n_4670),
.Y(n_4700)
);

HB1xp67_ASAP7_75t_L g4701 ( 
.A(n_4667),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4676),
.Y(n_4702)
);

O2A1O1Ixp5_ASAP7_75t_SL g4703 ( 
.A1(n_4672),
.A2(n_728),
.B(n_726),
.C(n_727),
.Y(n_4703)
);

AOI22xp33_ASAP7_75t_L g4704 ( 
.A1(n_4660),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_SL g4705 ( 
.A(n_4634),
.B(n_729),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4673),
.B(n_731),
.Y(n_4706)
);

AOI221xp5_ASAP7_75t_L g4707 ( 
.A1(n_4635),
.A2(n_4645),
.B1(n_4633),
.B2(n_4669),
.C(n_4644),
.Y(n_4707)
);

AOI21xp33_ASAP7_75t_L g4708 ( 
.A1(n_4664),
.A2(n_4678),
.B(n_4648),
.Y(n_4708)
);

AOI22xp33_ASAP7_75t_L g4709 ( 
.A1(n_4653),
.A2(n_4661),
.B1(n_4666),
.B2(n_4628),
.Y(n_4709)
);

OAI211xp5_ASAP7_75t_SL g4710 ( 
.A1(n_4668),
.A2(n_734),
.B(n_732),
.C(n_733),
.Y(n_4710)
);

AOI211xp5_ASAP7_75t_L g4711 ( 
.A1(n_4638),
.A2(n_736),
.B(n_733),
.C(n_735),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4632),
.Y(n_4712)
);

NAND2x1p5_ASAP7_75t_L g4713 ( 
.A(n_4663),
.B(n_737),
.Y(n_4713)
);

AOI221xp5_ASAP7_75t_L g4714 ( 
.A1(n_4642),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.C(n_740),
.Y(n_4714)
);

INVx1_ASAP7_75t_SL g4715 ( 
.A(n_4677),
.Y(n_4715)
);

AND3x4_ASAP7_75t_L g4716 ( 
.A(n_4686),
.B(n_4647),
.C(n_4636),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4686),
.Y(n_4717)
);

CKINVDCx20_ASAP7_75t_R g4718 ( 
.A(n_4683),
.Y(n_4718)
);

AOI22xp5_ASAP7_75t_L g4719 ( 
.A1(n_4700),
.A2(n_4680),
.B1(n_4671),
.B2(n_4675),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4701),
.Y(n_4720)
);

AO22x2_ASAP7_75t_L g4721 ( 
.A1(n_4689),
.A2(n_4665),
.B1(n_4650),
.B2(n_4659),
.Y(n_4721)
);

NAND2xp5_ASAP7_75t_L g4722 ( 
.A(n_4694),
.B(n_4679),
.Y(n_4722)
);

AOI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4695),
.A2(n_741),
.B1(n_739),
.B2(n_740),
.Y(n_4723)
);

AND2x2_ASAP7_75t_SL g4724 ( 
.A(n_4693),
.B(n_742),
.Y(n_4724)
);

OAI22xp5_ASAP7_75t_L g4725 ( 
.A1(n_4681),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_4725)
);

AND2x2_ASAP7_75t_L g4726 ( 
.A(n_4706),
.B(n_4682),
.Y(n_4726)
);

NOR2x1_ASAP7_75t_L g4727 ( 
.A(n_4696),
.B(n_743),
.Y(n_4727)
);

AO22x2_ASAP7_75t_L g4728 ( 
.A1(n_4712),
.A2(n_747),
.B1(n_745),
.B2(n_746),
.Y(n_4728)
);

NOR2x1_ASAP7_75t_L g4729 ( 
.A(n_4705),
.B(n_4710),
.Y(n_4729)
);

OAI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4692),
.A2(n_749),
.B1(n_747),
.B2(n_748),
.Y(n_4730)
);

NOR2x1_ASAP7_75t_L g4731 ( 
.A(n_4702),
.B(n_748),
.Y(n_4731)
);

OAI31xp33_ASAP7_75t_L g4732 ( 
.A1(n_4715),
.A2(n_4688),
.A3(n_4685),
.B(n_4713),
.Y(n_4732)
);

AOI22xp5_ASAP7_75t_L g4733 ( 
.A1(n_4687),
.A2(n_753),
.B1(n_749),
.B2(n_752),
.Y(n_4733)
);

AOI21xp5_ASAP7_75t_L g4734 ( 
.A1(n_4716),
.A2(n_4698),
.B(n_4707),
.Y(n_4734)
);

NOR2x1_ASAP7_75t_L g4735 ( 
.A(n_4718),
.B(n_4684),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4728),
.Y(n_4736)
);

NOR3xp33_ASAP7_75t_L g4737 ( 
.A(n_4720),
.B(n_4708),
.C(n_4697),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4717),
.B(n_4703),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4728),
.Y(n_4739)
);

NOR2x1_ASAP7_75t_L g4740 ( 
.A(n_4726),
.B(n_4725),
.Y(n_4740)
);

XOR2xp5_ASAP7_75t_L g4741 ( 
.A(n_4721),
.B(n_4690),
.Y(n_4741)
);

OR2x2_ASAP7_75t_L g4742 ( 
.A(n_4722),
.B(n_4704),
.Y(n_4742)
);

INVx3_ASAP7_75t_L g4743 ( 
.A(n_4724),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4731),
.Y(n_4744)
);

NOR2x1_ASAP7_75t_L g4745 ( 
.A(n_4729),
.B(n_4711),
.Y(n_4745)
);

OAI322xp33_ASAP7_75t_L g4746 ( 
.A1(n_4741),
.A2(n_4719),
.A3(n_4723),
.B1(n_4733),
.B2(n_4730),
.C1(n_4732),
.C2(n_4699),
.Y(n_4746)
);

OAI211xp5_ASAP7_75t_L g4747 ( 
.A1(n_4735),
.A2(n_4709),
.B(n_4714),
.C(n_4691),
.Y(n_4747)
);

AOI211xp5_ASAP7_75t_L g4748 ( 
.A1(n_4734),
.A2(n_4727),
.B(n_756),
.C(n_754),
.Y(n_4748)
);

AOI21xp5_ASAP7_75t_L g4749 ( 
.A1(n_4738),
.A2(n_755),
.B(n_757),
.Y(n_4749)
);

NOR3xp33_ASAP7_75t_L g4750 ( 
.A(n_4737),
.B(n_757),
.C(n_758),
.Y(n_4750)
);

AOI211xp5_ASAP7_75t_L g4751 ( 
.A1(n_4744),
.A2(n_760),
.B(n_758),
.C(n_759),
.Y(n_4751)
);

AOI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_4745),
.A2(n_759),
.B(n_760),
.Y(n_4752)
);

OAI22xp5_ASAP7_75t_L g4753 ( 
.A1(n_4740),
.A2(n_764),
.B1(n_761),
.B2(n_762),
.Y(n_4753)
);

AOI21xp5_ASAP7_75t_L g4754 ( 
.A1(n_4742),
.A2(n_761),
.B(n_762),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4753),
.Y(n_4755)
);

OA22x2_ASAP7_75t_L g4756 ( 
.A1(n_4747),
.A2(n_4739),
.B1(n_4736),
.B2(n_4743),
.Y(n_4756)
);

XNOR2x1_ASAP7_75t_L g4757 ( 
.A(n_4746),
.B(n_764),
.Y(n_4757)
);

XNOR2xp5_ASAP7_75t_L g4758 ( 
.A(n_4748),
.B(n_767),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4756),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4757),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4758),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4759),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4762),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4763),
.Y(n_4764)
);

AOI221xp5_ASAP7_75t_L g4765 ( 
.A1(n_4764),
.A2(n_4749),
.B1(n_4750),
.B2(n_4760),
.C(n_4761),
.Y(n_4765)
);

XNOR2xp5_ASAP7_75t_L g4766 ( 
.A(n_4765),
.B(n_4755),
.Y(n_4766)
);

OA21x2_ASAP7_75t_L g4767 ( 
.A1(n_4766),
.A2(n_4752),
.B(n_4754),
.Y(n_4767)
);

OAI22xp33_ASAP7_75t_L g4768 ( 
.A1(n_4767),
.A2(n_4751),
.B1(n_770),
.B2(n_768),
.Y(n_4768)
);

AOI22xp5_ASAP7_75t_SL g4769 ( 
.A1(n_4767),
.A2(n_771),
.B1(n_768),
.B2(n_769),
.Y(n_4769)
);

OAI211xp5_ASAP7_75t_L g4770 ( 
.A1(n_4769),
.A2(n_775),
.B(n_772),
.C(n_773),
.Y(n_4770)
);

AO221x2_ASAP7_75t_L g4771 ( 
.A1(n_4768),
.A2(n_778),
.B1(n_776),
.B2(n_777),
.C(n_779),
.Y(n_4771)
);

AOI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4771),
.A2(n_776),
.B(n_777),
.Y(n_4772)
);

AOI211xp5_ASAP7_75t_L g4773 ( 
.A1(n_4772),
.A2(n_4770),
.B(n_782),
.C(n_778),
.Y(n_4773)
);


endmodule