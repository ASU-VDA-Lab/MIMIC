module fake_jpeg_28540_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_20),
.B1(n_30),
.B2(n_21),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_7),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_52),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_67),
.B1(n_62),
.B2(n_40),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_24),
.B1(n_28),
.B2(n_35),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_56),
.B1(n_73),
.B2(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_18),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_29),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_43),
.B1(n_41),
.B2(n_17),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_43),
.B1(n_41),
.B2(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_22),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_22),
.CI(n_19),
.CON(n_91),
.SN(n_91)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_16),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_19),
.B(n_5),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_74),
.B(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_101),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_108),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_8),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_103),
.B1(n_112),
.B2(n_90),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_54),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_134),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_62),
.B(n_54),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_8),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_13),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_134),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_108),
.B(n_95),
.C(n_101),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_10),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_13),
.Y(n_156)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_144),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_84),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_155),
.B(n_128),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_161),
.C(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_83),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_163),
.B1(n_127),
.B2(n_120),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_86),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_124),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_154),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_129),
.A3(n_122),
.B1(n_116),
.B2(n_121),
.C1(n_128),
.C2(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_156),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_121),
.B1(n_123),
.B2(n_114),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_179),
.B1(n_161),
.B2(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_121),
.B1(n_123),
.B2(n_114),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_126),
.B1(n_128),
.B2(n_119),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_144),
.B1(n_142),
.B2(n_126),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_184),
.B(n_133),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_132),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_133),
.B(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_168),
.B1(n_172),
.B2(n_170),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_146),
.B1(n_150),
.B2(n_126),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_193),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_167),
.A3(n_181),
.B1(n_165),
.B2(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_150),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_198),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_159),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_197),
.C(n_200),
.Y(n_212)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_182),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_147),
.Y(n_197)
);

AO32x1_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_160),
.A3(n_137),
.B1(n_151),
.B2(n_153),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_198),
.A2(n_180),
.B1(n_168),
.B2(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_175),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_188),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_170),
.B1(n_145),
.B2(n_141),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_85),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_199),
.B(n_192),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_218),
.Y(n_228)
);

AOI31xp67_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_201),
.A3(n_197),
.B(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_209),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_188),
.C(n_163),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_222),
.C(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_189),
.C(n_94),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_223),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_196),
.C(n_127),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_208),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_204),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_220),
.A2(n_213),
.B1(n_209),
.B2(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_230),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_217),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

FAx1_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_205),
.CI(n_222),
.CON(n_235),
.SN(n_235)
);

AOI221xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_229),
.B1(n_225),
.B2(n_223),
.C(n_221),
.Y(n_237)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_10),
.B(n_100),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_214),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_236),
.A2(n_110),
.B(n_106),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_231),
.B1(n_202),
.B2(n_139),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_232),
.C(n_111),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_232),
.B(n_100),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_243),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_88),
.C(n_87),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_97),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_244),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_97),
.Y(n_248)
);


endmodule