module fake_netlist_5_1941_n_1946 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1946);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1946;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_SL g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_94),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_45),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_53),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_72),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_36),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_84),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_33),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_49),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_36),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_51),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_10),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_47),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_163),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_144),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_119),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_50),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_130),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_45),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_175),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_3),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_87),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_97),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_26),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_124),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_61),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_85),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_81),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_7),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_65),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_71),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_61),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_111),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_96),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_89),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_131),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_13),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_90),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_107),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_160),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_70),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_44),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_122),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_2),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_56),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_169),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_93),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_128),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_109),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_114),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_152),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_127),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_59),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_49),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_186),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_171),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_18),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_53),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_75),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_34),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_118),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_38),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_146),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_196),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_149),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_26),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_194),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_69),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_40),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_138),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_176),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_37),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_191),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_126),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_162),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_154),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_157),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_56),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_41),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_142),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_57),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_29),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_28),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_7),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_113),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_151),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_166),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_92),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_110),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_148),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_28),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_57),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_63),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_143),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_174),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_43),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_129),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_82),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_33),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_22),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_62),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_203),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_31),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_91),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_134),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_15),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_135),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_20),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_165),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_98),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_20),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_100),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_77),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_116),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_112),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_3),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_185),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_64),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_139),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_108),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_106),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_54),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_34),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_78),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_18),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_104),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_64),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_48),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_133),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_145),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_17),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_73),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_51),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_102),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_120),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_5),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_132),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_167),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_179),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_4),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_19),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_137),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_170),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_12),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_32),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_159),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_153),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_201),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_178),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_63),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_83),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_54),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_190),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_47),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_168),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_22),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_30),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_86),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_52),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_136),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_88),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_30),
.Y(n_399)
);

CKINVDCx12_ASAP7_75t_R g400 ( 
.A(n_16),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_23),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_74),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_2),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_12),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_65),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_79),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_40),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_23),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_316),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_240),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_236),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_271),
.B(n_1),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_275),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_246),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_316),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_249),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_251),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_243),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_266),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_209),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_243),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_268),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_304),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_204),
.B(n_1),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_269),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_263),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_217),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_217),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_217),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_217),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_270),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_217),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_360),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_248),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_263),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_234),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_333),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_379),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_234),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_333),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_204),
.B(n_4),
.Y(n_448)
);

BUFx6f_ASAP7_75t_SL g449 ( 
.A(n_362),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_209),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_291),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_214),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_248),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_263),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_248),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_395),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_6),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_248),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_248),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_292),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_257),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_296),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_407),
.B(n_8),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_257),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_207),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_406),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_257),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_302),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_260),
.B(n_8),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_238),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_257),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_305),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_362),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_310),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_241),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_245),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_312),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_257),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_211),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_337),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_242),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_278),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_280),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_317),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_281),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_250),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_260),
.B(n_9),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_282),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_324),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_407),
.B(n_10),
.Y(n_493)
);

XOR2x2_ASAP7_75t_L g494 ( 
.A(n_219),
.B(n_11),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_286),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_214),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_287),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_326),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_215),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_253),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_289),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_330),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_331),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_299),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_303),
.B(n_11),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_334),
.Y(n_506)
);

BUFx6f_ASAP7_75t_SL g507 ( 
.A(n_212),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_254),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_258),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_299),
.B(n_14),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_255),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_336),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_R g515 ( 
.A(n_410),
.B(n_205),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_410),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_SL g519 ( 
.A(n_463),
.B(n_215),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_472),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_477),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_427),
.B(n_206),
.Y(n_522)
);

INVxp33_ASAP7_75t_SL g523 ( 
.A(n_417),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_478),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_409),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_426),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_411),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_509),
.A2(n_346),
.B1(n_327),
.B2(n_315),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_444),
.B(n_206),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g533 ( 
.A(n_432),
.B(n_216),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_413),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_436),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_483),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_489),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_500),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_437),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_508),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_512),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_R g545 ( 
.A(n_417),
.B(n_256),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_447),
.B(n_208),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_419),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_452),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_419),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_475),
.B(n_205),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_416),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_423),
.B(n_208),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_441),
.B(n_273),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_494),
.A2(n_218),
.B1(n_220),
.B2(n_403),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_421),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_496),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_425),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_425),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_424),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_423),
.B(n_463),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_441),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_473),
.B(n_273),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_428),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_473),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_431),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_431),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_455),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_438),
.B(n_259),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_438),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_448),
.B(n_272),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_458),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_459),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_469),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_481),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_451),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_504),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_511),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_486),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_488),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_451),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_460),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_460),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_462),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_517),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_522),
.B(n_293),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_551),
.B(n_462),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_564),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_591),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_555),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_564),
.B(n_443),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_553),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_470),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_522),
.B(n_293),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_514),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_522),
.B(n_430),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_523),
.B(n_470),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_526),
.B(n_450),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_553),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_577),
.B(n_474),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_530),
.A2(n_490),
.B1(n_415),
.B2(n_471),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_517),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_566),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_530),
.B(n_474),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_530),
.B(n_476),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_518),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_555),
.B(n_546),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_518),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_566),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_515),
.A2(n_480),
.B1(n_487),
.B2(n_476),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_566),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_546),
.B(n_318),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_553),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_555),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_518),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_546),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_545),
.B(n_318),
.Y(n_634)
);

BUFx6f_ASAP7_75t_SL g635 ( 
.A(n_556),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_539),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_525),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_556),
.B(n_376),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_553),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_525),
.Y(n_640)
);

CKINVDCx14_ASAP7_75t_R g641 ( 
.A(n_562),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_575),
.B(n_376),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_562),
.B(n_505),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_574),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_534),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_R g646 ( 
.A(n_520),
.B(n_429),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_576),
.B(n_594),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_539),
.B(n_534),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_539),
.B(n_480),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_527),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_577),
.B(n_487),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_539),
.B(n_534),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_547),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_587),
.B(n_446),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_552),
.B(n_440),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_553),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_519),
.B(n_498),
.C(n_492),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_556),
.A2(n_505),
.B1(n_493),
.B2(n_401),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_533),
.B(n_492),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_574),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_556),
.A2(n_567),
.B1(n_536),
.B2(n_563),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_584),
.Y(n_663)
);

CKINVDCx16_ASAP7_75t_R g664 ( 
.A(n_529),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_450),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_536),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_567),
.A2(n_422),
.B1(n_510),
.B2(n_335),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_533),
.B(n_498),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_569),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_536),
.B(n_502),
.Y(n_671)
);

BUFx8_ASAP7_75t_SL g672 ( 
.A(n_521),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_563),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_563),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_567),
.B(n_502),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_584),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_553),
.Y(n_677)
);

BUFx4f_ASAP7_75t_L g678 ( 
.A(n_558),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_558),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_558),
.B(n_503),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_558),
.B(n_337),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_526),
.B(n_454),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_558),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_588),
.B(n_491),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_567),
.A2(n_343),
.B1(n_405),
.B2(n_352),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_581),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_529),
.B(n_468),
.C(n_465),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_572),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_581),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_590),
.A2(n_341),
.B1(n_394),
.B2(n_359),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g692 ( 
.A(n_549),
.B(n_218),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_550),
.B(n_503),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_569),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_576),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_516),
.B(n_506),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_590),
.B(n_592),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_588),
.B(n_501),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_596),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_572),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_590),
.A2(n_314),
.B1(n_393),
.B2(n_370),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_516),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_549),
.B(n_479),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_579),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_559),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_581),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_528),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_579),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_580),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_580),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_528),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_560),
.B(n_506),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_531),
.B(n_513),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_561),
.B(n_513),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_582),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_595),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_531),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_592),
.B(n_227),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_532),
.B(n_294),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_532),
.B(n_261),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_559),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_535),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_581),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_568),
.B(n_228),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_592),
.A2(n_399),
.B1(n_378),
.B2(n_457),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_571),
.B(n_433),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_593),
.A2(n_507),
.B1(n_497),
.B2(n_485),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_582),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_535),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_594),
.A2(n_442),
.B1(n_347),
.B2(n_373),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_573),
.B(n_230),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_569),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_586),
.B(n_449),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_537),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_581),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_524),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_583),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_537),
.B(n_262),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_538),
.B(n_265),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_538),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_542),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_569),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_593),
.B(n_449),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_540),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_449),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_542),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_601),
.A2(n_445),
.B1(n_456),
.B2(n_467),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_597),
.B(n_222),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_633),
.B(n_548),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_633),
.B(n_548),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_618),
.B(n_557),
.C(n_414),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_636),
.B(n_554),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_624),
.A2(n_494),
.B1(n_557),
.B2(n_396),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_636),
.B(n_624),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_631),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_631),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_604),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_604),
.B(n_235),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_636),
.B(n_554),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_624),
.B(n_604),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_607),
.B(n_565),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_602),
.B(n_337),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_599),
.A2(n_337),
.B1(n_397),
.B2(n_348),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_702),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_621),
.A2(n_353),
.B1(n_329),
.B2(n_325),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_598),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_610),
.B(n_570),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_694),
.B(n_626),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_717),
.B(n_570),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_717),
.B(n_239),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_685),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_R g774 ( 
.A(n_641),
.B(n_541),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_680),
.B(n_244),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_648),
.A2(n_589),
.B(n_585),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_649),
.B(n_247),
.Y(n_777)
);

AO22x1_ASAP7_75t_L g778 ( 
.A1(n_616),
.A2(n_391),
.B1(n_237),
.B2(n_382),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_685),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_605),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_707),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_707),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_748),
.B(n_622),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_651),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_662),
.B(n_337),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_665),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_627),
.B(n_354),
.C(n_338),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_737),
.B(n_252),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_543),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_670),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_698),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_603),
.B(n_264),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_612),
.B(n_267),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_671),
.B(n_337),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_670),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_697),
.B(n_337),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_619),
.B(n_466),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_605),
.B(n_654),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_697),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_599),
.A2(n_337),
.B1(n_397),
.B2(n_385),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_697),
.B(n_397),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_696),
.B(n_713),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_617),
.B(n_277),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_652),
.A2(n_589),
.B(n_585),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_638),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_620),
.B(n_279),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_628),
.B(n_283),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_689),
.B(n_284),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_700),
.B(n_285),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_670),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_732),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_704),
.B(n_295),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_675),
.B(n_495),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_665),
.B(n_361),
.C(n_358),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_654),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_703),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_656),
.A2(n_589),
.B(n_585),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_615),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_638),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_726),
.B(n_544),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_708),
.B(n_298),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_672),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_709),
.B(n_308),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_710),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_675),
.B(n_724),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_715),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_728),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_608),
.A2(n_344),
.B(n_322),
.C(n_342),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_734),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_739),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_705),
.B(n_721),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_724),
.B(n_210),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_635),
.A2(n_658),
.B1(n_668),
.B2(n_660),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_744),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_711),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_629),
.B(n_744),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_718),
.B(n_629),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_635),
.A2(n_668),
.B1(n_660),
.B2(n_731),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_744),
.B(n_319),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_638),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_600),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_711),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_600),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_643),
.A2(n_366),
.B1(n_367),
.B2(n_356),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_720),
.B(n_740),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_731),
.B(n_210),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_741),
.B(n_351),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_672),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_722),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_722),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_SL g852 ( 
.A(n_695),
.B(n_213),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_609),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_609),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_729),
.B(n_380),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_614),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_705),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_638),
.A2(n_397),
.B1(n_402),
.B2(n_403),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_646),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_735),
.B(n_742),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_742),
.B(n_274),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_643),
.B(n_213),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_L g863 ( 
.A(n_712),
.B(n_714),
.C(n_693),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_743),
.B(n_276),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_719),
.B(n_634),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_721),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_634),
.B(n_288),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_643),
.B(n_221),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_642),
.B(n_397),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_643),
.B(n_363),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_642),
.B(n_221),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_659),
.A2(n_226),
.B1(n_225),
.B2(n_398),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_614),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_611),
.B(n_223),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_653),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_677),
.B(n_290),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_684),
.B(n_297),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_718),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_681),
.B(n_300),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_681),
.B(n_301),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_637),
.B(n_307),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_635),
.A2(n_350),
.B1(n_309),
.B2(n_311),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_640),
.B(n_313),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_613),
.B(n_220),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_638),
.B(n_320),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_645),
.B(n_321),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_644),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_678),
.A2(n_339),
.B(n_340),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_641),
.B(n_364),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_666),
.B(n_323),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_682),
.A2(n_507),
.B(n_369),
.C(n_328),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_673),
.B(n_332),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_674),
.B(n_345),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_615),
.B(n_630),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_647),
.B(n_365),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_733),
.B(n_349),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_615),
.B(n_355),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_712),
.B(n_223),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_678),
.A2(n_357),
.B(n_371),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_615),
.B(n_372),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_615),
.B(n_225),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_630),
.B(n_226),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_630),
.B(n_229),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_644),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_683),
.B(n_224),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_657),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_667),
.B(n_368),
.C(n_408),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_623),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_639),
.B(n_229),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_657),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_802),
.B(n_638),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_750),
.B(n_714),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_797),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_802),
.B(n_747),
.Y(n_914)
);

OAI321xp33_ASAP7_75t_L g915 ( 
.A1(n_750),
.A2(n_730),
.A3(n_683),
.B1(n_647),
.B2(n_727),
.C(n_725),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_825),
.A2(n_832),
.B(n_847),
.C(n_813),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_768),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_799),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_825),
.A2(n_745),
.B(n_692),
.C(n_686),
.Y(n_919)
);

OAI321xp33_ASAP7_75t_L g920 ( 
.A1(n_832),
.A2(n_847),
.A3(n_874),
.B1(n_898),
.B2(n_753),
.C(n_767),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_875),
.B(n_746),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_831),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_756),
.A2(n_647),
.B1(n_678),
.B2(n_691),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_763),
.B(n_623),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_874),
.A2(n_647),
.B(n_231),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_754),
.A2(n_639),
.B(n_736),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_761),
.A2(n_639),
.B(n_736),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_764),
.A2(n_625),
.B(n_632),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_799),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_786),
.B(n_653),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_784),
.B(n_816),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_894),
.A2(n_762),
.B(n_836),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_859),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_762),
.A2(n_846),
.B(n_837),
.Y(n_934)
);

O2A1O1Ixp5_ASAP7_75t_L g935 ( 
.A1(n_794),
.A2(n_669),
.B(n_676),
.C(n_663),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_857),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_878),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_837),
.A2(n_818),
.B(n_770),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_805),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_865),
.B(n_625),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_783),
.B(n_632),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_759),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_769),
.B(n_661),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_SL g944 ( 
.A(n_805),
.B(n_232),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_794),
.A2(n_676),
.B(n_669),
.C(n_661),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_758),
.B(n_653),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_805),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_764),
.A2(n_663),
.B(n_736),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_780),
.B(n_699),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_780),
.B(n_699),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_766),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_776),
.A2(n_682),
.B(n_690),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_804),
.A2(n_690),
.B(n_701),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_818),
.A2(n_690),
.B(n_606),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_840),
.B(n_813),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_820),
.B(n_650),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_757),
.B(n_751),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_758),
.B(n_699),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_860),
.A2(n_738),
.B(n_706),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_752),
.B(n_706),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_879),
.A2(n_606),
.B(n_679),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_880),
.A2(n_606),
.B(n_679),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_758),
.B(n_706),
.Y(n_963)
);

O2A1O1Ixp5_ASAP7_75t_L g964 ( 
.A1(n_785),
.A2(n_692),
.B(n_507),
.C(n_723),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_758),
.B(n_706),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_759),
.B(n_716),
.Y(n_966)
);

AOI33xp33_ASAP7_75t_L g967 ( 
.A1(n_755),
.A2(n_664),
.A3(n_688),
.B1(n_237),
.B2(n_377),
.B3(n_382),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_876),
.A2(n_679),
.B(n_606),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_877),
.A2(n_679),
.B(n_606),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_863),
.B(n_388),
.C(n_233),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_805),
.B(n_738),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_785),
.A2(n_679),
.B(n_306),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_775),
.A2(n_771),
.B(n_777),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_819),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_781),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_781),
.A2(n_388),
.B(n_374),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_811),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_798),
.B(n_716),
.Y(n_978)
);

NOR2x1_ASAP7_75t_L g979 ( 
.A(n_814),
.B(n_655),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_798),
.B(n_716),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_885),
.A2(n_738),
.B(n_723),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_782),
.A2(n_386),
.B(n_374),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_866),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_788),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_819),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_838),
.A2(n_375),
.B1(n_384),
.B2(n_398),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_899),
.A2(n_723),
.B(n_687),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_828),
.A2(n_386),
.B(n_390),
.C(n_375),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_833),
.B(n_723),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_778),
.B(n_392),
.C(n_390),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_773),
.B(n_687),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_782),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_902),
.A2(n_687),
.B(n_392),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_779),
.B(n_687),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_903),
.A2(n_909),
.B(n_811),
.Y(n_995)
);

OAI21xp33_ASAP7_75t_L g996 ( 
.A1(n_755),
.A2(n_224),
.B(n_391),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_817),
.A2(n_687),
.B(n_384),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_819),
.B(n_383),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_897),
.A2(n_383),
.B(n_387),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_897),
.A2(n_900),
.B(n_795),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_900),
.A2(n_389),
.B(n_387),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_774),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_790),
.A2(n_389),
.B(n_377),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_810),
.A2(n_231),
.B(n_95),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_834),
.A2(n_202),
.B(n_200),
.Y(n_1005)
);

AO21x1_ASAP7_75t_L g1006 ( 
.A1(n_871),
.A2(n_869),
.B(n_901),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_861),
.A2(n_199),
.B(n_198),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_791),
.A2(n_193),
.B1(n_188),
.B2(n_183),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_871),
.A2(n_16),
.B(n_17),
.C(n_21),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_789),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_815),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_858),
.A2(n_181),
.B1(n_180),
.B2(n_173),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_760),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_905),
.B(n_24),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_824),
.B(n_25),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_826),
.B(n_827),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_864),
.A2(n_172),
.B(n_158),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_829),
.B(n_27),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_L g1019 ( 
.A(n_788),
.Y(n_1019)
);

NAND3xp33_ASAP7_75t_L g1020 ( 
.A(n_852),
.B(n_29),
.C(n_31),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_848),
.A2(n_32),
.B(n_35),
.C(n_37),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_830),
.B(n_35),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_835),
.B(n_39),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_883),
.A2(n_123),
.B(n_121),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_843),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_892),
.A2(n_117),
.B(n_115),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_850),
.B(n_41),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_851),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_893),
.A2(n_105),
.B(n_103),
.Y(n_1029)
);

NOR2x1p5_ASAP7_75t_L g1030 ( 
.A(n_822),
.B(n_42),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_819),
.B(n_99),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_870),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_772),
.B(n_46),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_787),
.B(n_50),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_792),
.B(n_52),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_867),
.B(n_55),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_881),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_908),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_841),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_896),
.B(n_58),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_884),
.B(n_66),
.C(n_67),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_828),
.A2(n_901),
.B(n_869),
.C(n_801),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_887),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_796),
.A2(n_801),
.B(n_839),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_862),
.A2(n_868),
.B(n_891),
.C(n_806),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_793),
.B(n_821),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_841),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_841),
.A2(n_749),
.B1(n_765),
.B2(n_800),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_808),
.B(n_823),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_904),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_842),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_841),
.A2(n_906),
.B(n_910),
.Y(n_1053)
);

OAI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_868),
.A2(n_872),
.B(n_907),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_809),
.B(n_812),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_881),
.A2(n_890),
.B(n_886),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_803),
.A2(n_807),
.B(n_855),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_886),
.A2(n_890),
.B(n_853),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_895),
.B(n_889),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_L g1060 ( 
.A1(n_844),
.A2(n_873),
.B(n_856),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_854),
.B(n_765),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_788),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_888),
.A2(n_800),
.B(n_845),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_882),
.A2(n_774),
.B(n_822),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_849),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_849),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_802),
.B(n_763),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_799),
.Y(n_1068)
);

NAND3xp33_ASAP7_75t_L g1069 ( 
.A(n_750),
.B(n_874),
.C(n_597),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_750),
.B(n_784),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_758),
.B(n_846),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_799),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_750),
.B(n_874),
.C(n_597),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_759),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_802),
.B(n_763),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_750),
.B(n_784),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_764),
.A2(n_761),
.B(n_754),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_750),
.B(n_784),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_797),
.B(n_831),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_L g1080 ( 
.A(n_768),
.B(n_746),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_758),
.B(n_802),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_750),
.B(n_784),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_756),
.A2(n_636),
.B(n_678),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_934),
.A2(n_911),
.B(n_1071),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1060),
.A2(n_981),
.B(n_945),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_935),
.A2(n_945),
.B(n_932),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_989),
.A2(n_935),
.B(n_1006),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_985),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1079),
.B(n_1070),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_951),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_912),
.A2(n_920),
.B1(n_1073),
.B2(n_1069),
.C(n_1082),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_L g1093 ( 
.A(n_970),
.B(n_1002),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_985),
.Y(n_1094)
);

OAI21xp33_ASAP7_75t_SL g1095 ( 
.A1(n_912),
.A2(n_1081),
.B(n_914),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_916),
.A2(n_1076),
.B1(n_1082),
.B2(n_1078),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_947),
.B(n_1031),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_921),
.B(n_1080),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1070),
.B(n_1076),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_917),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_939),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1078),
.A2(n_1055),
.B1(n_1050),
.B2(n_1047),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_995),
.A2(n_1083),
.B(n_1077),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1013),
.B(n_1032),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1071),
.A2(n_938),
.B(n_1045),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_943),
.B(n_941),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_973),
.A2(n_952),
.B(n_1063),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_989),
.A2(n_987),
.B(n_1000),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_917),
.B(n_1059),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_953),
.A2(n_960),
.B(n_940),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1053),
.A2(n_927),
.B(n_926),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_1059),
.B(n_1065),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1043),
.A2(n_924),
.B(n_1056),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_955),
.B(n_957),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1061),
.A2(n_964),
.B(n_1046),
.Y(n_1115)
);

AOI21x1_ASAP7_75t_L g1116 ( 
.A1(n_997),
.A2(n_1058),
.B(n_963),
.Y(n_1116)
);

AOI221xp5_ASAP7_75t_L g1117 ( 
.A1(n_1034),
.A2(n_1014),
.B1(n_915),
.B2(n_1009),
.C(n_1054),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_1034),
.A2(n_1014),
.B(n_955),
.Y(n_1118)
);

OA22x2_ASAP7_75t_L g1119 ( 
.A1(n_996),
.A2(n_913),
.B1(n_925),
.B2(n_986),
.Y(n_1119)
);

O2A1O1Ixp5_ASAP7_75t_L g1120 ( 
.A1(n_964),
.A2(n_998),
.B(n_944),
.C(n_993),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_931),
.B(n_1010),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_975),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_965),
.A2(n_947),
.B(n_1049),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_922),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_992),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_947),
.A2(n_998),
.B(n_994),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_949),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1066),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_961),
.A2(n_962),
.B(n_954),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_977),
.B(n_919),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_977),
.B(n_931),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_968),
.A2(n_969),
.B(n_971),
.Y(n_1132)
);

AO21x1_ASAP7_75t_L g1133 ( 
.A1(n_1012),
.A2(n_1033),
.B(n_1041),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1016),
.B(n_937),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_990),
.A2(n_1037),
.B1(n_923),
.B2(n_1013),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_971),
.A2(n_1057),
.B(n_991),
.Y(n_1136)
);

INVx6_ASAP7_75t_L g1137 ( 
.A(n_950),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1025),
.B(n_1028),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_983),
.Y(n_1139)
);

INVx8_ASAP7_75t_L g1140 ( 
.A(n_947),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_972),
.A2(n_1031),
.B(n_1040),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_930),
.B(n_983),
.Y(n_1142)
);

AO21x1_ASAP7_75t_L g1143 ( 
.A1(n_1035),
.A2(n_1023),
.B(n_1027),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1036),
.A2(n_1044),
.B(n_1051),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1072),
.A2(n_1052),
.B(n_1040),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_939),
.A2(n_1048),
.B(n_974),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_918),
.A2(n_929),
.B(n_1068),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_942),
.Y(n_1148)
);

AOI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_1015),
.A2(n_1022),
.B(n_1018),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_942),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_966),
.B(n_936),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1005),
.A2(n_1024),
.B(n_1029),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_958),
.A2(n_982),
.B(n_976),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1021),
.A2(n_1011),
.A3(n_1026),
.B(n_1017),
.Y(n_1154)
);

INVx11_ASAP7_75t_L g1155 ( 
.A(n_984),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1074),
.B(n_939),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1074),
.B(n_939),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1007),
.A2(n_1004),
.B(n_958),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_974),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_L g1160 ( 
.A1(n_946),
.A2(n_999),
.B(n_980),
.C(n_978),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_966),
.B(n_1019),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1062),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_974),
.B(n_1048),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1003),
.A2(n_1001),
.B(n_956),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_974),
.Y(n_1165)
);

INVx8_ASAP7_75t_L g1166 ( 
.A(n_1048),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1019),
.B(n_1062),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1064),
.A2(n_988),
.A3(n_1038),
.B(n_1042),
.Y(n_1168)
);

AOI21x1_ASAP7_75t_SL g1169 ( 
.A1(n_990),
.A2(n_1008),
.B(n_967),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1048),
.A2(n_979),
.B(n_1020),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1030),
.A2(n_928),
.B(n_948),
.Y(n_1171)
);

AOI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_933),
.A2(n_912),
.B(n_1069),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_959),
.A2(n_1071),
.B(n_989),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1065),
.B(n_1066),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_917),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_917),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1067),
.A2(n_1075),
.B1(n_1069),
.B2(n_1073),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1013),
.B(n_759),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1067),
.A2(n_1075),
.B(n_912),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1039),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_SL g1185 ( 
.A1(n_916),
.A2(n_911),
.B(n_1031),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_SL g1186 ( 
.A1(n_934),
.A2(n_1006),
.B(n_1056),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_939),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_928),
.A2(n_948),
.B(n_959),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_934),
.A2(n_911),
.B(n_1071),
.Y(n_1191)
);

CKINVDCx14_ASAP7_75t_R g1192 ( 
.A(n_1002),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_939),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1006),
.A2(n_916),
.A3(n_1046),
.B(n_987),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_947),
.B(n_985),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_917),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1067),
.A2(n_1075),
.B1(n_1069),
.B2(n_1073),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_928),
.A2(n_948),
.B(n_959),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_912),
.A2(n_916),
.B(n_1073),
.C(n_1069),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1013),
.B(n_759),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1069),
.B(n_1073),
.C(n_912),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1069),
.B(n_1073),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1208)
);

OAI22x1_ASAP7_75t_L g1209 ( 
.A1(n_912),
.A2(n_1073),
.B1(n_1069),
.B2(n_1070),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_928),
.A2(n_948),
.B(n_959),
.Y(n_1210)
);

O2A1O1Ixp5_ASAP7_75t_L g1211 ( 
.A1(n_1069),
.A2(n_1073),
.B(n_912),
.C(n_916),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_939),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_934),
.A2(n_636),
.B(n_756),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1006),
.A2(n_916),
.A3(n_1046),
.B(n_987),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_934),
.A2(n_911),
.B(n_1071),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_912),
.A2(n_750),
.B(n_1070),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1107),
.A2(n_1113),
.B(n_1110),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1216),
.B(n_1099),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1188),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1121),
.B(n_1109),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_R g1223 ( 
.A(n_1192),
.B(n_1098),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1211),
.A2(n_1118),
.B(n_1092),
.C(n_1117),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1090),
.B(n_1142),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1140),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1092),
.A2(n_1118),
.B1(n_1205),
.B2(n_1117),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1155),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1107),
.A2(n_1113),
.B(n_1110),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1179),
.B(n_1180),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1127),
.B(n_1099),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1176),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1091),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1177),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1198),
.Y(n_1235)
);

OAI21xp33_ASAP7_75t_L g1236 ( 
.A1(n_1180),
.A2(n_1187),
.B(n_1183),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1124),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1139),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1209),
.B(n_1151),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1188),
.Y(n_1240)
);

INVx8_ASAP7_75t_L g1241 ( 
.A(n_1166),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1100),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1104),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1181),
.B(n_1204),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1104),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1122),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1114),
.B(n_1181),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1125),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1183),
.B(n_1187),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1140),
.Y(n_1250)
);

OAI31xp33_ASAP7_75t_L g1251 ( 
.A1(n_1096),
.A2(n_1201),
.A3(n_1178),
.B(n_1102),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1128),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_1170),
.B(n_1162),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1175),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1175),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1114),
.B(n_1190),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1213),
.A2(n_1185),
.B(n_1105),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1204),
.B(n_1167),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1190),
.B(n_1193),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1140),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1087),
.A2(n_1191),
.B(n_1084),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1131),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1175),
.Y(n_1263)
);

AND2x6_ASAP7_75t_L g1264 ( 
.A(n_1089),
.B(n_1094),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1137),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1144),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1112),
.B(n_1161),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1166),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1206),
.A2(n_1172),
.B1(n_1093),
.B2(n_1207),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1166),
.B(n_1097),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1193),
.B(n_1196),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1089),
.B(n_1094),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1148),
.B(n_1134),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1137),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1199),
.B(n_1200),
.Y(n_1275)
);

INVx3_ASAP7_75t_SL g1276 ( 
.A(n_1137),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1131),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1186),
.A2(n_1215),
.B(n_1153),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1106),
.A2(n_1141),
.B(n_1199),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1188),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1200),
.A2(n_1207),
.B1(n_1208),
.B2(n_1134),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1208),
.B(n_1182),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1159),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1194),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_1097),
.B1(n_1135),
.B2(n_1130),
.Y(n_1285)
);

BUFx4_ASAP7_75t_SL g1286 ( 
.A(n_1150),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1172),
.B(n_1095),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1184),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1130),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1163),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1101),
.B(n_1165),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_1194),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1164),
.B(n_1212),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1119),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1149),
.B(n_1156),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1194),
.B(n_1212),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1157),
.B(n_1163),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1168),
.B(n_1157),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1212),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1168),
.B(n_1214),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1123),
.A2(n_1108),
.B(n_1120),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1197),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1143),
.B(n_1133),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1197),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1171),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1147),
.B(n_1168),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1111),
.A2(n_1126),
.B(n_1103),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1145),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1154),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1146),
.B(n_1154),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1129),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1195),
.B(n_1214),
.Y(n_1312)
);

NAND2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1136),
.B(n_1088),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1174),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_SL g1315 ( 
.A(n_1116),
.B(n_1160),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1088),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1169),
.A2(n_1132),
.B1(n_1085),
.B2(n_1189),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1195),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1214),
.A2(n_1154),
.B1(n_1202),
.B2(n_1210),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1086),
.A2(n_1067),
.B1(n_1075),
.B2(n_1173),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1216),
.A2(n_912),
.B1(n_1073),
.B2(n_1069),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1140),
.B(n_1166),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1089),
.B(n_1094),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1326)
);

NAND2x1_ASAP7_75t_L g1327 ( 
.A(n_1089),
.B(n_1094),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1176),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1216),
.B(n_1069),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1124),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1138),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1176),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1333)
);

NOR2xp67_ASAP7_75t_L g1334 ( 
.A(n_1100),
.B(n_768),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_1100),
.B(n_768),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1138),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1090),
.B(n_1079),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1181),
.B(n_1204),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1176),
.Y(n_1339)
);

AOI21xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1121),
.A2(n_912),
.B(n_750),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1140),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1216),
.A2(n_912),
.B1(n_1118),
.B2(n_1096),
.C(n_750),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1140),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1107),
.A2(n_1113),
.B(n_1110),
.Y(n_1345)
);

NOR3xp33_ASAP7_75t_L g1346 ( 
.A(n_1216),
.B(n_1073),
.C(n_1069),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1086),
.B(n_1173),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1181),
.B(n_1204),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1176),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1181),
.B(n_1204),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1086),
.A2(n_1067),
.B1(n_1075),
.B2(n_1173),
.Y(n_1351)
);

NOR2x1_ASAP7_75t_L g1352 ( 
.A(n_1121),
.B(n_737),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1203),
.A2(n_916),
.B(n_1118),
.C(n_1117),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1216),
.B(n_1069),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1216),
.B(n_1069),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1107),
.A2(n_1113),
.B(n_1110),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1176),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1099),
.B(n_650),
.Y(n_1358)
);

INVx3_ASAP7_75t_SL g1359 ( 
.A(n_1175),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1138),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1225),
.B(n_1337),
.Y(n_1361)
);

AO21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1303),
.A2(n_1282),
.B(n_1227),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1342),
.A2(n_1355),
.B1(n_1354),
.B2(n_1329),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1286),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1248),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1290),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1292),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1223),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1311),
.A2(n_1307),
.B(n_1301),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1228),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1292),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1342),
.A2(n_1346),
.B1(n_1251),
.B2(n_1322),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1246),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1330),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_SL g1375 ( 
.A1(n_1285),
.A2(n_1295),
.B(n_1282),
.Y(n_1375)
);

AO21x1_ASAP7_75t_L g1376 ( 
.A1(n_1251),
.A2(n_1287),
.B(n_1340),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1344),
.B(n_1292),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1358),
.B(n_1231),
.Y(n_1378)
);

INVx5_ASAP7_75t_L g1379 ( 
.A(n_1324),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1257),
.A2(n_1356),
.B(n_1217),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1242),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1247),
.B(n_1244),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1241),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1219),
.A2(n_1294),
.B1(n_1321),
.B2(n_1351),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1274),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1236),
.A2(n_1321),
.B1(n_1351),
.B2(n_1281),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1288),
.Y(n_1388)
);

BUFx2_ASAP7_75t_R g1389 ( 
.A(n_1237),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1352),
.A2(n_1267),
.B1(n_1269),
.B2(n_1222),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1273),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1279),
.A2(n_1224),
.B(n_1285),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1276),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1235),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1290),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_SL g1396 ( 
.A(n_1332),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1297),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1359),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1297),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1281),
.A2(n_1360),
.B1(n_1331),
.B2(n_1336),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1232),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1218),
.B(n_1220),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1241),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1328),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1298),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1217),
.A2(n_1356),
.B(n_1345),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1339),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1267),
.A2(n_1258),
.B1(n_1239),
.B2(n_1333),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1234),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1244),
.B(n_1338),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1229),
.A2(n_1303),
.B(n_1318),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1344),
.B(n_1226),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1349),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1277),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1218),
.A2(n_1220),
.B1(n_1347),
.B2(n_1230),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1273),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1241),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1238),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1357),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1324),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1234),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1324),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1221),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1262),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1313),
.A2(n_1266),
.B(n_1305),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1262),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1320),
.A2(n_1310),
.B(n_1295),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1317),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1283),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1256),
.Y(n_1431)
);

CKINVDCx6p67_ASAP7_75t_R g1432 ( 
.A(n_1252),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1230),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1249),
.A2(n_1343),
.B1(n_1347),
.B2(n_1326),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1313),
.A2(n_1305),
.B(n_1320),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1245),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1258),
.A2(n_1275),
.B1(n_1343),
.B2(n_1323),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1249),
.A2(n_1333),
.B1(n_1326),
.B2(n_1275),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1259),
.A2(n_1323),
.B1(n_1271),
.B2(n_1316),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1319),
.A2(n_1300),
.B(n_1312),
.Y(n_1440)
);

BUFx4f_ASAP7_75t_SL g1441 ( 
.A(n_1221),
.Y(n_1441)
);

INVx3_ASAP7_75t_SL g1442 ( 
.A(n_1296),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1259),
.A2(n_1271),
.B1(n_1289),
.B2(n_1306),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1264),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1243),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1254),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1253),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1255),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1334),
.A2(n_1335),
.B1(n_1263),
.B2(n_1291),
.Y(n_1449)
);

CKINVDCx6p67_ASAP7_75t_R g1450 ( 
.A(n_1268),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1240),
.Y(n_1451)
);

BUFx8_ASAP7_75t_SL g1452 ( 
.A(n_1280),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1306),
.A2(n_1309),
.B1(n_1353),
.B2(n_1310),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1291),
.B(n_1264),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1278),
.A2(n_1293),
.B1(n_1261),
.B2(n_1314),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1296),
.B(n_1299),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1272),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1270),
.B(n_1293),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1278),
.A2(n_1261),
.B1(n_1314),
.B2(n_1270),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1270),
.B(n_1268),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1314),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1250),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1315),
.A2(n_1325),
.B1(n_1304),
.B2(n_1302),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1327),
.B(n_1304),
.Y(n_1464)
);

INVxp67_ASAP7_75t_SL g1465 ( 
.A(n_1308),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1284),
.B(n_1260),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1260),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1341),
.A2(n_1301),
.B(n_1115),
.Y(n_1468)
);

INVx6_ASAP7_75t_L g1469 ( 
.A(n_1341),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1238),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1233),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1233),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1225),
.B(n_1337),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1344),
.B(n_1292),
.Y(n_1474)
);

INVx4_ASAP7_75t_SL g1475 ( 
.A(n_1264),
.Y(n_1475)
);

AO21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1303),
.A2(n_1282),
.B(n_1227),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1342),
.A2(n_1216),
.B1(n_912),
.B2(n_1118),
.Y(n_1477)
);

BUFx4f_ASAP7_75t_L g1478 ( 
.A(n_1241),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1292),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1301),
.A2(n_1115),
.B(n_1217),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_SL g1481 ( 
.A(n_1228),
.B(n_672),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1233),
.Y(n_1482)
);

INVx8_ASAP7_75t_L g1483 ( 
.A(n_1241),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1264),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1244),
.B(n_1338),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1218),
.A2(n_1069),
.B1(n_1073),
.B2(n_912),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1225),
.B(n_1337),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1366),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1440),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1440),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1429),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1392),
.B(n_1375),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1429),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1402),
.B(n_1433),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1405),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1362),
.B(n_1476),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1405),
.B(n_1376),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1428),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1366),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1443),
.B(n_1378),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1411),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1411),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1395),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1458),
.B(n_1465),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1435),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1426),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1406),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_SL g1510 ( 
.A(n_1389),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1373),
.Y(n_1511)
);

OAI222xp33_ASAP7_75t_L g1512 ( 
.A1(n_1363),
.A2(n_1372),
.B1(n_1477),
.B2(n_1385),
.C1(n_1439),
.C2(n_1486),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1369),
.A2(n_1380),
.B(n_1465),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1468),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1387),
.A2(n_1455),
.B(n_1453),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1443),
.B(n_1385),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1387),
.B(n_1480),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1415),
.B(n_1437),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1372),
.B(n_1439),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1453),
.B(n_1431),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1425),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1477),
.A2(n_1390),
.B(n_1447),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1388),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1455),
.A2(n_1459),
.B(n_1444),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1400),
.B(n_1415),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1400),
.B(n_1361),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1427),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1365),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1434),
.B(n_1438),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1471),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1458),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1472),
.Y(n_1532)
);

AOI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1461),
.A2(n_1454),
.B(n_1457),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1473),
.B(n_1487),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1458),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1482),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1379),
.B(n_1421),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1459),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1370),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_SL g1540 ( 
.A(n_1368),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1408),
.B(n_1430),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1417),
.B(n_1391),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1379),
.B(n_1421),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1409),
.B(n_1382),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1463),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1463),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1414),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1460),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1445),
.B(n_1456),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1470),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1460),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1470),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1393),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1467),
.A2(n_1449),
.B(n_1466),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1423),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1422),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_SL g1557 ( 
.A(n_1364),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1419),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1484),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1475),
.Y(n_1560)
);

CKINVDCx6p67_ASAP7_75t_R g1561 ( 
.A(n_1374),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1464),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1475),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1446),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1464),
.Y(n_1565)
);

AO21x1_ASAP7_75t_L g1566 ( 
.A1(n_1423),
.A2(n_1474),
.B(n_1377),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1404),
.B(n_1407),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1464),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1475),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1462),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1483),
.B(n_1412),
.Y(n_1571)
);

AO21x2_ASAP7_75t_L g1572 ( 
.A1(n_1410),
.A2(n_1416),
.B(n_1485),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1413),
.B(n_1420),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1377),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1367),
.Y(n_1575)
);

INVxp33_ASAP7_75t_L g1576 ( 
.A(n_1394),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1371),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1489),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1517),
.B(n_1448),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1517),
.B(n_1384),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1512),
.B(n_1384),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1495),
.B(n_1432),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1538),
.B(n_1442),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1490),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1519),
.A2(n_1436),
.B1(n_1420),
.B2(n_1413),
.Y(n_1585)
);

NOR4xp25_ASAP7_75t_SL g1586 ( 
.A(n_1553),
.B(n_1545),
.C(n_1546),
.D(n_1535),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1519),
.A2(n_1436),
.B1(n_1386),
.B2(n_1398),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1524),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1501),
.B(n_1424),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1491),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1529),
.B(n_1424),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1495),
.B(n_1381),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1516),
.A2(n_1386),
.B1(n_1398),
.B2(n_1401),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1493),
.B(n_1451),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1554),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1522),
.B(n_1393),
.C(n_1374),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1526),
.B(n_1469),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1500),
.B(n_1371),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1511),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1492),
.A2(n_1513),
.B(n_1509),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1524),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1497),
.B(n_1371),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1497),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1520),
.B(n_1418),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1508),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1562),
.B(n_1418),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1496),
.B(n_1396),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1502),
.B(n_1479),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1502),
.B(n_1498),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1492),
.B(n_1483),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1515),
.B(n_1479),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1515),
.B(n_1383),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1498),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1515),
.B(n_1523),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_SL g1616 ( 
.A(n_1561),
.B(n_1478),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1515),
.B(n_1383),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1488),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1492),
.B(n_1403),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1492),
.B(n_1403),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1528),
.B(n_1450),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1528),
.B(n_1481),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1541),
.B(n_1396),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1580),
.B(n_1525),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1580),
.B(n_1525),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1581),
.B(n_1541),
.C(n_1545),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1618),
.B(n_1521),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1625),
.B(n_1576),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1597),
.A2(n_1516),
.B1(n_1496),
.B2(n_1518),
.Y(n_1633)
);

OAI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1597),
.A2(n_1546),
.B1(n_1573),
.B2(n_1556),
.C(n_1494),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1581),
.A2(n_1562),
.B(n_1568),
.Y(n_1635)
);

OAI21xp33_ASAP7_75t_L g1636 ( 
.A1(n_1585),
.A2(n_1534),
.B(n_1544),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1572),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1572),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1618),
.B(n_1527),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1579),
.B(n_1622),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1625),
.B(n_1623),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1579),
.B(n_1547),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1601),
.B(n_1554),
.C(n_1565),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1622),
.B(n_1547),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1587),
.A2(n_1563),
.B(n_1560),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1599),
.B(n_1550),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1552),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1615),
.B(n_1513),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1601),
.A2(n_1503),
.B(n_1504),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1623),
.B(n_1574),
.C(n_1565),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1583),
.B(n_1554),
.C(n_1568),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1612),
.B(n_1513),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1590),
.A2(n_1596),
.B(n_1610),
.Y(n_1654)
);

NAND2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1586),
.B(n_1560),
.Y(n_1655)
);

NOR3xp33_ASAP7_75t_L g1656 ( 
.A(n_1592),
.B(n_1574),
.C(n_1569),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1514),
.Y(n_1657)
);

OAI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1616),
.A2(n_1531),
.B1(n_1561),
.B2(n_1571),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1613),
.B(n_1617),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1589),
.B(n_1558),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1594),
.A2(n_1564),
.B1(n_1567),
.B2(n_1569),
.C(n_1563),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1603),
.B(n_1532),
.Y(n_1662)
);

OAI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1594),
.A2(n_1531),
.B1(n_1551),
.B2(n_1548),
.C(n_1555),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1585),
.A2(n_1587),
.B1(n_1531),
.B2(n_1605),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1621),
.B(n_1566),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_SL g1666 ( 
.A(n_1624),
.B(n_1566),
.C(n_1510),
.D(n_1549),
.Y(n_1666)
);

OAI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1590),
.A2(n_1542),
.B(n_1533),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1611),
.B(n_1506),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1592),
.B(n_1532),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1608),
.A2(n_1537),
.B(n_1543),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1610),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1626),
.B(n_1514),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1616),
.A2(n_1551),
.B1(n_1548),
.B2(n_1555),
.C(n_1571),
.Y(n_1673)
);

XOR2xp5_ASAP7_75t_L g1674 ( 
.A(n_1598),
.B(n_1539),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1582),
.A2(n_1557),
.B1(n_1548),
.B2(n_1551),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1600),
.B(n_1577),
.C(n_1575),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1626),
.B(n_1507),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1619),
.A2(n_1537),
.B(n_1543),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1609),
.B(n_1536),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1596),
.B(n_1506),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1588),
.B(n_1570),
.C(n_1559),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1671),
.B(n_1614),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1677),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1677),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1630),
.B(n_1607),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1640),
.B(n_1578),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1658),
.B(n_1607),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1679),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1632),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1646),
.B(n_1649),
.Y(n_1690)
);

INVx3_ASAP7_75t_SL g1691 ( 
.A(n_1665),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1659),
.B(n_1588),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1680),
.B(n_1578),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1672),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1646),
.B(n_1588),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1588),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1653),
.B(n_1657),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1650),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1672),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1649),
.B(n_1637),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1578),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1644),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1680),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1642),
.Y(n_1704)
);

NAND2x1_ASAP7_75t_L g1705 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1669),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1673),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1666),
.A2(n_1611),
.B1(n_1619),
.B2(n_1620),
.Y(n_1708)
);

AND2x4_ASAP7_75t_SL g1709 ( 
.A(n_1668),
.B(n_1611),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1650),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1662),
.B(n_1614),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1631),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1639),
.B(n_1584),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1667),
.B(n_1591),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1665),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1682),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1682),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1717),
.B(n_1656),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1700),
.B(n_1652),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1634),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1683),
.Y(n_1723)
);

INVxp67_ASAP7_75t_SL g1724 ( 
.A(n_1698),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1683),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1697),
.B(n_1641),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1717),
.B(n_1647),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1698),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1709),
.B(n_1643),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1695),
.B(n_1651),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1684),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1684),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1695),
.B(n_1635),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1697),
.B(n_1678),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1702),
.B(n_1648),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1697),
.B(n_1611),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1713),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1710),
.Y(n_1739)
);

INVxp33_ASAP7_75t_L g1740 ( 
.A(n_1714),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1705),
.B(n_1685),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1702),
.B(n_1591),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1690),
.B(n_1593),
.Y(n_1745)
);

AOI33xp33_ASAP7_75t_L g1746 ( 
.A1(n_1712),
.A2(n_1633),
.A3(n_1664),
.B1(n_1586),
.B2(n_1549),
.B3(n_1624),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1710),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1681),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1692),
.B(n_1696),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1705),
.B(n_1606),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1713),
.Y(n_1751)
);

NOR2xp67_ASAP7_75t_L g1752 ( 
.A(n_1716),
.B(n_1670),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1701),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1693),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1707),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1735),
.B(n_1691),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1722),
.A2(n_1708),
.B(n_1707),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1745),
.B(n_1714),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1720),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1755),
.A2(n_1691),
.B1(n_1707),
.B2(n_1661),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1727),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

NAND2x1p5_ASAP7_75t_L g1764 ( 
.A(n_1748),
.B(n_1687),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1755),
.B(n_1712),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1740),
.B(n_1704),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1723),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1723),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1752),
.A2(n_1663),
.B1(n_1645),
.B2(n_1674),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1735),
.B(n_1692),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1721),
.B(n_1715),
.Y(n_1771)
);

OAI21xp33_ASAP7_75t_L g1772 ( 
.A1(n_1746),
.A2(n_1636),
.B(n_1715),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1720),
.B(n_1704),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1725),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1725),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1727),
.Y(n_1776)
);

AND2x2_ASAP7_75t_SL g1777 ( 
.A(n_1730),
.B(n_1709),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1728),
.B(n_1706),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1752),
.A2(n_1674),
.B1(n_1703),
.B2(n_1636),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1728),
.B(n_1706),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1729),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1741),
.B(n_1736),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1732),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1741),
.B(n_1688),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1732),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1738),
.B(n_1711),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1736),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1749),
.B(n_1692),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1733),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1742),
.A2(n_1716),
.B(n_1675),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1733),
.Y(n_1791)
);

NOR4xp25_ASAP7_75t_SL g1792 ( 
.A(n_1724),
.B(n_1655),
.C(n_1699),
.D(n_1694),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1729),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1749),
.B(n_1737),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1738),
.B(n_1711),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1745),
.B(n_1686),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1743),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1743),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1726),
.B(n_1688),
.Y(n_1800)
);

NAND2x1p5_ASAP7_75t_L g1801 ( 
.A(n_1748),
.B(n_1703),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1750),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1764),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1785),
.Y(n_1804)
);

AOI222xp33_ASAP7_75t_L g1805 ( 
.A1(n_1772),
.A2(n_1730),
.B1(n_1734),
.B2(n_1731),
.C1(n_1718),
.C2(n_1719),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1760),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1785),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1758),
.B(n_1731),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1782),
.B(n_1718),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1742),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1770),
.B(n_1730),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1765),
.B(n_1731),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1761),
.B(n_1719),
.C(n_1751),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1756),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1777),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1767),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1756),
.B(n_1742),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1779),
.A2(n_1742),
.B1(n_1748),
.B2(n_1734),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1768),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1769),
.A2(n_1748),
.B1(n_1734),
.B2(n_1751),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1757),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1774),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1773),
.B(n_1726),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1775),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1795),
.B(n_1764),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1757),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1783),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1789),
.Y(n_1828)
);

AO21x2_ASAP7_75t_L g1829 ( 
.A1(n_1762),
.A2(n_1724),
.B(n_1729),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1791),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1795),
.B(n_1737),
.Y(n_1831)
);

INVx4_ASAP7_75t_L g1832 ( 
.A(n_1801),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1762),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1763),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1763),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1770),
.B(n_1801),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1776),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1793),
.B(n_1754),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1815),
.B(n_1793),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1806),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1836),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1804),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1804),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1807),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1807),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1826),
.B(n_1771),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1821),
.B(n_1814),
.Y(n_1848)
);

AOI32xp33_ASAP7_75t_L g1849 ( 
.A1(n_1808),
.A2(n_1793),
.A3(n_1771),
.B1(n_1802),
.B2(n_1798),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1816),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1820),
.A2(n_1790),
.B1(n_1792),
.B2(n_1787),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1816),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1819),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1818),
.A2(n_1750),
.B1(n_1799),
.B2(n_1802),
.C(n_1766),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1813),
.A2(n_1778),
.B1(n_1780),
.B2(n_1802),
.C(n_1784),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1815),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1803),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1810),
.A2(n_1759),
.B1(n_1800),
.B2(n_1750),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1825),
.B(n_1788),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1819),
.Y(n_1860)
);

OAI31xp33_ASAP7_75t_L g1861 ( 
.A1(n_1810),
.A2(n_1655),
.A3(n_1750),
.B(n_1627),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1825),
.B(n_1786),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1836),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1817),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1822),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1832),
.B(n_1796),
.C(n_1786),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1840),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1840),
.B(n_1817),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1841),
.B(n_1823),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1850),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1841),
.B(n_1831),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1847),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1852),
.Y(n_1873)
);

AND2x4_ASAP7_75t_SL g1874 ( 
.A(n_1842),
.B(n_1832),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1848),
.B(n_1812),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1856),
.B(n_1831),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1863),
.B(n_1811),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1864),
.B(n_1811),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1853),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_SL g1880 ( 
.A1(n_1851),
.A2(n_1832),
.B1(n_1811),
.B2(n_1839),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1859),
.B(n_1839),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1843),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1844),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1857),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1862),
.B(n_1839),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1860),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1845),
.B(n_1809),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1855),
.B(n_1822),
.Y(n_1888)
);

OAI21xp33_ASAP7_75t_L g1889 ( 
.A1(n_1880),
.A2(n_1884),
.B(n_1871),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1871),
.B(n_1846),
.Y(n_1890)
);

AOI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1888),
.A2(n_1849),
.B1(n_1866),
.B2(n_1854),
.C(n_1865),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1868),
.B(n_1837),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_SL g1893 ( 
.A(n_1869),
.B(n_1861),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1869),
.B(n_1809),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1872),
.A2(n_1861),
.B(n_1858),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1867),
.A2(n_1827),
.B(n_1828),
.C(n_1824),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1878),
.A2(n_1837),
.B1(n_1797),
.B2(n_1830),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1872),
.A2(n_1827),
.B(n_1824),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1876),
.A2(n_1830),
.B(n_1828),
.Y(n_1899)
);

AOI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1875),
.A2(n_1834),
.B(n_1833),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1889),
.B(n_1867),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1892),
.B(n_1868),
.Y(n_1902)
);

AO22x1_ASAP7_75t_L g1903 ( 
.A1(n_1895),
.A2(n_1877),
.B1(n_1883),
.B2(n_1882),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1890),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_L g1905 ( 
.A(n_1891),
.B(n_1877),
.C(n_1882),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1894),
.B(n_1885),
.Y(n_1906)
);

AND4x1_ASAP7_75t_L g1907 ( 
.A(n_1893),
.B(n_1870),
.C(n_1886),
.D(n_1873),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1896),
.B(n_1883),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1899),
.B(n_1885),
.Y(n_1909)
);

INVxp67_ASAP7_75t_L g1910 ( 
.A(n_1897),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1900),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1883),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1902),
.B(n_1881),
.Y(n_1913)
);

NAND4xp75_ASAP7_75t_L g1914 ( 
.A(n_1901),
.B(n_1898),
.C(n_1881),
.D(n_1879),
.Y(n_1914)
);

OAI211xp5_ASAP7_75t_L g1915 ( 
.A1(n_1905),
.A2(n_1875),
.B(n_1887),
.C(n_1874),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1903),
.B(n_1887),
.C(n_1874),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_1834),
.C(n_1833),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1912),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1913),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1914),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1917),
.Y(n_1921)
);

CKINVDCx20_ASAP7_75t_R g1922 ( 
.A(n_1915),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1916),
.Y(n_1923)
);

NOR3xp33_ASAP7_75t_SL g1924 ( 
.A(n_1915),
.B(n_1904),
.C(n_1909),
.Y(n_1924)
);

NAND4xp75_ASAP7_75t_L g1925 ( 
.A(n_1924),
.B(n_1911),
.C(n_1906),
.D(n_1907),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1918),
.B(n_1922),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1923),
.B(n_1919),
.Y(n_1927)
);

NAND3xp33_ASAP7_75t_SL g1928 ( 
.A(n_1924),
.B(n_1910),
.C(n_1838),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1920),
.B(n_1796),
.Y(n_1929)
);

AOI31xp33_ASAP7_75t_L g1930 ( 
.A1(n_1921),
.A2(n_1540),
.A3(n_1835),
.B(n_1838),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1927),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1926),
.Y(n_1932)
);

XNOR2x1_ASAP7_75t_L g1933 ( 
.A(n_1925),
.B(n_1627),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1931),
.Y(n_1934)
);

OAI322xp33_ASAP7_75t_L g1935 ( 
.A1(n_1934),
.A2(n_1932),
.A3(n_1933),
.B1(n_1931),
.B2(n_1928),
.C1(n_1930),
.C2(n_1929),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1935),
.A2(n_1934),
.B1(n_1835),
.B2(n_1829),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1935),
.B(n_1829),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1937),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1936),
.A2(n_1829),
.B1(n_1794),
.B2(n_1781),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1938),
.A2(n_1794),
.B1(n_1781),
.B2(n_1776),
.Y(n_1940)
);

AOI221x1_ASAP7_75t_L g1941 ( 
.A1(n_1939),
.A2(n_1739),
.B1(n_1744),
.B2(n_1747),
.C(n_1754),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1940),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_L g1943 ( 
.A(n_1941),
.B(n_1744),
.C(n_1739),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1942),
.A2(n_1747),
.B1(n_1744),
.B2(n_1739),
.Y(n_1944)
);

OAI221xp5_ASAP7_75t_R g1945 ( 
.A1(n_1944),
.A2(n_1943),
.B1(n_1441),
.B2(n_1747),
.C(n_1754),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1582),
.B(n_1595),
.C(n_1753),
.Y(n_1946)
);


endmodule