module fake_aes_8080_n_794 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_794);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_794;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_L g101 ( .A(n_33), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_1), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_38), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_23), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_66), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_40), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_88), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_43), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_4), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_99), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_16), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_30), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_95), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_61), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_81), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_83), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_85), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_31), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_9), .Y(n_120) );
BUFx5_ASAP7_75t_L g121 ( .A(n_71), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_82), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_69), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_26), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_58), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_68), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_41), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_9), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_18), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_8), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_51), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_26), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_64), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_91), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_23), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_5), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_13), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_4), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_96), .Y(n_139) );
BUFx10_ASAP7_75t_L g140 ( .A(n_65), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_22), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_20), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_59), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_131), .B(n_0), .Y(n_145) );
BUFx8_ASAP7_75t_SL g146 ( .A(n_126), .Y(n_146) );
BUFx12f_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_107), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_101), .B(n_0), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_102), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_123), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_121), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_141), .B(n_1), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_118), .Y(n_161) );
BUFx12f_ASAP7_75t_L g162 ( .A(n_123), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_112), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_102), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_141), .Y(n_167) );
OAI22xp33_ASAP7_75t_L g168 ( .A1(n_161), .A2(n_103), .B1(n_143), .B2(n_104), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_162), .Y(n_169) );
OAI22xp33_ASAP7_75t_L g170 ( .A1(n_161), .A2(n_103), .B1(n_143), .B2(n_104), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_161), .A2(n_124), .B1(n_120), .B2(n_119), .Y(n_171) );
OR2x6_ASAP7_75t_L g172 ( .A(n_147), .B(n_106), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_161), .A2(n_109), .B1(n_142), .B2(n_136), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_150), .A2(n_137), .B1(n_113), .B2(n_138), .Y(n_175) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_152), .B(n_125), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_150), .B(n_135), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_150), .B(n_111), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_165), .A2(n_132), .B1(n_129), .B2(n_130), .Y(n_180) );
OAI22xp33_ASAP7_75t_SL g181 ( .A1(n_145), .A2(n_128), .B1(n_139), .B2(n_108), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_165), .B(n_105), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_165), .A2(n_105), .B1(n_139), .B2(n_108), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_149), .A2(n_115), .B1(n_144), .B2(n_133), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_152), .B(n_115), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_145), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_145), .A2(n_134), .B1(n_127), .B2(n_122), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_152), .B(n_157), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_152), .B(n_2), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_152), .B(n_110), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_149), .A2(n_117), .B1(n_116), .B2(n_114), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_149), .A2(n_121), .B1(n_6), .B2(n_7), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
BUFx6f_ASAP7_75t_SL g194 ( .A(n_152), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_146), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
BUFx6f_ASAP7_75t_SL g197 ( .A(n_152), .Y(n_197) );
AO22x2_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_3), .B1(n_6), .B2(n_7), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_159), .A2(n_121), .B1(n_10), .B2(n_11), .Y(n_200) );
NAND3x1_ASAP7_75t_L g201 ( .A(n_146), .B(n_8), .C(n_10), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_121), .B1(n_12), .B2(n_13), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_159), .A2(n_11), .B1(n_12), .B2(n_14), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_152), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_205) );
AOI22x1_ASAP7_75t_SL g206 ( .A1(n_146), .A2(n_15), .B1(n_17), .B2(n_18), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_157), .B(n_17), .Y(n_208) );
NAND3x1_ASAP7_75t_L g209 ( .A(n_148), .B(n_19), .C(n_20), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_157), .B(n_19), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_157), .A2(n_21), .B1(n_22), .B2(n_24), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_157), .B(n_42), .Y(n_212) );
OR2x6_ASAP7_75t_L g213 ( .A(n_147), .B(n_21), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_147), .A2(n_24), .B1(n_25), .B2(n_27), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_182), .B(n_157), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_185), .B(n_157), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_172), .B(n_157), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_179), .B(n_147), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
XOR2x2_ASAP7_75t_L g220 ( .A(n_171), .B(n_147), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_196), .Y(n_221) );
XNOR2xp5_ASAP7_75t_L g222 ( .A(n_168), .B(n_148), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_202), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_207), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_200), .B(n_151), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_200), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_172), .B(n_148), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_203), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_203), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_204), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_169), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_183), .B(n_148), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_191), .B(n_163), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_172), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_176), .B(n_163), .Y(n_236) );
XNOR2x2_ASAP7_75t_L g237 ( .A(n_186), .B(n_163), .Y(n_237) );
XOR2xp5_ASAP7_75t_L g238 ( .A(n_195), .B(n_25), .Y(n_238) );
XNOR2xp5_ASAP7_75t_L g239 ( .A(n_170), .B(n_163), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_178), .B(n_151), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_198), .Y(n_241) );
NAND2x1p5_ASAP7_75t_L g242 ( .A(n_189), .B(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_198), .Y(n_244) );
INVxp33_ASAP7_75t_L g245 ( .A(n_180), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g246 ( .A(n_194), .B(n_151), .Y(n_246) );
NAND2xp33_ASAP7_75t_SL g247 ( .A(n_194), .B(n_151), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_173), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_191), .B(n_162), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_213), .Y(n_252) );
XOR2x2_ASAP7_75t_L g253 ( .A(n_201), .B(n_27), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_188), .B(n_151), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_184), .B(n_151), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_192), .B(n_151), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_184), .B(n_155), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_190), .B(n_167), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_210), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_197), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_197), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_193), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_214), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_211), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_199), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_174), .B(n_28), .Y(n_271) );
INVxp33_ASAP7_75t_L g272 ( .A(n_175), .Y(n_272) );
AND2x6_ASAP7_75t_L g273 ( .A(n_212), .B(n_155), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_206), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_181), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_187), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_233), .B(n_167), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_227), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_257), .B(n_155), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_256), .B(n_155), .Y(n_280) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_227), .B(n_154), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_219), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_232), .B(n_167), .Y(n_283) );
NAND3xp33_ASAP7_75t_SL g284 ( .A(n_274), .B(n_160), .C(n_156), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_221), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_265), .B(n_155), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_227), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_257), .B(n_217), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_231), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_217), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_217), .B(n_155), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_264), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_242), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_257), .B(n_155), .Y(n_298) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_226), .B(n_154), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_256), .B(n_155), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_236), .B(n_154), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_259), .B(n_154), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_236), .B(n_154), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_231), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_240), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_249), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_240), .B(n_156), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_215), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_264), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_259), .B(n_156), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_225), .B(n_156), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_276), .B(n_156), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_218), .B(n_167), .Y(n_316) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_226), .B(n_160), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_261), .B(n_160), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_276), .B(n_160), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_242), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_269), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_269), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_225), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_225), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_215), .B(n_160), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_216), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_288), .B(n_228), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_289), .B(n_241), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_228), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_322), .B(n_229), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_289), .B(n_230), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_288), .B(n_229), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_322), .B(n_230), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_282), .B(n_235), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_290), .Y(n_340) );
BUFx8_ASAP7_75t_SL g341 ( .A(n_289), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_288), .B(n_245), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_288), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_282), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_290), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_281), .B(n_235), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_282), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_281), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_285), .Y(n_349) );
INVx4_ASAP7_75t_L g350 ( .A(n_295), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_285), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_285), .Y(n_352) );
INVx6_ASAP7_75t_L g353 ( .A(n_295), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_295), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_281), .B(n_258), .Y(n_356) );
INVx6_ASAP7_75t_SL g357 ( .A(n_289), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_278), .B(n_241), .Y(n_358) );
NOR2xp33_ASAP7_75t_SL g359 ( .A(n_281), .B(n_244), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_329), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_353), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_344), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_344), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_329), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_350), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_350), .B(n_324), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_329), .Y(n_368) );
BUFx6f_ASAP7_75t_SL g369 ( .A(n_334), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_329), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_255), .B1(n_325), .B2(n_324), .Y(n_376) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_348), .B(n_324), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_329), .Y(n_378) );
BUFx6f_ASAP7_75t_SL g379 ( .A(n_334), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_346), .A2(n_266), .B1(n_237), .B2(n_275), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
INVx5_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
INVx8_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_346), .B(n_289), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_355), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_353), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_340), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_382), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_380), .A2(n_348), .B1(n_346), .B2(n_356), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_374), .Y(n_391) );
BUFx12f_ASAP7_75t_L g392 ( .A(n_382), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_369), .A2(n_237), .B1(n_359), .B2(n_356), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_382), .Y(n_394) );
CKINVDCx11_ASAP7_75t_R g395 ( .A(n_383), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_380), .A2(n_356), .B1(n_328), .B2(n_337), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_369), .A2(n_359), .B1(n_331), .B2(n_289), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_360), .Y(n_399) );
AOI22x1_ASAP7_75t_SL g400 ( .A1(n_383), .A2(n_248), .B1(n_251), .B2(n_252), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
AND2x4_ASAP7_75t_SL g402 ( .A(n_366), .B(n_350), .Y(n_402) );
INVx5_ASAP7_75t_L g403 ( .A(n_382), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_383), .A2(n_337), .B1(n_328), .B2(n_331), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_360), .Y(n_406) );
CKINVDCx6p67_ASAP7_75t_R g407 ( .A(n_382), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_383), .A2(n_337), .B1(n_328), .B2(n_331), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_363), .B(n_332), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_383), .A2(n_328), .B1(n_337), .B2(n_336), .Y(n_410) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_370), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_374), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_379), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_370), .Y(n_415) );
BUFx10_ASAP7_75t_L g416 ( .A(n_369), .Y(n_416) );
INVx5_ASAP7_75t_L g417 ( .A(n_382), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_383), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_369), .A2(n_299), .B1(n_317), .B2(n_337), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_383), .A2(n_328), .B1(n_337), .B2(n_336), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_373), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_363), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_383), .A2(n_338), .B1(n_332), .B2(n_339), .Y(n_423) );
BUFx10_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_363), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_367), .Y(n_426) );
INVx6_ASAP7_75t_L g427 ( .A(n_382), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_328), .B1(n_336), .B2(n_253), .Y(n_430) );
INVx6_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_369), .A2(n_253), .B1(n_275), .B2(n_299), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_430), .A2(n_369), .B1(n_379), .B2(n_382), .Y(n_433) );
CKINVDCx6p67_ASAP7_75t_R g434 ( .A(n_403), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_423), .A2(n_379), .B1(n_342), .B2(n_384), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_399), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_432), .A2(n_382), .B1(n_379), .B2(n_377), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_399), .B(n_364), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
OAI222xp33_ASAP7_75t_L g441 ( .A1(n_430), .A2(n_238), .B1(n_385), .B2(n_366), .C1(n_367), .C2(n_376), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_432), .A2(n_379), .B1(n_377), .B2(n_342), .Y(n_442) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_395), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_405), .B(n_364), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_416), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_403), .B(n_366), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_402), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_391), .B(n_375), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_423), .A2(n_379), .B1(n_377), .B2(n_357), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_419), .A2(n_377), .B1(n_366), .B2(n_385), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_419), .A2(n_377), .B1(n_357), .B2(n_384), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_401), .B(n_388), .Y(n_452) );
BUFx12f_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_390), .A2(n_271), .B1(n_268), .B2(n_267), .C1(n_239), .C2(n_222), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_393), .A2(n_239), .B(n_222), .Y(n_456) );
BUFx4f_ASAP7_75t_SL g457 ( .A(n_392), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_406), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_413), .A2(n_366), .B1(n_385), .B2(n_376), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_413), .A2(n_366), .B1(n_385), .B2(n_271), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_403), .A2(n_366), .B1(n_385), .B2(n_338), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_389), .A2(n_272), .B(n_270), .C(n_376), .Y(n_462) );
OAI21xp33_ASAP7_75t_L g463 ( .A1(n_393), .A2(n_385), .B(n_388), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_401), .B(n_388), .Y(n_464) );
OAI222xp33_ASAP7_75t_L g465 ( .A1(n_398), .A2(n_238), .B1(n_367), .B2(n_364), .C1(n_350), .C2(n_330), .Y(n_465) );
INVx5_ASAP7_75t_SL g466 ( .A(n_407), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_407), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_403), .A2(n_367), .B1(n_384), .B2(n_362), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_406), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_401), .B(n_367), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_403), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_412), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_412), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_396), .A2(n_357), .B1(n_317), .B2(n_299), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_412), .B(n_373), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_403), .A2(n_339), .B1(n_354), .B2(n_334), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_390), .A2(n_357), .B1(n_299), .B2(n_317), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g481 ( .A1(n_404), .A2(n_354), .B(n_284), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_403), .A2(n_243), .B1(n_220), .B2(n_277), .C1(n_283), .C2(n_298), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_425), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_417), .A2(n_362), .B1(n_387), .B2(n_334), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_394), .A2(n_220), .B(n_340), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_417), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_407), .A2(n_357), .B1(n_277), .B2(n_330), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_417), .A2(n_325), .B1(n_324), .B2(n_347), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_417), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_404), .A2(n_330), .B1(n_283), .B2(n_341), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_408), .A2(n_330), .B1(n_358), .B2(n_316), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_408), .A2(n_330), .B1(n_358), .B2(n_316), .Y(n_492) );
BUFx4f_ASAP7_75t_SL g493 ( .A(n_418), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_417), .Y(n_494) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_394), .A2(n_345), .B(n_284), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g496 ( .A1(n_394), .A2(n_345), .B(n_330), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_417), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_414), .B(n_373), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_414), .B(n_373), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_414), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_457), .A2(n_427), .B1(n_431), .B2(n_417), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_482), .A2(n_417), .B1(n_410), .B2(n_420), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_471), .B(n_421), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_466), .A2(n_431), .B1(n_427), .B2(n_389), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_456), .A2(n_420), .B1(n_410), .B2(n_428), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_485), .A2(n_428), .B1(n_431), .B2(n_427), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_466), .A2(n_431), .B1(n_427), .B2(n_389), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_435), .A2(n_409), .B1(n_426), .B2(n_429), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_433), .A2(n_426), .B1(n_424), .B2(n_416), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_455), .A2(n_424), .B1(n_416), .B2(n_409), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_435), .A2(n_426), .B1(n_416), .B2(n_424), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g512 ( .A1(n_465), .A2(n_402), .B(n_426), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_460), .A2(n_424), .B1(n_330), .B2(n_358), .Y(n_513) );
OAI222xp33_ASAP7_75t_L g514 ( .A1(n_459), .A2(n_400), .B1(n_429), .B2(n_421), .C1(n_365), .C2(n_386), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_448), .B(n_429), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_441), .B(n_250), .C(n_362), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_449), .A2(n_424), .B1(n_402), .B2(n_358), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_442), .A2(n_358), .B1(n_362), .B2(n_387), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_438), .A2(n_358), .B1(n_387), .B2(n_325), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_477), .A2(n_387), .B1(n_352), .B2(n_351), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_448), .B(n_452), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_480), .A2(n_400), .B1(n_347), .B2(n_352), .Y(n_522) );
OAI222xp33_ASAP7_75t_L g523 ( .A1(n_450), .A2(n_365), .B1(n_386), .B2(n_415), .C1(n_373), .C2(n_381), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_451), .A2(n_349), .B1(n_353), .B2(n_335), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_462), .A2(n_415), .B1(n_353), .B2(n_386), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_452), .B(n_381), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_466), .A2(n_371), .B1(n_361), .B2(n_368), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_464), .B(n_381), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_491), .A2(n_353), .B1(n_343), .B2(n_335), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_492), .A2(n_343), .B1(n_335), .B2(n_361), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_462), .A2(n_365), .B1(n_333), .B2(n_381), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_490), .A2(n_343), .B1(n_368), .B2(n_361), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_463), .A2(n_368), .B1(n_361), .B2(n_371), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_463), .A2(n_368), .B1(n_361), .B2(n_371), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_496), .A2(n_371), .B1(n_294), .B2(n_314), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_481), .A2(n_333), .B1(n_381), .B2(n_345), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_466), .A2(n_411), .B1(n_397), .B2(n_378), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_481), .A2(n_345), .B1(n_355), .B2(n_378), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_434), .A2(n_411), .B1(n_397), .B2(n_355), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_484), .B(n_153), .C(n_158), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_434), .A2(n_355), .B1(n_370), .B2(n_378), .Y(n_541) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_467), .A2(n_314), .B1(n_298), .B2(n_279), .C1(n_294), .C2(n_311), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_453), .A2(n_287), .B1(n_291), .B2(n_314), .Y(n_543) );
OAI222xp33_ASAP7_75t_L g544 ( .A1(n_468), .A2(n_314), .B1(n_298), .B2(n_279), .C1(n_311), .C2(n_167), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_437), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_453), .A2(n_287), .B1(n_291), .B2(n_298), .Y(n_546) );
OAI222xp33_ASAP7_75t_L g547 ( .A1(n_447), .A2(n_298), .B1(n_279), .B2(n_311), .C1(n_167), .C2(n_286), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_479), .A2(n_411), .B1(n_397), .B2(n_355), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_487), .A2(n_411), .B1(n_397), .B2(n_355), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_436), .A2(n_493), .B1(n_489), .B2(n_486), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_494), .A2(n_378), .B1(n_372), .B2(n_370), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_447), .A2(n_378), .B1(n_372), .B2(n_370), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_494), .A2(n_372), .B1(n_378), .B2(n_311), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_497), .A2(n_372), .B1(n_295), .B2(n_297), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_443), .A2(n_372), .B1(n_300), .B2(n_278), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_461), .A2(n_372), .B1(n_295), .B2(n_297), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_440), .B(n_153), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_458), .A2(n_153), .B1(n_158), .B2(n_164), .C(n_166), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_476), .B(n_153), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_445), .A2(n_320), .B1(n_295), .B2(n_297), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_445), .A2(n_297), .B1(n_320), .B2(n_310), .Y(n_561) );
OAI222xp33_ASAP7_75t_L g562 ( .A1(n_446), .A2(n_167), .B1(n_286), .B2(n_292), .C1(n_300), .C2(n_278), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_488), .A2(n_306), .B1(n_297), .B2(n_320), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_446), .A2(n_278), .B1(n_297), .B2(n_320), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_446), .A2(n_297), .B1(n_320), .B2(n_292), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_474), .A2(n_297), .B1(n_320), .B2(n_312), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_445), .A2(n_320), .B1(n_296), .B2(n_286), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_458), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_469), .B(n_153), .Y(n_569) );
OAI222xp33_ASAP7_75t_L g570 ( .A1(n_454), .A2(n_167), .B1(n_296), .B2(n_313), .C1(n_312), .C2(n_303), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_470), .B(n_28), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_474), .A2(n_313), .B1(n_306), .B2(n_273), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_470), .A2(n_167), .B1(n_315), .B2(n_319), .C1(n_313), .C2(n_304), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_474), .A2(n_273), .B1(n_315), .B2(n_319), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_454), .A2(n_293), .B1(n_290), .B2(n_305), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_474), .A2(n_273), .B1(n_323), .B2(n_321), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_472), .A2(n_153), .B1(n_158), .B2(n_164), .C(n_166), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_454), .B(n_29), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_500), .A2(n_472), .B1(n_483), .B2(n_473), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_473), .A2(n_273), .B1(n_323), .B2(n_321), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_495), .A2(n_293), .B1(n_303), .B2(n_301), .C(n_280), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_512), .A2(n_495), .B(n_500), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_521), .B(n_478), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_512), .A2(n_514), .B(n_501), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_536), .A2(n_444), .B1(n_439), .B2(n_164), .C(n_153), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_545), .B(n_478), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_503), .B(n_498), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_510), .A2(n_475), .B1(n_167), .B2(n_499), .C(n_498), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_578), .B(n_510), .C(n_579), .Y(n_589) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_504), .A2(n_499), .B(n_475), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_545), .B(n_29), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_571), .B(n_153), .C(n_158), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_516), .B(n_153), .C(n_158), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_538), .B(n_167), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_536), .B(n_158), .C(n_164), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_522), .B(n_30), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_568), .B(n_31), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_568), .B(n_32), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_502), .A2(n_293), .B1(n_290), .B2(n_305), .Y(n_599) );
OA211x2_ASAP7_75t_L g600 ( .A1(n_550), .A2(n_32), .B(n_33), .C(n_34), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_538), .B(n_167), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_503), .B(n_34), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_515), .B(n_35), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_508), .A2(n_158), .B1(n_164), .B2(n_166), .C(n_167), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_540), .B(n_158), .C(n_164), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_508), .A2(n_158), .B1(n_164), .B2(n_166), .C(n_304), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_526), .B(n_35), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g608 ( .A1(n_505), .A2(n_280), .B1(n_301), .B2(n_302), .C(n_304), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_569), .B(n_36), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_540), .B(n_164), .C(n_166), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_528), .B(n_37), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_531), .A2(n_164), .B1(n_166), .B2(n_302), .C(n_304), .Y(n_612) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_531), .A2(n_302), .B1(n_262), .B2(n_263), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_561), .B(n_166), .C(n_318), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_513), .B(n_38), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_560), .B(n_166), .C(n_318), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_555), .B(n_577), .C(n_558), .Y(n_617) );
NOR2x1_ASAP7_75t_SL g618 ( .A(n_565), .B(n_305), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_557), .B(n_307), .C(n_309), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_559), .B(n_39), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_537), .B(n_246), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_520), .A2(n_309), .B1(n_307), .B2(n_302), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_559), .B(n_40), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_506), .B(n_246), .C(n_247), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_44), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_543), .A2(n_247), .B1(n_262), .B2(n_263), .C(n_327), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_533), .B(n_45), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_529), .A2(n_323), .B1(n_321), .B2(n_273), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_535), .B(n_308), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_534), .B(n_46), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_530), .A2(n_323), .B1(n_321), .B2(n_273), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_573), .B(n_308), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_573), .B(n_308), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_542), .A2(n_326), .B(n_327), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_552), .B(n_47), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_507), .A2(n_326), .B(n_327), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_563), .B(n_48), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_547), .B(n_260), .C(n_49), .Y(n_638) );
OAI221xp5_ASAP7_75t_SL g639 ( .A1(n_543), .A2(n_546), .B1(n_524), .B2(n_519), .C(n_518), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_517), .B(n_50), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_523), .A2(n_52), .B1(n_53), .B2(n_54), .C(n_55), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_552), .B(n_56), .Y(n_642) );
OA21x2_ASAP7_75t_L g643 ( .A1(n_548), .A2(n_57), .B(n_60), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_527), .B(n_62), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_532), .B(n_63), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_509), .B(n_67), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_544), .B(n_72), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_581), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_525), .B(n_76), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_565), .B(n_77), .C(n_78), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_549), .B(n_79), .C(n_80), .Y(n_651) );
OA211x2_ASAP7_75t_L g652 ( .A1(n_556), .A2(n_84), .B(n_86), .C(n_87), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_541), .B(n_89), .C(n_90), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_567), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_541), .B(n_98), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g656 ( .A1(n_570), .A2(n_100), .B(n_562), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_564), .A2(n_575), .B(n_539), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_553), .B(n_551), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_554), .B(n_575), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_583), .B(n_566), .Y(n_660) );
AO21x1_ASAP7_75t_SL g661 ( .A1(n_582), .A2(n_572), .B(n_574), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_586), .Y(n_662) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_584), .B(n_576), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_656), .A2(n_580), .B(n_636), .C(n_644), .Y(n_664) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_618), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_589), .A2(n_615), .B(n_657), .C(n_602), .Y(n_666) );
NOR3xp33_ASAP7_75t_SL g667 ( .A(n_644), .B(n_596), .C(n_639), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_596), .B(n_603), .C(n_598), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_590), .B(n_619), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_593), .B(n_617), .C(n_641), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_648), .B(n_658), .C(n_592), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_591), .B(n_597), .C(n_620), .Y(n_672) );
NAND4xp75_ASAP7_75t_L g673 ( .A(n_600), .B(n_652), .C(n_607), .D(n_611), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_648), .B(n_595), .C(n_613), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_585), .B(n_616), .C(n_604), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_608), .B(n_623), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_655), .B(n_642), .Y(n_677) );
NAND4xp75_ASAP7_75t_L g678 ( .A(n_659), .B(n_625), .C(n_643), .D(n_634), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_594), .B(n_601), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_609), .B(n_626), .C(n_647), .Y(n_680) );
NOR3xp33_ASAP7_75t_SL g681 ( .A(n_647), .B(n_614), .C(n_650), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_638), .B(n_640), .C(n_649), .Y(n_682) );
NAND4xp75_ASAP7_75t_L g683 ( .A(n_643), .B(n_635), .C(n_601), .D(n_621), .Y(n_683) );
NAND4xp75_ASAP7_75t_L g684 ( .A(n_621), .B(n_612), .C(n_630), .D(n_627), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_637), .B(n_646), .C(n_653), .Y(n_685) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_654), .B(n_645), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_599), .A2(n_633), .B1(n_632), .B2(n_629), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_606), .B(n_654), .C(n_605), .Y(n_688) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_610), .B(n_651), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_622), .A2(n_631), .B(n_628), .C(n_624), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_588), .A2(n_589), .B1(n_516), .B2(n_502), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_656), .A2(n_584), .B(n_644), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_584), .B(n_589), .C(n_657), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_588), .A2(n_589), .B1(n_516), .B2(n_502), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_584), .B(n_589), .C(n_657), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_596), .B(n_656), .C(n_584), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_589), .B(n_443), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_588), .A2(n_589), .B1(n_516), .B2(n_502), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_656), .A2(n_584), .B(n_644), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_587), .B(n_583), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_589), .A2(n_456), .B1(n_510), .B2(n_430), .Y(n_701) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_584), .B(n_644), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_587), .B(n_583), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_587), .B(n_583), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_584), .A2(n_656), .B(n_636), .C(n_512), .Y(n_705) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_584), .B(n_644), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_588), .A2(n_589), .B1(n_516), .B2(n_502), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_584), .B(n_589), .C(n_657), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_587), .B(n_583), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g710 ( .A1(n_584), .A2(n_656), .B(n_512), .C(n_636), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_586), .Y(n_711) );
NOR4xp25_ASAP7_75t_L g712 ( .A(n_693), .B(n_708), .C(n_695), .D(n_666), .Y(n_712) );
XOR2x2_ASAP7_75t_L g713 ( .A(n_702), .B(n_706), .Y(n_713) );
NOR4xp25_ASAP7_75t_L g714 ( .A(n_666), .B(n_705), .C(n_697), .D(n_692), .Y(n_714) );
NOR4xp25_ASAP7_75t_L g715 ( .A(n_705), .B(n_699), .C(n_701), .D(n_664), .Y(n_715) );
XOR2xp5_ASAP7_75t_L g716 ( .A(n_701), .B(n_673), .Y(n_716) );
XNOR2x1_ASAP7_75t_L g717 ( .A(n_678), .B(n_684), .Y(n_717) );
XNOR2x2_ASAP7_75t_L g718 ( .A(n_683), .B(n_674), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_662), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_670), .B(n_696), .C(n_710), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_711), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_665), .B(n_696), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_700), .B(n_703), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_704), .B(n_709), .Y(n_724) );
INVx4_ASAP7_75t_SL g725 ( .A(n_677), .Y(n_725) );
OAI31xp33_ASAP7_75t_L g726 ( .A1(n_664), .A2(n_690), .A3(n_669), .B(n_663), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_660), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_679), .Y(n_728) );
NAND4xp75_ASAP7_75t_L g729 ( .A(n_667), .B(n_686), .C(n_681), .D(n_689), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_671), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_672), .B(n_668), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_672), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_668), .B(n_687), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_691), .B(n_707), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_686), .Y(n_735) );
BUFx3_ASAP7_75t_L g736 ( .A(n_688), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_736), .B(n_676), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_722), .Y(n_738) );
INVxp67_ASAP7_75t_L g739 ( .A(n_731), .Y(n_739) );
INVxp67_ASAP7_75t_L g740 ( .A(n_732), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_729), .A2(n_680), .B1(n_698), .B2(n_694), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_727), .B(n_730), .Y(n_742) );
INVx1_ASAP7_75t_SL g743 ( .A(n_713), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_719), .Y(n_744) );
XNOR2x1_ASAP7_75t_L g745 ( .A(n_729), .B(n_675), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_725), .Y(n_746) );
OA22x2_ASAP7_75t_L g747 ( .A1(n_716), .A2(n_690), .B1(n_661), .B2(n_680), .Y(n_747) );
INVx4_ASAP7_75t_L g748 ( .A(n_713), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_721), .Y(n_749) );
XOR2x2_ASAP7_75t_L g750 ( .A(n_716), .B(n_682), .Y(n_750) );
INVx4_ASAP7_75t_L g751 ( .A(n_713), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_728), .B(n_685), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_732), .Y(n_753) );
AOI22x1_ASAP7_75t_SL g754 ( .A1(n_748), .A2(n_751), .B1(n_743), .B2(n_730), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_747), .A2(n_720), .B1(n_717), .B2(n_715), .Y(n_755) );
INVx1_ASAP7_75t_SL g756 ( .A(n_752), .Y(n_756) );
OA22x2_ASAP7_75t_L g757 ( .A1(n_748), .A2(n_735), .B1(n_734), .B2(n_718), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_751), .A2(n_717), .B1(n_724), .B2(n_723), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_744), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_751), .A2(n_717), .B1(n_724), .B2(n_723), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_749), .Y(n_761) );
INVx3_ASAP7_75t_L g762 ( .A(n_746), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_747), .A2(n_715), .B1(n_714), .B2(n_712), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_755), .A2(n_738), .B1(n_747), .B2(n_746), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_759), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_761), .Y(n_766) );
BUFx2_ASAP7_75t_L g767 ( .A(n_762), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_756), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_762), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_768), .Y(n_770) );
OAI22x1_ASAP7_75t_L g771 ( .A1(n_767), .A2(n_763), .B1(n_754), .B2(n_741), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_767), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_769), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_764), .A2(n_745), .B1(n_760), .B2(n_758), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_772), .Y(n_775) );
AND4x1_ASAP7_75t_L g776 ( .A(n_774), .B(n_714), .C(n_712), .D(n_726), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_770), .Y(n_777) );
OR2x2_ASAP7_75t_L g778 ( .A(n_775), .B(n_742), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_775), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_777), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_780), .A2(n_771), .B1(n_745), .B2(n_757), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_778), .Y(n_782) );
AO22x1_ASAP7_75t_L g783 ( .A1(n_782), .A2(n_779), .B1(n_737), .B2(n_736), .Y(n_783) );
AND4x1_ASAP7_75t_L g784 ( .A(n_781), .B(n_726), .C(n_737), .D(n_776), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_783), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_784), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_785), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_787), .Y(n_788) );
NAND4xp25_ASAP7_75t_L g789 ( .A(n_788), .B(n_786), .C(n_736), .D(n_773), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_789), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_790), .A2(n_739), .B1(n_750), .B2(n_757), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_791), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_792), .A2(n_740), .B1(n_753), .B2(n_765), .C(n_766), .Y(n_793) );
AOI211xp5_ASAP7_75t_L g794 ( .A1(n_793), .A2(n_733), .B(n_752), .C(n_750), .Y(n_794) );
endmodule