module fake_jpeg_15661_n_70 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_26),
.B(n_29),
.C(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_41),
.B1(n_21),
.B2(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_26),
.B1(n_15),
.B2(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_2),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_3),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_6),
.Y(n_55)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_47),
.C(n_59),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_50),
.B(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_58),
.B1(n_61),
.B2(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_64),
.B1(n_58),
.B2(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_12),
.B1(n_14),
.B2(n_18),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_20),
.Y(n_70)
);


endmodule