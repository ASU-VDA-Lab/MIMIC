module fake_jpeg_2817_n_690 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_690);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_690;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_62),
.Y(n_171)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_71),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_66),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_23),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_70),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_73),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_20),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_74),
.B(n_33),
.Y(n_161)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_82),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_23),
.A2(n_31),
.B1(n_26),
.B2(n_22),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_84),
.A2(n_45),
.B1(n_49),
.B2(n_52),
.Y(n_151)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_85),
.Y(n_223)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_91),
.Y(n_229)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_92),
.Y(n_154)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_98),
.Y(n_226)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_25),
.B(n_9),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_131),
.Y(n_157)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_24),
.B(n_19),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

BUFx2_ASAP7_75t_SL g215 ( 
.A(n_132),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_135),
.A2(n_156),
.B(n_174),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_23),
.B1(n_45),
.B2(n_49),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_141),
.A2(n_153),
.B1(n_202),
.B2(n_221),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_66),
.B(n_57),
.C(n_55),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_143),
.B(n_12),
.C(n_14),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_74),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_144),
.A2(n_152),
.B1(n_158),
.B2(n_160),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_151),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_110),
.B1(n_104),
.B2(n_106),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_49),
.B1(n_34),
.B2(n_24),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_69),
.B(n_57),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_65),
.A2(n_25),
.B1(n_28),
.B2(n_35),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_71),
.A2(n_55),
.B1(n_41),
.B2(n_47),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_161),
.B(n_163),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_47),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_168),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_109),
.A2(n_33),
.B1(n_46),
.B2(n_52),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_170),
.A2(n_172),
.B1(n_182),
.B2(n_187),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_111),
.A2(n_48),
.B1(n_34),
.B2(n_28),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_94),
.B(n_32),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_59),
.B(n_35),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_179),
.B(n_184),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_60),
.A2(n_50),
.B1(n_32),
.B2(n_48),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_67),
.B(n_50),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_70),
.A2(n_98),
.B1(n_72),
.B2(n_73),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_120),
.A2(n_30),
.B(n_34),
.C(n_54),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_101),
.B(n_19),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_81),
.B(n_9),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_216),
.B(n_224),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_82),
.A2(n_11),
.B1(n_18),
.B2(n_17),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_217),
.A2(n_219),
.B1(n_224),
.B2(n_231),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_87),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_132),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_116),
.B(n_8),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_117),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_233),
.Y(n_334)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_138),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_237),
.B(n_263),
.Y(n_326)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_238),
.Y(n_360)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

AO22x1_ASAP7_75t_SL g243 ( 
.A1(n_168),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_243),
.Y(n_322)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_244),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_186),
.B(n_12),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_245),
.B(n_253),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_246),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_248),
.B(n_250),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_249),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_252),
.B(n_282),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_147),
.B(n_12),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_254),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_139),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_255),
.B(n_259),
.Y(n_345)
);

OR2x2_ASAP7_75t_SL g256 ( 
.A(n_156),
.B(n_13),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_256),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_215),
.Y(n_257)
);

INVx4_ASAP7_75t_SL g337 ( 
.A(n_257),
.Y(n_337)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_260),
.A2(n_274),
.B1(n_319),
.B2(n_257),
.Y(n_368)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_261),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_145),
.Y(n_262)
);

INVx8_ASAP7_75t_L g373 ( 
.A(n_262),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_194),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_140),
.B(n_157),
.C(n_166),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_267),
.B(n_314),
.C(n_275),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_202),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_269),
.B(n_287),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_136),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_270),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_272),
.B(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_144),
.B(n_1),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_273),
.B(n_299),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_170),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_195),
.B(n_4),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_275),
.Y(n_355)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_154),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_276),
.Y(n_381)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_176),
.Y(n_278)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_226),
.Y(n_279)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_232),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_293),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_154),
.B(n_4),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_209),
.Y(n_285)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_285),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_223),
.A2(n_5),
.B1(n_218),
.B2(n_167),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_286),
.A2(n_292),
.B1(n_304),
.B2(n_310),
.Y(n_349)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_201),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_288),
.B(n_295),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_152),
.A2(n_5),
.B1(n_187),
.B2(n_231),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_289),
.A2(n_308),
.B1(n_271),
.B2(n_282),
.Y(n_353)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_205),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_298),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_134),
.A2(n_5),
.B1(n_173),
.B2(n_177),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_232),
.Y(n_293)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_133),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_296),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_171),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_301),
.Y(n_354)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_178),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_199),
.B(n_206),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_307),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_171),
.A2(n_228),
.B1(n_137),
.B2(n_230),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_303),
.A2(n_316),
.B1(n_213),
.B2(n_262),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_155),
.A2(n_164),
.B1(n_159),
.B2(n_133),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_150),
.B(n_229),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_305),
.B(n_306),
.Y(n_364)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_153),
.A2(n_141),
.B1(n_221),
.B2(n_210),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_190),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_311),
.Y(n_343)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_137),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_190),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_145),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_312),
.A2(n_313),
.B1(n_315),
.B2(n_318),
.Y(n_351)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_149),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_150),
.B(n_229),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_192),
.A2(n_210),
.B1(n_188),
.B2(n_226),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_149),
.A2(n_230),
.B1(n_189),
.B2(n_200),
.Y(n_316)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_188),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_213),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_SL g320 ( 
.A(n_252),
.B(n_189),
.C(n_200),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_344),
.C(n_313),
.Y(n_393)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_290),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_324),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_340),
.B1(n_346),
.B2(n_353),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_272),
.A2(n_283),
.B1(n_273),
.B2(n_317),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_236),
.A2(n_247),
.B(n_267),
.C(n_239),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_341),
.B(n_362),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_317),
.A2(n_236),
.B1(n_281),
.B2(n_234),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_256),
.A2(n_275),
.B(n_282),
.C(n_243),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_289),
.A2(n_268),
.B1(n_314),
.B2(n_310),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_366),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_318),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_268),
.A2(n_299),
.B1(n_303),
.B2(n_316),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_370),
.B1(n_233),
.B2(n_244),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_268),
.A2(n_243),
.B1(n_235),
.B2(n_238),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_319),
.A2(n_268),
.B1(n_309),
.B2(n_311),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_371),
.A2(n_382),
.B1(n_337),
.B2(n_380),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_314),
.A2(n_307),
.B1(n_261),
.B2(n_300),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g415 ( 
.A1(n_372),
.A2(n_279),
.B1(n_349),
.B2(n_337),
.Y(n_415)
);

OAI22x1_ASAP7_75t_L g377 ( 
.A1(n_296),
.A2(n_278),
.B1(n_241),
.B2(n_264),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_377),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_265),
.A2(n_302),
.B(n_277),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_380),
.A2(n_249),
.B(n_246),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_325),
.B(n_342),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_383),
.B(n_385),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_384),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_298),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_374),
.A2(n_240),
.B(n_266),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_386),
.A2(n_399),
.B(n_418),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_343),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_396),
.Y(n_438)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g469 ( 
.A(n_389),
.B(n_427),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_251),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_390),
.B(n_411),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_295),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_417),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_329),
.C(n_359),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_394),
.Y(n_457)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_378),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_397),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_353),
.A2(n_306),
.B1(n_312),
.B2(n_288),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_400),
.B1(n_414),
.B2(n_422),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_374),
.A2(n_242),
.B(n_285),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_401),
.B(n_404),
.Y(n_441)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_378),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_328),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_405),
.B(n_416),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_254),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_L g440 ( 
.A1(n_406),
.A2(n_421),
.B(n_326),
.Y(n_440)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_415),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_364),
.B(n_284),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_370),
.A2(n_276),
.B(n_294),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_413),
.A2(n_377),
.B(n_339),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_322),
.A2(n_287),
.B1(n_291),
.B2(n_258),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_320),
.B(n_344),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_SL g418 ( 
.A(n_355),
.B(n_322),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_420),
.Y(n_474)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_357),
.B(n_338),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_348),
.A2(n_346),
.B1(n_369),
.B2(n_332),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_348),
.A2(n_332),
.B1(n_362),
.B2(n_376),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_423),
.A2(n_330),
.B1(n_365),
.B2(n_360),
.Y(n_471)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_323),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_424),
.B(n_430),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_331),
.A2(n_332),
.B1(n_341),
.B2(n_376),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_432),
.B1(n_422),
.B2(n_429),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_426),
.A2(n_381),
.B(n_338),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_336),
.B(n_379),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

BUFx5_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_345),
.A2(n_350),
.B1(n_382),
.B2(n_354),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_379),
.C(n_359),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_444),
.C(n_454),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_435),
.A2(n_471),
.B1(n_431),
.B2(n_430),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_391),
.A2(n_351),
.B1(n_367),
.B2(n_326),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_439),
.A2(n_442),
.B1(n_460),
.B2(n_473),
.Y(n_489)
);

OAI21xp33_ASAP7_75t_L g481 ( 
.A1(n_440),
.A2(n_432),
.B(n_421),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_391),
.A2(n_367),
.B1(n_357),
.B2(n_373),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_446),
.A2(n_448),
.B(n_458),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_409),
.A2(n_381),
.B(n_356),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_356),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_427),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_393),
.B(n_329),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_409),
.A2(n_347),
.B(n_361),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_387),
.B(n_334),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_470),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_400),
.A2(n_373),
.B1(n_352),
.B2(n_337),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_427),
.Y(n_463)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_383),
.B(n_385),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_465),
.B(n_450),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_395),
.B(n_347),
.C(n_334),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_475),
.C(n_420),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_360),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_425),
.A2(n_373),
.B1(n_365),
.B2(n_361),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_403),
.B(n_404),
.C(n_401),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_455),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_476),
.B(n_479),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_418),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_444),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_480),
.B(n_485),
.C(n_486),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_481),
.B(n_491),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_461),
.B(n_405),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_482),
.B(n_494),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_483),
.B(n_488),
.Y(n_535)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_484),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_433),
.B(n_396),
.C(n_407),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_410),
.C(n_392),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_447),
.Y(n_487)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_411),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_474),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_386),
.C(n_406),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_492),
.B(n_502),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_436),
.A2(n_413),
.B1(n_394),
.B2(n_406),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_493),
.A2(n_439),
.B1(n_463),
.B2(n_457),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_451),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_495),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_469),
.A2(n_399),
.B(n_389),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_496),
.A2(n_501),
.B(n_449),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_416),
.C(n_419),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_500),
.C(n_437),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_451),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_499),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_390),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_434),
.A2(n_394),
.B1(n_427),
.B2(n_414),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_507),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_438),
.B(n_427),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_458),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_SL g505 ( 
.A(n_437),
.B(n_388),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_510),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_424),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_467),
.B(n_397),
.Y(n_508)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_447),
.Y(n_509)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

XNOR2x2_ASAP7_75t_L g511 ( 
.A(n_435),
.B(n_431),
.Y(n_511)
);

A2O1A1O1Ixp25_ASAP7_75t_L g551 ( 
.A1(n_511),
.A2(n_456),
.B(n_428),
.C(n_402),
.D(n_339),
.Y(n_551)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_443),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_515),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_467),
.B(n_358),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_513),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_459),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_514),
.Y(n_537)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

OAI22x1_ASAP7_75t_L g516 ( 
.A1(n_501),
.A2(n_434),
.B1(n_441),
.B2(n_469),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_516),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_476),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_523),
.A2(n_525),
.B1(n_539),
.B2(n_544),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_478),
.B(n_441),
.C(n_464),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_528),
.C(n_529),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_489),
.A2(n_442),
.B1(n_434),
.B2(n_438),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_445),
.C(n_464),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_480),
.B(n_445),
.C(n_448),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_489),
.A2(n_434),
.B1(n_436),
.B2(n_452),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_534),
.B(n_488),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_536),
.B(n_479),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_493),
.A2(n_452),
.B1(n_473),
.B2(n_457),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_486),
.B(n_462),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_540),
.B(n_548),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_507),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_541),
.B(n_542),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_497),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_483),
.B(n_466),
.C(n_471),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_543),
.B(n_519),
.C(n_520),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_484),
.A2(n_462),
.B1(n_468),
.B2(n_470),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_496),
.A2(n_460),
.B1(n_453),
.B2(n_446),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_546),
.A2(n_550),
.B1(n_552),
.B2(n_539),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_547),
.A2(n_506),
.B(n_477),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_485),
.B(n_449),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_497),
.A2(n_431),
.B1(n_472),
.B2(n_456),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_551),
.A2(n_506),
.B(n_504),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_511),
.A2(n_412),
.B1(n_358),
.B2(n_330),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_554),
.A2(n_555),
.B(n_518),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_522),
.B(n_498),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_556),
.B(n_568),
.Y(n_589)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_517),
.Y(n_557)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_557),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_558),
.B(n_570),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_538),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_571),
.Y(n_590)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_538),
.Y(n_560)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_560),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_527),
.Y(n_561)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_561),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_562),
.B(n_574),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_525),
.A2(n_477),
.B1(n_490),
.B2(n_492),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_565),
.A2(n_573),
.B1(n_577),
.B2(n_583),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_566),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_530),
.B(n_502),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_526),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_585),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_535),
.B(n_500),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_547),
.A2(n_515),
.B(n_512),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_523),
.A2(n_487),
.B1(n_495),
.B2(n_509),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_549),
.B(n_412),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_535),
.B(n_408),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_575),
.B(n_576),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_521),
.B(n_520),
.Y(n_576)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_579),
.Y(n_605)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_580),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_581),
.B(n_584),
.C(n_549),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_537),
.B(n_532),
.Y(n_582)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_582),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_546),
.A2(n_518),
.B1(n_553),
.B2(n_534),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_543),
.B(n_528),
.C(n_548),
.Y(n_584)
);

AND3x1_ASAP7_75t_L g585 ( 
.A(n_516),
.B(n_536),
.C(n_551),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_545),
.Y(n_591)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_591),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_572),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_593),
.B(n_602),
.Y(n_626)
);

XNOR2x1_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_555),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_564),
.A2(n_518),
.B1(n_529),
.B2(n_540),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_599),
.A2(n_606),
.B1(n_610),
.B2(n_573),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_576),
.B(n_524),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_601),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_581),
.B(n_519),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_570),
.B(n_533),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_604),
.B(n_609),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_583),
.A2(n_526),
.B1(n_533),
.B2(n_560),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_579),
.B(n_561),
.Y(n_608)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_608),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_578),
.B(n_558),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_554),
.A2(n_565),
.B1(n_566),
.B2(n_571),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_590),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_612),
.B(n_613),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_589),
.B(n_575),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_596),
.B(n_569),
.Y(n_614)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_614),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_615),
.B(n_620),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_594),
.A2(n_585),
.B(n_567),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_616),
.A2(n_622),
.B(n_587),
.Y(n_636)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_596),
.Y(n_621)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_621),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_598),
.A2(n_578),
.B(n_563),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_611),
.Y(n_623)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_623),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_606),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_624),
.B(n_631),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_586),
.A2(n_563),
.B1(n_584),
.B2(n_574),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_602),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_601),
.C(n_592),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_628),
.B(n_592),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_604),
.B(n_562),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_609),
.Y(n_651)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_607),
.Y(n_630)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_630),
.Y(n_649)
);

BUFx24_ASAP7_75t_SL g631 ( 
.A(n_595),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_SL g632 ( 
.A(n_603),
.B(n_610),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_SL g639 ( 
.A(n_632),
.B(n_603),
.Y(n_639)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_588),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_633),
.B(n_605),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_599),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_634),
.B(n_635),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_636),
.B(n_641),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_639),
.B(n_642),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_615),
.A2(n_598),
.B(n_597),
.Y(n_641)
);

AOI21x1_ASAP7_75t_SL g655 ( 
.A1(n_641),
.A2(n_616),
.B(n_614),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_629),
.B(n_586),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_643),
.B(n_644),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_625),
.B(n_595),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_618),
.B(n_628),
.C(n_627),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_645),
.B(n_618),
.Y(n_661)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_648),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g654 ( 
.A(n_651),
.B(n_622),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_654),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_655),
.A2(n_636),
.B(n_637),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_634),
.B(n_620),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_656),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_650),
.A2(n_617),
.B1(n_619),
.B2(n_626),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_657),
.B(n_659),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_638),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_661),
.B(n_663),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_642),
.B(n_632),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_662),
.Y(n_673)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_640),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_664),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_645),
.B(n_643),
.C(n_646),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_665),
.B(n_644),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_658),
.B(n_649),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_668),
.B(n_672),
.Y(n_681)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_671),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_660),
.B(n_647),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_675),
.B(n_652),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_SL g676 ( 
.A1(n_667),
.A2(n_664),
.B(n_655),
.C(n_659),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_676),
.B(n_677),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_670),
.B(n_656),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_SL g682 ( 
.A1(n_678),
.A2(n_679),
.B(n_674),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_666),
.A2(n_637),
.B1(n_654),
.B2(n_653),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_682),
.B(n_676),
.Y(n_685)
);

O2A1O1Ixp5_ASAP7_75t_L g684 ( 
.A1(n_680),
.A2(n_674),
.B(n_639),
.C(n_673),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_684),
.B(n_681),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_SL g687 ( 
.A1(n_685),
.A2(n_686),
.B1(n_683),
.B2(n_669),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_653),
.B(n_662),
.Y(n_688)
);

XNOR2x2_ASAP7_75t_SL g689 ( 
.A(n_688),
.B(n_651),
.Y(n_689)
);

BUFx24_ASAP7_75t_SL g690 ( 
.A(n_689),
.Y(n_690)
);


endmodule