module fake_jpeg_6014_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_18),
.B(n_20),
.Y(n_23)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_28),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_18),
.C(n_14),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_33),
.C(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_36),
.Y(n_39)
);

AO22x1_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_22),
.B1(n_16),
.B2(n_17),
.Y(n_33)
);

FAx1_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_16),
.CI(n_19),
.CON(n_34),
.SN(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_15),
.B(n_8),
.C(n_9),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_35),
.B1(n_33),
.B2(n_15),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_19),
.C(n_22),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_46),
.B(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_34),
.B1(n_24),
.B2(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_38),
.B1(n_10),
.B2(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_43),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.C(n_2),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_1),
.B(n_10),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.C(n_6),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_2),
.C(n_6),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_7),
.Y(n_57)
);


endmodule