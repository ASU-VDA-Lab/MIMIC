module fake_jpeg_10688_n_420 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_420);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_420;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_0),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_19),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_58),
.B(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_63),
.B(n_65),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_28),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_38),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_29),
.B1(n_18),
.B2(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_1),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_32),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

INVx11_ASAP7_75t_SL g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_13),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_120),
.B1(n_18),
.B2(n_29),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_103),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_23),
.B1(n_36),
.B2(n_35),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_100),
.A2(n_52),
.B(n_39),
.C(n_20),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_117),
.Y(n_141)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_31),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_66),
.B1(n_64),
.B2(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_12),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_12),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_83),
.B1(n_70),
.B2(n_73),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_128),
.A2(n_129),
.B1(n_143),
.B2(n_150),
.Y(n_189)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_130),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_137),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_53),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_157),
.B(n_26),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_87),
.Y(n_133)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_91),
.A2(n_47),
.B(n_59),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_135),
.A2(n_163),
.B(n_106),
.Y(n_194)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_93),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_71),
.B1(n_50),
.B2(n_51),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_39),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_159),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_86),
.A2(n_43),
.B1(n_55),
.B2(n_60),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_153),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_44),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_68),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_95),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_22),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_22),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_165),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_43),
.B1(n_79),
.B2(n_36),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_45),
.B1(n_74),
.B2(n_115),
.Y(n_169)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_33),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_84),
.B1(n_115),
.B2(n_108),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_169),
.B1(n_172),
.B2(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_105),
.C(n_122),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_178),
.C(n_132),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_157),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_126),
.B1(n_87),
.B2(n_121),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_131),
.A2(n_126),
.B1(n_121),
.B2(n_98),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_105),
.C(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_192),
.Y(n_198)
);

NAND2x1_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_110),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_194),
.B(n_163),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_119),
.A3(n_125),
.B1(n_57),
.B2(n_110),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_125),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_95),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_144),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_199),
.B(n_209),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_165),
.B1(n_162),
.B2(n_143),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_208),
.B1(n_211),
.B2(n_215),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_204),
.C(n_188),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_135),
.C(n_155),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_221),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_129),
.B1(n_163),
.B2(n_133),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_142),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_212),
.B(n_227),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_163),
.B1(n_133),
.B2(n_148),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_151),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_213),
.B(n_216),
.Y(n_244)
);

OAI221xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_149),
.B1(n_130),
.B2(n_163),
.C(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_90),
.B1(n_145),
.B2(n_139),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_139),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_147),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_90),
.B1(n_160),
.B2(n_164),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_220),
.B1(n_169),
.B2(n_167),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_158),
.B1(n_146),
.B2(n_138),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_249),
.C(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_192),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_230),
.B(n_254),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_227),
.A3(n_198),
.B1(n_199),
.B2(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_255),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_206),
.B1(n_200),
.B2(n_204),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_235),
.A2(n_248),
.B1(n_136),
.B2(n_106),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_246),
.B1(n_214),
.B2(n_226),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_172),
.B1(n_176),
.B2(n_178),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_181),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_191),
.B1(n_197),
.B2(n_158),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_173),
.C(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_173),
.C(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_182),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_207),
.B(n_181),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_182),
.C(n_170),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_193),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_280),
.C(n_285),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_232),
.A2(n_205),
.B1(n_215),
.B2(n_221),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_258),
.A2(n_266),
.B1(n_273),
.B2(n_286),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_210),
.B(n_211),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_259),
.A2(n_261),
.B(n_264),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_210),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_213),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_263),
.B(n_239),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_220),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_265),
.A2(n_269),
.B1(n_272),
.B2(n_245),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_225),
.B1(n_201),
.B2(n_205),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_251),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_218),
.B1(n_184),
.B2(n_170),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_174),
.B(n_193),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_282),
.B(n_283),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_174),
.B1(n_146),
.B2(n_134),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_119),
.B1(n_193),
.B2(n_33),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_242),
.B(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_33),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_242),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_244),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_26),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_234),
.A2(n_26),
.B(n_22),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_20),
.B(n_3),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_92),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_235),
.A2(n_36),
.B1(n_20),
.B2(n_27),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_249),
.C(n_250),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_300),
.C(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_233),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_294),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_279),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_296),
.B(n_298),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_256),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_243),
.C(n_240),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_252),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_304),
.C(n_308),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_240),
.C(n_239),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_305),
.B(n_281),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_241),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_288),
.B(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_243),
.C(n_247),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_238),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_286),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_282),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_264),
.A2(n_245),
.B1(n_241),
.B2(n_36),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_271),
.B(n_308),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_318),
.B(n_333),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_273),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_334),
.Y(n_343)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_325),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_284),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_324),
.Y(n_342)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_326),
.A2(n_321),
.B1(n_324),
.B2(n_336),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_297),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_336),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_299),
.A2(n_264),
.B1(n_272),
.B2(n_269),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_329),
.A2(n_307),
.B1(n_282),
.B2(n_287),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_275),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_332),
.A2(n_274),
.B1(n_287),
.B2(n_300),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_306),
.B(n_304),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_270),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_333),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_292),
.C(n_289),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_340),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_303),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_344),
.A2(n_345),
.B1(n_349),
.B2(n_2),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_330),
.A2(n_323),
.B1(n_329),
.B2(n_332),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_318),
.A2(n_307),
.B(n_270),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_262),
.B(n_3),
.C(n_4),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_321),
.A2(n_305),
.B1(n_262),
.B2(n_27),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_316),
.C(n_327),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_353),
.C(n_317),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_327),
.C(n_331),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_355),
.A2(n_325),
.B1(n_320),
.B2(n_319),
.Y(n_366)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_358),
.B(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_346),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_361),
.Y(n_378)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_343),
.B(n_334),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_341),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_365),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_314),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_364),
.B(n_366),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_339),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_351),
.C(n_350),
.Y(n_372)
);

O2A1O1Ixp33_ASAP7_75t_SL g376 ( 
.A1(n_368),
.A2(n_370),
.B(n_341),
.C(n_349),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_369),
.A2(n_354),
.B(n_348),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_SL g370 ( 
.A1(n_347),
.A2(n_92),
.B(n_5),
.C(n_6),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_371),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_373),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_358),
.A2(n_348),
.B(n_352),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_374),
.A2(n_342),
.B(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_352),
.C(n_343),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_370),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_376),
.A2(n_383),
.B1(n_370),
.B2(n_5),
.Y(n_395)
);

INVx11_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_359),
.C(n_364),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_386),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_384),
.C(n_374),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_6),
.B(n_7),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_373),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_394),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_383),
.B(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_391),
.B(n_396),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_377),
.A2(n_378),
.B(n_382),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_392),
.A2(n_7),
.B(n_8),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_4),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_381),
.A2(n_378),
.B1(n_376),
.B2(n_6),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_387),
.A2(n_381),
.B(n_5),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_399),
.A2(n_404),
.B(n_8),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_401),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_9),
.B(n_11),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_390),
.B(n_395),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_408),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_398),
.B(n_393),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_411),
.Y(n_415)
);

O2A1O1Ixp33_ASAP7_75t_SL g410 ( 
.A1(n_403),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_410)
);

O2A1O1Ixp33_ASAP7_75t_SL g412 ( 
.A1(n_410),
.A2(n_402),
.B(n_400),
.C(n_11),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_414),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_406),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g417 ( 
.A(n_413),
.B(n_402),
.CI(n_9),
.CON(n_417),
.SN(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_417),
.B(n_415),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_417),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_416),
.Y(n_420)
);


endmodule