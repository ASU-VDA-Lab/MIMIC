module fake_aes_2409_n_659 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_659);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_659;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g79 ( .A(n_55), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_30), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_22), .Y(n_81) );
BUFx3_ASAP7_75t_L g82 ( .A(n_76), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_67), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_72), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_29), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_26), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_8), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_46), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_37), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_18), .Y(n_92) );
INVxp33_ASAP7_75t_L g93 ( .A(n_27), .Y(n_93) );
BUFx2_ASAP7_75t_L g94 ( .A(n_16), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_16), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_22), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_62), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_43), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_34), .Y(n_100) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_31), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_45), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_35), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_77), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_17), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_9), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_4), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_32), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_39), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_70), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_13), .B(n_36), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_6), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_60), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_56), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_38), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_5), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_42), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_73), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_41), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_4), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_115), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_101), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_79), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_94), .B(n_0), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
NOR2xp33_ASAP7_75t_R g133 ( .A(n_102), .B(n_24), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_94), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
NAND2xp33_ASAP7_75t_SL g136 ( .A(n_93), .B(n_109), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_107), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_122), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_119), .Y(n_139) );
NOR2xp33_ASAP7_75t_R g140 ( .A(n_82), .B(n_25), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_82), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_80), .B(n_0), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
NOR2xp67_ASAP7_75t_L g146 ( .A(n_92), .B(n_1), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_92), .B(n_2), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_82), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_108), .B(n_2), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_81), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_108), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_112), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_112), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_113), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_95), .B(n_3), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_87), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_84), .B(n_3), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_113), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_84), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_83), .B(n_47), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_88), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_80), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_87), .B(n_5), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_169), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_130), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_131), .B(n_104), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_128), .B(n_104), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_131), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_169), .B(n_125), .Y(n_176) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_169), .B(n_125), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_134), .B(n_106), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_151), .B(n_103), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_151), .B(n_103), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_153), .B(n_100), .Y(n_186) );
INVx8_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_169), .B(n_106), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_168), .B(n_90), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_153), .B(n_90), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_130), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_168), .B(n_97), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_155), .B(n_97), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_155), .B(n_105), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_157), .B(n_118), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_156), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_143), .B(n_105), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_130), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_148), .B(n_100), .Y(n_202) );
NAND3xp33_ASAP7_75t_L g203 ( .A(n_156), .B(n_118), .C(n_111), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_130), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_157), .B(n_99), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_148), .B(n_99), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_141), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_129), .B(n_110), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_129), .B(n_110), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_138), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_163), .A2(n_98), .B1(n_85), .B2(n_121), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_163), .B(n_98), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_145), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_152), .B(n_111), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_127), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_139), .B(n_96), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_152), .B(n_146), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_154), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_161), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_162), .B(n_96), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_170), .A2(n_144), .B(n_165), .C(n_149), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_175), .B(n_127), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_205), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_205), .B(n_139), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_172), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_196), .B(n_147), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_196), .B(n_191), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_223), .B(n_136), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_176), .A2(n_159), .B1(n_160), .B2(n_86), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_210), .B(n_116), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_190), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_198), .A2(n_114), .B1(n_85), .B2(n_86), .C(n_121), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_175), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_172), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_176), .B(n_166), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_176), .B(n_166), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_217), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_177), .Y(n_250) );
BUFx4_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
BUFx8_ASAP7_75t_L g252 ( .A(n_196), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_218), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_177), .B(n_166), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_177), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_218), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_191), .A2(n_166), .B1(n_124), .B2(n_91), .Y(n_257) );
NAND3xp33_ASAP7_75t_SL g258 ( .A(n_215), .B(n_140), .C(n_133), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_191), .B(n_166), .Y(n_259) );
AO22x1_ASAP7_75t_L g260 ( .A1(n_199), .A2(n_166), .B1(n_117), .B2(n_91), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_190), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_226), .Y(n_262) );
AND2x6_ASAP7_75t_L g263 ( .A(n_170), .B(n_117), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_191), .A2(n_89), .B1(n_123), .B2(n_120), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_192), .B(n_137), .Y(n_265) );
INVx5_ASAP7_75t_L g266 ( .A(n_170), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g267 ( .A(n_222), .B(n_6), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_211), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_226), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_195), .A2(n_89), .B1(n_120), .B2(n_123), .Y(n_270) );
AND2x6_ASAP7_75t_L g271 ( .A(n_188), .B(n_123), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_198), .B(n_120), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_227), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_195), .B(n_88), .Y(n_274) );
AND3x1_ASAP7_75t_L g275 ( .A(n_215), .B(n_88), .C(n_8), .Y(n_275) );
AO22x1_ASAP7_75t_L g276 ( .A1(n_195), .A2(n_84), .B1(n_9), .B2(n_10), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_192), .B(n_7), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_188), .B(n_84), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_187), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_187), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_188), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_203), .B(n_7), .C(n_10), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
BUFx8_ASAP7_75t_L g284 ( .A(n_195), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_174), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_188), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_174), .B(n_84), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_187), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_173), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_174), .B(n_11), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_229), .B(n_51), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_229), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_216), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_231), .B(n_180), .Y(n_295) );
INVx4_ASAP7_75t_L g296 ( .A(n_271), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_238), .A2(n_184), .B1(n_180), .B2(n_181), .Y(n_297) );
O2A1O1Ixp5_ASAP7_75t_L g298 ( .A1(n_260), .A2(n_186), .B(n_197), .C(n_207), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_289), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_252), .Y(n_300) );
BUFx4_ASAP7_75t_SL g301 ( .A(n_244), .Y(n_301) );
BUFx4f_ASAP7_75t_SL g302 ( .A(n_252), .Y(n_302) );
NAND3x1_ASAP7_75t_L g303 ( .A(n_264), .B(n_200), .C(n_202), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_247), .Y(n_304) );
BUFx4f_ASAP7_75t_SL g305 ( .A(n_284), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_249), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_246), .A2(n_213), .B(n_208), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_271), .A2(n_229), .B1(n_180), .B2(n_208), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_284), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_271), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_250), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_253), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_294), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
INVx5_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_262), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_269), .Y(n_317) );
BUFx12f_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_273), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_255), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_233), .B(n_221), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_266), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_235), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_237), .B(n_225), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_237), .B(n_225), .Y(n_328) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_255), .B(n_213), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_271), .Y(n_330) );
BUFx10_ASAP7_75t_L g331 ( .A(n_238), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_291), .B(n_225), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_281), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_281), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_277), .A2(n_211), .B1(n_221), .B2(n_182), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_266), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_279), .B(n_221), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_246), .A2(n_213), .B(n_214), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_285), .B(n_182), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_245), .B(n_183), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_261), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_251), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_248), .A2(n_214), .B(n_228), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_308), .A2(n_293), .B1(n_274), .B2(n_245), .Y(n_347) );
NAND2xp33_ASAP7_75t_R g348 ( .A(n_320), .B(n_280), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_308), .A2(n_274), .B1(n_270), .B2(n_272), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_304), .A2(n_236), .B1(n_263), .B2(n_287), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_311), .B(n_288), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_344), .B(n_265), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_307), .A2(n_278), .B(n_292), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_320), .B(n_234), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_336), .A2(n_272), .B1(n_290), .B2(n_292), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_318), .A2(n_240), .B1(n_234), .B2(n_267), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_318), .A2(n_240), .B1(n_258), .B2(n_259), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_313), .Y(n_358) );
NAND2xp33_ASAP7_75t_L g359 ( .A(n_310), .B(n_263), .Y(n_359) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_300), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_332), .A2(n_275), .B1(n_258), .B2(n_239), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_304), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_332), .A2(n_232), .B1(n_241), .B2(n_263), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_287), .Y(n_364) );
AND2x6_ASAP7_75t_L g365 ( .A(n_310), .B(n_259), .Y(n_365) );
INVx4_ASAP7_75t_SL g366 ( .A(n_310), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_305), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_309), .B(n_266), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_295), .A2(n_263), .B1(n_243), .B2(n_266), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_306), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_295), .A2(n_263), .B1(n_243), .B2(n_257), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_304), .A2(n_228), .B1(n_194), .B2(n_173), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_302), .A2(n_276), .B1(n_278), .B2(n_248), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_312), .A2(n_178), .B1(n_189), .B2(n_183), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_322), .B(n_230), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g376 ( .A1(n_298), .A2(n_319), .B(n_306), .C(n_314), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_312), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g378 ( .A(n_367), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_377), .B(n_341), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_361), .A2(n_297), .B1(n_327), .B2(n_328), .C(n_338), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_347), .A2(n_311), .B1(n_296), .B2(n_330), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_349), .A2(n_303), .B1(n_296), .B2(n_332), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_356), .A2(n_332), .B1(n_295), .B2(n_319), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_295), .B1(n_316), .B2(n_317), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_339), .B(n_345), .Y(n_386) );
OR2x6_ASAP7_75t_L g387 ( .A(n_351), .B(n_296), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_375), .A2(n_312), .B(n_303), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_372), .A2(n_296), .B1(n_317), .B2(n_316), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_321), .B1(n_314), .B2(n_340), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_321), .B1(n_340), .B2(n_341), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_351), .B(n_299), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_376), .A2(n_254), .B(n_282), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_340), .B1(n_333), .B2(n_334), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_355), .A2(n_330), .B1(n_329), .B2(n_310), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_340), .B1(n_333), .B2(n_334), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_329), .B1(n_310), .B2(n_338), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_363), .A2(n_333), .B1(n_334), .B2(n_323), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_374), .A2(n_329), .B1(n_310), .B2(n_338), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_354), .A2(n_338), .B1(n_282), .B2(n_323), .C(n_335), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_359), .A2(n_254), .B(n_342), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_346), .B(n_338), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_374), .A2(n_315), .B1(n_299), .B2(n_189), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_380), .B(n_373), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_383), .A2(n_358), .B(n_368), .C(n_364), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_386), .A2(n_324), .B(n_337), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_392), .B(n_373), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_392), .Y(n_410) );
AOI222xp33_ASAP7_75t_SL g411 ( .A1(n_390), .A2(n_360), .B1(n_301), .B2(n_14), .C1(n_15), .C2(n_17), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_380), .B(n_343), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_350), .B(n_342), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_389), .A2(n_350), .B(n_325), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_387), .Y(n_416) );
OA21x2_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_325), .B(n_326), .Y(n_417) );
OR2x6_ASAP7_75t_L g418 ( .A(n_387), .B(n_299), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_379), .B(n_178), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_387), .B(n_366), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_179), .B(n_194), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_384), .B(n_179), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_402), .B(n_324), .C(n_337), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_381), .A2(n_348), .B1(n_365), .B2(n_315), .Y(n_426) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_391), .A2(n_324), .B(n_337), .C(n_343), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_393), .A2(n_335), .B1(n_324), .B2(n_337), .C(n_326), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_387), .B(n_366), .Y(n_429) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_400), .A2(n_185), .B(n_193), .C(n_201), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_397), .A2(n_315), .B1(n_299), .B2(n_268), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_404), .Y(n_433) );
NOR4xp25_ASAP7_75t_SL g434 ( .A(n_394), .B(n_366), .C(n_315), .D(n_14), .Y(n_434) );
BUFx10_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
OAI31xp33_ASAP7_75t_L g436 ( .A1(n_399), .A2(n_331), .A3(n_315), .B(n_15), .Y(n_436) );
OR2x6_ASAP7_75t_L g437 ( .A(n_401), .B(n_299), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_404), .B(n_299), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_410), .B(n_395), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_409), .B(n_395), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_410), .B(n_395), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_417), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_424), .B(n_396), .Y(n_445) );
OAI31xp33_ASAP7_75t_L g446 ( .A1(n_436), .A2(n_405), .A3(n_398), .B(n_403), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_409), .B(n_405), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_424), .B(n_382), .Y(n_448) );
AOI21xp33_ASAP7_75t_SL g449 ( .A1(n_436), .A2(n_12), .B(n_13), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_415), .B(n_12), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_406), .A2(n_378), .B1(n_365), .B2(n_315), .C1(n_331), .C2(n_23), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_435), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_435), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_406), .B(n_18), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_433), .B(n_365), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_417), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_421), .A2(n_365), .B(n_206), .Y(n_457) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_420), .B(n_185), .Y(n_458) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_438), .Y(n_459) );
AND4x1_ASAP7_75t_L g460 ( .A(n_407), .B(n_19), .C(n_20), .D(n_21), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_412), .B(n_331), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_407), .B(n_365), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_439), .B(n_21), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_440), .B(n_66), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_412), .A2(n_206), .B1(n_224), .B2(n_193), .C(n_219), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_426), .B(n_331), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_425), .A2(n_220), .B1(n_209), .B2(n_171), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_440), .B(n_23), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_423), .B(n_40), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_423), .B(n_48), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_416), .B(n_438), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_423), .B(n_49), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_411), .B(n_220), .C(n_209), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_435), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_416), .B(n_50), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_408), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_435), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_432), .B(n_52), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_416), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_432), .B(n_53), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_432), .B(n_54), .Y(n_484) );
XOR2x2_ASAP7_75t_L g485 ( .A(n_426), .B(n_57), .Y(n_485) );
INVx5_ASAP7_75t_L g486 ( .A(n_418), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_408), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_463), .A2(n_411), .A3(n_431), .B1(n_430), .B2(n_224), .B3(n_219), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_442), .B(n_437), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_459), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_460), .B(n_429), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_413), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_485), .Y(n_493) );
INVx8_ASAP7_75t_L g494 ( .A(n_486), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_442), .B(n_437), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_441), .B(n_413), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_444), .Y(n_497) );
NAND2xp33_ASAP7_75t_R g498 ( .A(n_453), .B(n_434), .Y(n_498) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_453), .B(n_420), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_473), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g501 ( .A(n_477), .B(n_420), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_448), .B(n_413), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_486), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_444), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_456), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_454), .B(n_419), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_448), .B(n_413), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_473), .B(n_437), .Y(n_509) );
OAI33xp33_ASAP7_75t_L g510 ( .A1(n_463), .A2(n_431), .A3(n_204), .B1(n_201), .B2(n_434), .B3(n_427), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_476), .B(n_414), .Y(n_511) );
NAND2x1_ASAP7_75t_L g512 ( .A(n_453), .B(n_420), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_450), .B(n_422), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_485), .B(n_429), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_450), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_456), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_452), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_452), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_445), .B(n_422), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_456), .Y(n_521) );
NAND4xp25_ASAP7_75t_L g522 ( .A(n_451), .B(n_428), .C(n_421), .D(n_204), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_445), .B(n_414), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_443), .B(n_447), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_443), .B(n_437), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_469), .B(n_414), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_469), .B(n_414), .Y(n_527) );
OAI211xp5_ASAP7_75t_SL g528 ( .A1(n_451), .A2(n_437), .B(n_418), .C(n_63), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_485), .B(n_418), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_486), .B(n_418), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_453), .A2(n_59), .B1(n_61), .B2(n_64), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_460), .B(n_65), .Y(n_532) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_486), .B(n_68), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_480), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_447), .B(n_69), .Y(n_535) );
OAI33xp33_ASAP7_75t_L g536 ( .A1(n_475), .A2(n_71), .A3(n_75), .B1(n_220), .B2(n_209), .B3(n_171), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_465), .B(n_220), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_480), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_461), .B(n_171), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_455), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_519), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_515), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_500), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_493), .A2(n_462), .B1(n_467), .B2(n_475), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g546 ( .A1(n_491), .A2(n_462), .B(n_477), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_538), .B(n_482), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_540), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g549 ( .A(n_493), .B(n_486), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_516), .B(n_449), .Y(n_550) );
INVxp33_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_494), .Y(n_552) );
OAI22xp33_ASAP7_75t_L g553 ( .A1(n_529), .A2(n_449), .B1(n_486), .B2(n_478), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_488), .A2(n_486), .B1(n_458), .B2(n_478), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_520), .B(n_465), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_524), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_507), .A2(n_457), .B1(n_481), .B2(n_464), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_524), .B(n_470), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_532), .B(n_446), .C(n_458), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_499), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_528), .A2(n_464), .B1(n_457), .B2(n_483), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_503), .B(n_470), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_499), .A2(n_464), .B1(n_468), .B2(n_481), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_518), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_508), .B(n_464), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_534), .B(n_472), .Y(n_568) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_512), .A2(n_479), .B(n_487), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_502), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_502), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_501), .B(n_479), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_508), .B(n_472), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_509), .B(n_479), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_498), .B(n_466), .C(n_484), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_509), .B(n_471), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_505), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_501), .B(n_504), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_506), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_533), .A2(n_471), .B(n_483), .Y(n_580) );
NAND3xp33_ASAP7_75t_SL g581 ( .A(n_512), .B(n_474), .C(n_484), .Y(n_581) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_533), .B(n_474), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_535), .A2(n_171), .B1(n_209), .B2(n_220), .Y(n_583) );
AOI211xp5_ASAP7_75t_SL g584 ( .A1(n_504), .A2(n_171), .B(n_209), .C(n_535), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_542), .B(n_504), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_557), .B(n_523), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_553), .B(n_494), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_573), .B(n_523), .Y(n_588) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_578), .B(n_530), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_555), .Y(n_590) );
AOI221x1_ASAP7_75t_L g591 ( .A1(n_560), .A2(n_522), .B1(n_539), .B2(n_537), .C(n_521), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_544), .B(n_496), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_563), .B(n_492), .Y(n_593) );
NOR2x1p5_ASAP7_75t_L g594 ( .A(n_581), .B(n_489), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_543), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_566), .B(n_492), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_578), .A2(n_536), .B(n_510), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_541), .B(n_511), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_559), .Y(n_599) );
NOR3xp33_ASAP7_75t_SL g600 ( .A(n_553), .B(n_513), .C(n_494), .Y(n_600) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_552), .A2(n_494), .B(n_489), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_584), .A2(n_531), .B(n_495), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_541), .B(n_517), .C(n_521), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_567), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g605 ( .A(n_582), .B(n_495), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_545), .A2(n_525), .B1(n_511), .B2(n_526), .C(n_527), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_577), .B(n_526), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_565), .B(n_527), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_571), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_556), .B(n_537), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_551), .B(n_550), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_574), .B(n_577), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_575), .A2(n_554), .B(n_581), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_547), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_599), .B(n_548), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_614), .A2(n_546), .B(n_558), .C(n_572), .Y(n_618) );
OAI21xp5_ASAP7_75t_SL g619 ( .A1(n_591), .A2(n_562), .B(n_561), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_613), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_615), .B(n_576), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_607), .A2(n_558), .B1(n_568), .B2(n_572), .C(n_564), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_589), .B(n_569), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_612), .A2(n_568), .B1(n_583), .B2(n_549), .C(n_580), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_613), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_593), .B(n_596), .Y(n_626) );
AOI31xp33_ASAP7_75t_L g627 ( .A1(n_587), .A2(n_601), .A3(n_585), .B(n_597), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_605), .A2(n_594), .B1(n_602), .B2(n_609), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_591), .A2(n_600), .B(n_605), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_608), .A2(n_598), .B1(n_592), .B2(n_611), .C1(n_603), .C2(n_595), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_620), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_617), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_629), .A2(n_608), .B(n_586), .C(n_606), .Y(n_633) );
NAND2xp33_ASAP7_75t_SL g634 ( .A(n_629), .B(n_588), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_627), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_630), .B(n_588), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_621), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_619), .B(n_610), .C(n_604), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_628), .A2(n_610), .B(n_604), .Y(n_639) );
NAND2xp33_ASAP7_75t_SL g640 ( .A(n_625), .B(n_616), .Y(n_640) );
AOI31xp33_ASAP7_75t_L g641 ( .A1(n_622), .A2(n_590), .A3(n_624), .B(n_623), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_618), .B(n_590), .C(n_623), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_626), .A2(n_627), .B(n_629), .C(n_628), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_620), .Y(n_644) );
NOR3xp33_ASAP7_75t_SL g645 ( .A(n_629), .B(n_619), .C(n_614), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_619), .B(n_618), .C(n_629), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_632), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_640), .Y(n_648) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_631), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_637), .Y(n_650) );
NOR2xp33_ASAP7_75t_R g651 ( .A(n_635), .B(n_634), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_650), .B(n_646), .C(n_643), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_648), .B(n_645), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_651), .B(n_642), .C(n_638), .D(n_636), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_652), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_641), .B1(n_654), .B2(n_650), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_655), .B1(n_649), .B2(n_647), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_649), .B1(n_639), .B2(n_633), .C(n_644), .Y(n_659) );
endmodule