module fake_jpeg_25136_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_41),
.Y(n_47)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_32),
.B1(n_26),
.B2(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_38),
.B1(n_39),
.B2(n_32),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_38),
.B1(n_36),
.B2(n_18),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_31),
.B(n_21),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_32),
.B1(n_26),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_38),
.B1(n_36),
.B2(n_56),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_44),
.C(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_70),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_44),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_41),
.C(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_96),
.B1(n_36),
.B2(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_79),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_32),
.B1(n_24),
.B2(n_25),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_90),
.B(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_87),
.C(n_36),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_61),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_30),
.C(n_27),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_17),
.B1(n_34),
.B2(n_27),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_98),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_108),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_42),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_110),
.B1(n_93),
.B2(n_97),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_36),
.B1(n_39),
.B2(n_18),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_126),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_0),
.B(n_1),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_60),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_66),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_1),
.B(n_22),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_87),
.B1(n_70),
.B2(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_133),
.B1(n_134),
.B2(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_19),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_132),
.B(n_144),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_87),
.B1(n_85),
.B2(n_95),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_68),
.B1(n_97),
.B2(n_89),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_153),
.B1(n_106),
.B2(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_139),
.A2(n_150),
.B(n_22),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_147),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_68),
.B1(n_98),
.B2(n_18),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_29),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_22),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_29),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_154),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_23),
.B1(n_27),
.B2(n_67),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_22),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_19),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_143),
.B1(n_148),
.B2(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_141),
.B1(n_155),
.B2(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_165),
.A2(n_172),
.B1(n_178),
.B2(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_105),
.B(n_125),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_110),
.B(n_120),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_112),
.B1(n_115),
.B2(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_177),
.B(n_181),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_115),
.B1(n_126),
.B2(n_121),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_123),
.B(n_76),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_2),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_186),
.B(n_151),
.C(n_30),
.D(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

NOR4xp25_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_33),
.C(n_16),
.D(n_30),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_139),
.A2(n_42),
.B(n_121),
.C(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_42),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_27),
.B1(n_43),
.B2(n_37),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_144),
.B1(n_132),
.B2(n_142),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_193),
.B(n_195),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_215),
.B1(n_199),
.B2(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_219),
.B(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_179),
.C(n_173),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_203),
.C(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_34),
.B1(n_17),
.B2(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_160),
.B1(n_164),
.B2(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_159),
.B1(n_174),
.B2(n_184),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_230),
.B1(n_210),
.B2(n_197),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_217),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_169),
.B1(n_161),
.B2(n_189),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_219),
.B1(n_204),
.B2(n_202),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_207),
.A2(n_192),
.B1(n_189),
.B2(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_207),
.C(n_203),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_205),
.C(n_208),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_192),
.B(n_189),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_218),
.B(n_92),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_258),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_248),
.B1(n_259),
.B2(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_211),
.B(n_212),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_255),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_92),
.C(n_69),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_228),
.C(n_238),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_33),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_34),
.B1(n_17),
.B2(n_5),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_34),
.B1(n_17),
.B2(n_16),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_16),
.B1(n_4),
.B2(n_6),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_244),
.B1(n_229),
.B2(n_230),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_240),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_237),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_273),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_235),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_270),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_241),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_233),
.B(n_231),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_239),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_16),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_246),
.C(n_257),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_30),
.B1(n_4),
.B2(n_7),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_288),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_249),
.B(n_252),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_285),
.B(n_9),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_256),
.C(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_289),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_265),
.A2(n_262),
.B(n_256),
.Y(n_285)
);

OAI322xp33_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_263),
.A3(n_245),
.B1(n_261),
.B2(n_8),
.C1(n_9),
.C2(n_11),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_3),
.B(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_43),
.C(n_37),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_43),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_277),
.B1(n_279),
.B2(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

OAI21x1_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_3),
.B(n_7),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_8),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_283),
.C(n_284),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_287),
.B(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_284),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_11),
.B(n_13),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_286),
.A3(n_16),
.B1(n_15),
.B2(n_30),
.C1(n_43),
.C2(n_37),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_300),
.C(n_297),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_310),
.B(n_299),
.Y(n_315)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_305),
.C(n_301),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_318),
.B(n_313),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_311),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_320),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_316),
.B(n_317),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_15),
.B(n_43),
.Y(n_324)
);


endmodule