module fake_jpeg_8923_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_29),
.B1(n_26),
.B2(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_19),
.B1(n_28),
.B2(n_20),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_17),
.B1(n_22),
.B2(n_30),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_34),
.B1(n_18),
.B2(n_24),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_18),
.B1(n_34),
.B2(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_40),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_82),
.B1(n_64),
.B2(n_54),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_35),
.C(n_40),
.D(n_38),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_23),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_39),
.B1(n_36),
.B2(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_88),
.B1(n_65),
.B2(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_25),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_85),
.Y(n_109)
);

AO22x2_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_37),
.B1(n_42),
.B2(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_91),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_65),
.B1(n_27),
.B2(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_31),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_99),
.Y(n_120)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_66),
.C(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_103),
.C(n_108),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_105),
.B1(n_114),
.B2(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_118),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_57),
.C(n_45),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_4),
.B(n_5),
.Y(n_141)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_107),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_23),
.Y(n_108)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_23),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_73),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_1),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_3),
.Y(n_135)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_45),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_100),
.B1(n_95),
.B2(n_110),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_130),
.Y(n_149)
);

NOR4xp25_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_85),
.C(n_75),
.D(n_79),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_77),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_79),
.B1(n_90),
.B2(n_69),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_101),
.B1(n_105),
.B2(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_53),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_69),
.B1(n_45),
.B2(n_87),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_138),
.B1(n_106),
.B2(n_89),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_141),
.B(n_111),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_91),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_84),
.B1(n_93),
.B2(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_144),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_158),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_162),
.B1(n_165),
.B2(n_131),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_110),
.B1(n_115),
.B2(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_164),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_168),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_117),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_173),
.B(n_128),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_94),
.B(n_63),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_183),
.B1(n_197),
.B2(n_148),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_182),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_127),
.B1(n_136),
.B2(n_128),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_122),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_190),
.C(n_194),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_148),
.Y(n_211)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_191),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_122),
.C(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_193),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_144),
.C(n_142),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_173),
.B(n_167),
.C(n_158),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_123),
.B1(n_84),
.B2(n_93),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_153),
.B1(n_166),
.B2(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_151),
.CI(n_149),
.CON(n_202),
.SN(n_202)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_206),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_162),
.B1(n_123),
.B2(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_154),
.C(n_147),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_214),
.C(n_188),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_196),
.B(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_213),
.B1(n_188),
.B2(n_187),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_194),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_78),
.B1(n_63),
.B2(n_60),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_4),
.C(n_5),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_175),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_4),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_211),
.B(n_185),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_216),
.B1(n_201),
.B2(n_203),
.Y(n_235)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_228),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_214),
.C(n_198),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_223),
.B(n_227),
.C(n_8),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_200),
.C(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_242),
.C(n_243),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_181),
.C(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_246),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_202),
.C(n_207),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

AOI321xp33_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_226),
.A3(n_219),
.B1(n_229),
.B2(n_207),
.C(n_202),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_241),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_251),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_207),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_231),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_227),
.B1(n_7),
.B2(n_8),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_254),
.C(n_256),
.Y(n_258)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_253),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_264),
.C(n_250),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_263),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_9),
.B(n_10),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_264),
.C(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_6),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_269),
.A2(n_259),
.B(n_258),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_272),
.A3(n_273),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_266),
.B(n_267),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_16),
.B(n_11),
.Y(n_273)
);

AOI321xp33_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_275),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_14),
.Y(n_278)
);


endmodule