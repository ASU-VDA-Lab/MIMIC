module fake_jpeg_12944_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_17),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_2),
.B1(n_4),
.B2(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_32),
.B(n_33),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_16),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_19),
.B1(n_12),
.B2(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_9),
.B2(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_26),
.B1(n_20),
.B2(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_31),
.B(n_24),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_40),
.B1(n_35),
.B2(n_10),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_40),
.CON(n_43),
.SN(n_43)
);


endmodule