module fake_jpeg_32053_n_381 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_381);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_381;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_19),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_51),
.A2(n_18),
.B1(n_17),
.B2(n_36),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_32),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_16),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_73),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_19),
.B1(n_38),
.B2(n_32),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_104),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_32),
.B(n_31),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_18),
.B1(n_17),
.B2(n_36),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_18),
.B1(n_17),
.B2(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_30),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_107),
.B1(n_114),
.B2(n_77),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_33),
.B1(n_19),
.B2(n_37),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_113),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_42),
.A2(n_28),
.B1(n_39),
.B2(n_33),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_46),
.A2(n_21),
.B1(n_31),
.B2(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_112),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_54),
.A2(n_41),
.B1(n_23),
.B2(n_29),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_34),
.B1(n_41),
.B2(n_23),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_45),
.A2(n_41),
.B1(n_23),
.B2(n_29),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_55),
.A2(n_26),
.B1(n_34),
.B2(n_37),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_73),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_130),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_34),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_122),
.B(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_108),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_65),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_131),
.A2(n_64),
.B1(n_50),
.B2(n_43),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_142),
.B1(n_151),
.B2(n_127),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_29),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_80),
.B(n_30),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_136),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_152),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_48),
.B1(n_69),
.B2(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_80),
.B(n_63),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_149),
.Y(n_183)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_81),
.B(n_39),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_78),
.A2(n_90),
.B1(n_111),
.B2(n_39),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_20),
.B1(n_87),
.B2(n_62),
.Y(n_167)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

BUFx4f_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_58),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_105),
.B(n_13),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_11),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_78),
.B1(n_90),
.B2(n_102),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_167),
.B1(n_150),
.B2(n_132),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_133),
.B(n_140),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_165),
.A2(n_173),
.B(n_147),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_134),
.B(n_71),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_122),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_188),
.B1(n_126),
.B2(n_158),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_89),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_89),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_88),
.C(n_83),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_192),
.C(n_193),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_88),
.C(n_83),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_92),
.C(n_84),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_92),
.B1(n_60),
.B2(n_20),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_128),
.B1(n_47),
.B2(n_63),
.Y(n_212)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_149),
.B1(n_153),
.B2(n_139),
.Y(n_200)
);

HB1xp67_ASAP7_75t_SL g258 ( 
.A(n_200),
.Y(n_258)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_119),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_212),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_117),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_124),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_126),
.C(n_152),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_213),
.C(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_137),
.B1(n_118),
.B2(n_144),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_216),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_162),
.B(n_177),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_156),
.B1(n_157),
.B2(n_66),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_164),
.A2(n_10),
.B1(n_58),
.B2(n_3),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_146),
.C(n_145),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_165),
.A2(n_40),
.B(n_146),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_188),
.B(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_176),
.B(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_176),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_178),
.B1(n_163),
.B2(n_175),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_40),
.B1(n_146),
.B2(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_230),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_40),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_236),
.B(n_222),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_189),
.B(n_193),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_255),
.B1(n_218),
.B2(n_212),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_192),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_251),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_249),
.A2(n_252),
.B(n_259),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_162),
.C(n_181),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_162),
.B(n_173),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_240),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_167),
.B1(n_175),
.B2(n_171),
.Y(n_255)
);

XOR2x1_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_168),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_210),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_262),
.A2(n_276),
.B1(n_279),
.B2(n_245),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_266),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_196),
.B1(n_199),
.B2(n_203),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_278),
.B(n_231),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_223),
.B1(n_224),
.B2(n_216),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_201),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_213),
.B1(n_221),
.B2(n_196),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_241),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_283),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_273),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_227),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_220),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_214),
.B1(n_205),
.B2(n_229),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_168),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_197),
.B1(n_179),
.B2(n_172),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_194),
.B1(n_172),
.B2(n_179),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_190),
.B1(n_166),
.B2(n_40),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_1),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_235),
.A2(n_190),
.B1(n_154),
.B2(n_5),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_285),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_190),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_1),
.C(n_4),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_242),
.B(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_6),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_294),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_295),
.B1(n_298),
.B2(n_250),
.Y(n_321)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_250),
.B1(n_252),
.B2(n_236),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_263),
.C(n_239),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_305),
.C(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_251),
.C(n_249),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_250),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_265),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_285),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_311),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_313),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_242),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_264),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_323),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_264),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_318),
.C(n_322),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_268),
.C(n_238),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_291),
.A2(n_262),
.B1(n_278),
.B2(n_276),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_320),
.A2(n_304),
.B1(n_247),
.B2(n_293),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_279),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_238),
.C(n_281),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_306),
.B(n_291),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_298),
.B(n_259),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_289),
.B(n_296),
.Y(n_327)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_SL g326 ( 
.A(n_310),
.B(n_287),
.C(n_294),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_331),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_337),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_296),
.B(n_300),
.Y(n_328)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_259),
.B(n_300),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_330),
.A2(n_280),
.B(n_255),
.Y(n_351)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_288),
.C(n_299),
.Y(n_331)
);

AOI221xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_303),
.B1(n_283),
.B2(n_304),
.C(n_299),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_334),
.A2(n_335),
.B(n_340),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_322),
.B(n_245),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_318),
.C(n_323),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_341),
.B(n_342),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_313),
.C(n_317),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_315),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_344),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_314),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_309),
.C(n_246),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_350),
.C(n_333),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_237),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_233),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_246),
.C(n_257),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_351),
.B(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_348),
.B(n_342),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_356),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_345),
.B(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_341),
.B(n_244),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_359),
.B(n_362),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_348),
.A2(n_332),
.B1(n_334),
.B2(n_244),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_360),
.A2(n_350),
.B(n_243),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_243),
.C(n_154),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_233),
.B1(n_282),
.B2(n_257),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_367),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_355),
.A2(n_154),
.B(n_7),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_7),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_354),
.C(n_353),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_371),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_365),
.B(n_357),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_373),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_SL g374 ( 
.A(n_369),
.B(n_360),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_375),
.A2(n_364),
.B(n_370),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_377),
.Y(n_378)
);

A2O1A1O1Ixp25_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_374),
.B(n_363),
.C(n_372),
.D(n_367),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_372),
.C(n_376),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_7),
.Y(n_381)
);


endmodule