module real_aes_884_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_713;
wire n_728;
wire n_598;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_481;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g245 ( .A(n_0), .B(n_152), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_2), .B(n_141), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_3), .B(n_150), .Y(n_502) );
INVx1_ASAP7_75t_L g140 ( .A(n_4), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_5), .B(n_141), .Y(n_198) );
NAND2xp33_ASAP7_75t_SL g191 ( .A(n_6), .B(n_147), .Y(n_191) );
INVx1_ASAP7_75t_L g171 ( .A(n_7), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
AND2x2_ASAP7_75t_L g196 ( .A(n_9), .B(n_131), .Y(n_196) );
AND2x2_ASAP7_75t_L g495 ( .A(n_10), .B(n_188), .Y(n_495) );
AND2x2_ASAP7_75t_L g504 ( .A(n_11), .B(n_163), .Y(n_504) );
INVx2_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_13), .B(n_150), .Y(n_557) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_14), .Y(n_114) );
AOI221x1_ASAP7_75t_L g185 ( .A1(n_15), .A2(n_135), .B1(n_186), .B2(n_188), .C(n_190), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_16), .B(n_141), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_17), .B(n_141), .Y(n_542) );
INVx1_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_19), .A2(n_93), .B1(n_141), .B2(n_173), .Y(n_483) );
AOI221xp5_ASAP7_75t_SL g134 ( .A1(n_20), .A2(n_35), .B1(n_135), .B2(n_141), .C(n_148), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_21), .A2(n_135), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_22), .B(n_152), .Y(n_201) );
OR2x2_ASAP7_75t_L g133 ( .A(n_23), .B(n_92), .Y(n_133) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_23), .A2(n_92), .B(n_132), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_24), .B(n_150), .Y(n_162) );
INVxp67_ASAP7_75t_L g184 ( .A(n_25), .Y(n_184) );
AND2x2_ASAP7_75t_L g234 ( .A(n_26), .B(n_130), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_27), .A2(n_135), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_28), .A2(n_188), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_29), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_30), .A2(n_135), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_31), .B(n_150), .Y(n_537) );
AND2x2_ASAP7_75t_L g136 ( .A(n_32), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g147 ( .A(n_32), .B(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g180 ( .A(n_32), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g111 ( .A(n_33), .B(n_112), .C(n_114), .Y(n_111) );
OR2x6_ASAP7_75t_L g455 ( .A(n_33), .B(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_34), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_34), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_36), .B(n_141), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_37), .A2(n_85), .B1(n_135), .B2(n_178), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_38), .B(n_150), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_39), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_40), .B(n_141), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_41), .B(n_152), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_42), .A2(n_135), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_43), .A2(n_75), .B1(n_759), .B2(n_760), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_43), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_44), .A2(n_754), .B1(n_764), .B2(n_766), .Y(n_763) );
AND2x2_ASAP7_75t_L g248 ( .A(n_45), .B(n_130), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_46), .B(n_152), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_47), .B(n_130), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_48), .B(n_141), .Y(n_554) );
INVx1_ASAP7_75t_L g139 ( .A(n_49), .Y(n_139) );
INVx1_ASAP7_75t_L g144 ( .A(n_49), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_50), .B(n_150), .Y(n_493) );
OAI22x1_ASAP7_75t_R g442 ( .A1(n_51), .A2(n_443), .B1(n_446), .B2(n_447), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_51), .Y(n_446) );
AOI22xp5_ASAP7_75t_SL g754 ( .A1(n_52), .A2(n_755), .B1(n_761), .B2(n_762), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_52), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_53), .Y(n_771) );
AND2x2_ASAP7_75t_L g523 ( .A(n_54), .B(n_130), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_55), .B(n_141), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_56), .B(n_152), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_57), .B(n_152), .Y(n_536) );
AND2x2_ASAP7_75t_L g212 ( .A(n_58), .B(n_130), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_59), .B(n_141), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_60), .B(n_150), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_61), .B(n_141), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_62), .A2(n_135), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_63), .B(n_131), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_64), .B(n_152), .Y(n_209) );
AND2x2_ASAP7_75t_L g548 ( .A(n_65), .B(n_131), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_66), .A2(n_135), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_67), .B(n_150), .Y(n_202) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_68), .B(n_163), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_69), .B(n_152), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_70), .A2(n_73), .B1(n_444), .B2(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_70), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_71), .B(n_152), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_72), .A2(n_95), .B1(n_135), .B2(n_178), .Y(n_484) );
INVx1_ASAP7_75t_L g445 ( .A(n_73), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_74), .B(n_150), .Y(n_545) );
INVx1_ASAP7_75t_L g760 ( .A(n_75), .Y(n_760) );
INVx1_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_76), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_77), .B(n_152), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_78), .A2(n_135), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_79), .A2(n_135), .B(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_80), .A2(n_135), .B(n_556), .Y(n_555) );
XNOR2x1_ASAP7_75t_SL g122 ( .A(n_81), .B(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g539 ( .A(n_81), .B(n_131), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_82), .B(n_130), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_83), .B(n_141), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_84), .A2(n_87), .B1(n_141), .B2(n_173), .Y(n_217) );
INVx1_ASAP7_75t_L g109 ( .A(n_86), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_88), .B(n_152), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_89), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g516 ( .A(n_90), .B(n_163), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_91), .A2(n_135), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_94), .B(n_150), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_96), .A2(n_135), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_97), .B(n_150), .Y(n_514) );
INVxp67_ASAP7_75t_L g187 ( .A(n_98), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_99), .B(n_141), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_100), .B(n_150), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_101), .A2(n_135), .B(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g547 ( .A(n_102), .Y(n_547) );
BUFx2_ASAP7_75t_L g120 ( .A(n_103), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_103), .B(n_457), .Y(n_460) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_115), .B(n_770), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g772 ( .A(n_106), .Y(n_772) );
INVx3_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_109), .B(n_110), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_114), .B(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_SL g466 ( .A(n_114), .B(n_455), .Y(n_466) );
OR2x6_ASAP7_75t_SL g469 ( .A(n_114), .B(n_454), .Y(n_469) );
OR2x2_ASAP7_75t_L g769 ( .A(n_114), .B(n_455), .Y(n_769) );
OA22x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B1(n_460), .B2(n_461), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_449), .B(n_457), .Y(n_121) );
OAI22x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_441), .B1(n_442), .B2(n_448), .Y(n_123) );
INVx2_ASAP7_75t_L g448 ( .A(n_124), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_124), .A2(n_467), .B1(n_471), .B2(n_765), .Y(n_764) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_354), .Y(n_124) );
NAND3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_264), .C(n_304), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_166), .B(n_193), .C(n_220), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_127), .B(n_269), .Y(n_303) );
NOR2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_155), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g239 ( .A(n_129), .Y(n_239) );
INVx2_ASAP7_75t_L g255 ( .A(n_129), .Y(n_255) );
OR2x2_ASAP7_75t_L g267 ( .A(n_129), .B(n_156), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_129), .B(n_240), .Y(n_281) );
INVx1_ASAP7_75t_L g309 ( .A(n_129), .Y(n_309) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_129), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_129), .B(n_156), .Y(n_415) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_130), .Y(n_211) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_130), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_130), .A2(n_511), .B(n_512), .Y(n_510) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x4_ASAP7_75t_L g172 ( .A(n_132), .B(n_133), .Y(n_172) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
BUFx3_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
AND2x6_ASAP7_75t_L g152 ( .A(n_137), .B(n_143), .Y(n_152) );
INVx2_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
AND2x4_ASAP7_75t_L g178 ( .A(n_138), .B(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g150 ( .A(n_139), .B(n_145), .Y(n_150) );
INVx2_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
INVx1_ASAP7_75t_L g192 ( .A(n_142), .Y(n_192) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx5_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B(n_153), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_152), .B(n_547), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_153), .A2(n_161), .B(n_162), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_153), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_153), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_153), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_153), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_153), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_153), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_153), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_153), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_153), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_153), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_153), .A2(n_557), .B(n_558), .Y(n_556) );
OR2x2_ASAP7_75t_L g236 ( .A(n_155), .B(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_155), .Y(n_371) );
AND2x2_ASAP7_75t_L g376 ( .A(n_155), .B(n_238), .Y(n_376) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g166 ( .A(n_156), .B(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g235 ( .A(n_156), .B(n_168), .Y(n_235) );
OR2x2_ASAP7_75t_L g254 ( .A(n_156), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g283 ( .A(n_156), .Y(n_283) );
AND2x4_ASAP7_75t_SL g322 ( .A(n_156), .B(n_168), .Y(n_322) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_156), .Y(n_326) );
OR2x2_ASAP7_75t_L g343 ( .A(n_156), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g353 ( .A(n_156), .B(n_260), .Y(n_353) );
INVx1_ASAP7_75t_L g382 ( .A(n_156), .Y(n_382) );
OR2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_165), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_163), .Y(n_157) );
INVx2_ASAP7_75t_SL g215 ( .A(n_163), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_163), .A2(n_542), .B(n_543), .Y(n_541) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g189 ( .A(n_164), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_166), .B(n_311), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_167), .B(n_240), .Y(n_257) );
AND2x2_ASAP7_75t_L g269 ( .A(n_167), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g287 ( .A(n_167), .B(n_254), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_167), .B(n_308), .Y(n_307) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g260 ( .A(n_168), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g282 ( .A(n_168), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g317 ( .A(n_168), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_168), .B(n_240), .Y(n_341) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_185), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B1(n_178), .B2(n_183), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_172), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_172), .B(n_187), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g190 ( .A(n_172), .B(n_191), .C(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_172), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_172), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_172), .A2(n_554), .B(n_555), .Y(n_553) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_177), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g532 ( .A(n_188), .Y(n_532) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_189), .A2(n_242), .B(n_248), .Y(n_241) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_189), .A2(n_489), .B(n_495), .Y(n_488) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_194), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g290 ( .A(n_194), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_194), .B(n_204), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_194), .B(n_311), .C(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g358 ( .A(n_194), .B(n_263), .Y(n_358) );
INVx5_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g225 ( .A(n_195), .B(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_SL g262 ( .A(n_195), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g278 ( .A(n_195), .Y(n_278) );
OR2x2_ASAP7_75t_L g301 ( .A(n_195), .B(n_291), .Y(n_301) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_195), .Y(n_318) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_195), .B(n_224), .Y(n_336) );
AND2x4_ASAP7_75t_L g351 ( .A(n_195), .B(n_227), .Y(n_351) );
AND2x2_ASAP7_75t_L g365 ( .A(n_195), .B(n_204), .Y(n_365) );
OR2x2_ASAP7_75t_L g386 ( .A(n_195), .B(n_213), .Y(n_386) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_L g440 ( .A(n_203), .B(n_318), .Y(n_440) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
AND2x4_ASAP7_75t_L g263 ( .A(n_204), .B(n_226), .Y(n_263) );
INVx2_ASAP7_75t_L g274 ( .A(n_204), .Y(n_274) );
AND2x2_ASAP7_75t_L g279 ( .A(n_204), .B(n_224), .Y(n_279) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_204), .Y(n_312) );
OR2x2_ASAP7_75t_L g335 ( .A(n_204), .B(n_227), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_204), .B(n_227), .Y(n_338) );
INVx1_ASAP7_75t_L g347 ( .A(n_204), .Y(n_347) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_211), .B(n_212), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_211), .A2(n_228), .B(n_234), .Y(n_227) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_211), .A2(n_228), .B(n_234), .Y(n_291) );
AOI21x1_ASAP7_75t_L g497 ( .A1(n_211), .A2(n_498), .B(n_504), .Y(n_497) );
AND2x2_ASAP7_75t_L g250 ( .A(n_213), .B(n_227), .Y(n_250) );
BUFx2_ASAP7_75t_L g299 ( .A(n_213), .Y(n_299) );
AND2x2_ASAP7_75t_L g394 ( .A(n_213), .B(n_274), .Y(n_394) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
AOI21x1_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_219), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_235), .B1(n_236), .B2(n_249), .C(n_251), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
NOR2x1_ASAP7_75t_L g296 ( .A(n_223), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_223), .B(n_290), .Y(n_330) );
OR2x2_ASAP7_75t_L g342 ( .A(n_223), .B(n_338), .Y(n_342) );
OR2x2_ASAP7_75t_L g345 ( .A(n_223), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g434 ( .A(n_223), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_L g273 ( .A(n_224), .B(n_274), .Y(n_273) );
OA33x2_ASAP7_75t_L g306 ( .A1(n_224), .A2(n_267), .A3(n_307), .B1(n_310), .B2(n_313), .B3(n_316), .Y(n_306) );
OR2x2_ASAP7_75t_L g337 ( .A(n_224), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g361 ( .A(n_224), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g369 ( .A(n_224), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g389 ( .A(n_224), .B(n_263), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_224), .B(n_278), .Y(n_427) );
INVx2_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
AOI322xp5_ASAP7_75t_L g367 ( .A1(n_225), .A2(n_280), .A3(n_368), .B1(n_371), .B2(n_372), .C1(n_374), .C2(n_376), .Y(n_367) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_227), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
OR2x2_ASAP7_75t_L g349 ( .A(n_235), .B(n_328), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_235), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g422 ( .A(n_235), .Y(n_422) );
INVx1_ASAP7_75t_SL g288 ( .A(n_236), .Y(n_288) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g321 ( .A(n_238), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g261 ( .A(n_240), .Y(n_261) );
INVx1_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
INVx1_ASAP7_75t_L g311 ( .A(n_240), .Y(n_311) );
OR2x2_ASAP7_75t_L g328 ( .A(n_240), .B(n_255), .Y(n_328) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_240), .Y(n_403) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_250), .B(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_258), .B(n_262), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_252), .A2(n_326), .B(n_327), .C(n_329), .Y(n_325) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g390 ( .A(n_254), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_255), .Y(n_259) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g414 ( .A(n_257), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_260), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g391 ( .A(n_260), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_260), .B(n_382), .Y(n_399) );
INVx3_ASAP7_75t_SL g324 ( .A(n_263), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_271), .B1(n_275), .B2(n_280), .C(n_284), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_270), .Y(n_315) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_273), .A2(n_300), .B(n_372), .Y(n_378) );
AND2x2_ASAP7_75t_L g404 ( .A(n_273), .B(n_351), .Y(n_404) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_274), .Y(n_292) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g413 ( .A(n_278), .B(n_335), .Y(n_413) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g362 ( .A(n_281), .Y(n_362) );
OAI21xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B(n_293), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx2_ASAP7_75t_L g435 ( .A(n_290), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_291), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g364 ( .A(n_291), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_292), .B(n_314), .Y(n_313) );
OAI31xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .A3(n_298), .B(n_302), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_297), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g375 ( .A(n_299), .B(n_301), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_299), .B(n_351), .Y(n_430) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR5xp2_ASAP7_75t_L g304 ( .A(n_305), .B(n_319), .C(n_331), .D(n_340), .E(n_348), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_309), .B(n_311), .Y(n_344) );
INVx1_ASAP7_75t_L g384 ( .A(n_309), .Y(n_384) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_309), .Y(n_421) );
INVx1_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OAI321xp33_ASAP7_75t_L g356 ( .A1(n_317), .A2(n_357), .A3(n_359), .B1(n_363), .B2(n_366), .C(n_367), .Y(n_356) );
INVx1_ASAP7_75t_L g410 ( .A(n_318), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B(n_325), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_321), .A2(n_394), .B1(n_401), .B2(n_404), .Y(n_400) );
AND2x2_ASAP7_75t_L g429 ( .A(n_322), .B(n_403), .Y(n_429) );
INVx1_ASAP7_75t_L g339 ( .A(n_327), .Y(n_339) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_337), .B(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_338), .A2(n_349), .B1(n_350), .B2(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g411 ( .A(n_338), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_343), .B2(n_345), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_347), .B(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_349), .A2(n_426), .B1(n_428), .B2(n_430), .C(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_349), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_350), .A2(n_407), .B1(n_414), .B2(n_416), .C(n_417), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_352), .A2(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_405), .Y(n_354) );
NOR3xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_377), .C(n_395), .Y(n_355) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_358), .Y(n_424) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_368), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g416 ( .A(n_376), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_385), .B(n_387), .Y(n_379) );
INVxp67_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g392 ( .A(n_383), .Y(n_392) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B1(n_392), .B2(n_393), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_400), .Y(n_395) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_425), .C(n_436), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_412), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_423), .B(n_424), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_429), .A2(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g447 ( .A(n_443), .Y(n_447) );
OA22x2_ASAP7_75t_L g462 ( .A1(n_448), .A2(n_463), .B1(n_467), .B2(n_470), .Y(n_462) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g459 ( .A(n_453), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
OAI21xp33_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_754), .B(n_763), .Y(n_461) );
CKINVDCx6p67_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_SL g765 ( .A(n_464), .Y(n_765) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
CKINVDCx11_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_691), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_607), .C(n_644), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_575), .C(n_590), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_520), .B1(n_549), .B2(n_561), .C(n_562), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_477), .B(n_505), .Y(n_476) );
OAI22xp33_ASAP7_75t_SL g635 ( .A1(n_477), .A2(n_599), .B1(n_636), .B2(n_639), .Y(n_635) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
OAI21xp33_ASAP7_75t_SL g645 ( .A1(n_478), .A2(n_646), .B(n_652), .Y(n_645) );
OR2x2_ASAP7_75t_L g674 ( .A(n_478), .B(n_507), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_478), .B(n_594), .Y(n_675) );
INVx2_ASAP7_75t_L g706 ( .A(n_478), .Y(n_706) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_479), .B(n_566), .Y(n_687) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g561 ( .A(n_480), .B(n_488), .Y(n_561) );
BUFx3_ASAP7_75t_L g587 ( .A(n_480), .Y(n_587) );
AND2x2_ASAP7_75t_L g723 ( .A(n_480), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g746 ( .A(n_480), .B(n_508), .Y(n_746) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x4_ASAP7_75t_L g519 ( .A(n_481), .B(n_482), .Y(n_519) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_486), .B(n_508), .Y(n_666) );
INVx1_ASAP7_75t_L g703 ( .A(n_486), .Y(n_703) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
AND2x2_ASAP7_75t_L g518 ( .A(n_487), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g724 ( .A(n_487), .Y(n_724) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g567 ( .A(n_488), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_488), .B(n_496), .Y(n_568) );
AND2x2_ASAP7_75t_L g589 ( .A(n_488), .B(n_509), .Y(n_589) );
AND2x2_ASAP7_75t_L g671 ( .A(n_488), .B(n_497), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
AND2x4_ASAP7_75t_SL g564 ( .A(n_496), .B(n_509), .Y(n_564) );
INVx1_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
INVx2_ASAP7_75t_L g603 ( .A(n_496), .Y(n_603) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_496), .Y(n_627) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_497), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_518), .Y(n_505) );
AND2x2_ASAP7_75t_L g742 ( .A(n_506), .B(n_605), .Y(n_742) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_508), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g653 ( .A(n_508), .B(n_568), .Y(n_653) );
AND2x2_ASAP7_75t_L g670 ( .A(n_508), .B(n_671), .Y(n_670) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_L g594 ( .A(n_509), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g610 ( .A(n_509), .Y(n_610) );
AND2x2_ASAP7_75t_L g654 ( .A(n_509), .B(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g661 ( .A(n_509), .B(n_662), .Y(n_661) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_509), .B(n_567), .Y(n_676) );
BUFx2_ASAP7_75t_L g686 ( .A(n_509), .Y(n_686) );
AND2x2_ASAP7_75t_L g711 ( .A(n_509), .B(n_671), .Y(n_711) );
AND2x2_ASAP7_75t_L g732 ( .A(n_509), .B(n_733), .Y(n_732) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g663 ( .A(n_517), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_518), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g693 ( .A(n_518), .B(n_564), .Y(n_693) );
INVx3_ASAP7_75t_L g600 ( .A(n_519), .Y(n_600) );
AND2x2_ASAP7_75t_L g733 ( .A(n_519), .B(n_655), .Y(n_733) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_521), .A2(n_563), .B1(n_568), .B2(n_569), .Y(n_562) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_530), .Y(n_521) );
INVx4_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
INVx2_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
NAND2x1_ASAP7_75t_L g623 ( .A(n_522), .B(n_540), .Y(n_623) );
OR2x2_ASAP7_75t_L g638 ( .A(n_522), .B(n_573), .Y(n_638) );
OR2x2_ASAP7_75t_SL g665 ( .A(n_522), .B(n_637), .Y(n_665) );
AND2x2_ASAP7_75t_L g678 ( .A(n_522), .B(n_552), .Y(n_678) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_522), .Y(n_699) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g578 ( .A(n_530), .Y(n_578) );
AND2x2_ASAP7_75t_L g710 ( .A(n_530), .B(n_684), .Y(n_710) );
NOR2x1_ASAP7_75t_SL g530 ( .A(n_531), .B(n_540), .Y(n_530) );
AND2x2_ASAP7_75t_L g551 ( .A(n_531), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g727 ( .A(n_531), .B(n_650), .Y(n_727) );
AO21x1_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_533), .B(n_539), .Y(n_531) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_532), .A2(n_533), .B(n_539), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
OR2x2_ASAP7_75t_L g559 ( .A(n_540), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g570 ( .A(n_540), .B(n_560), .Y(n_570) );
AND2x2_ASAP7_75t_L g616 ( .A(n_540), .B(n_573), .Y(n_616) );
OR2x2_ASAP7_75t_L g637 ( .A(n_540), .B(n_552), .Y(n_637) );
INVx2_ASAP7_75t_SL g643 ( .A(n_540), .Y(n_643) );
AND2x2_ASAP7_75t_L g649 ( .A(n_540), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g659 ( .A(n_540), .B(n_642), .Y(n_659) );
BUFx2_ASAP7_75t_L g681 ( .A(n_540), .Y(n_681) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_548), .Y(n_540) );
INVx2_ASAP7_75t_L g728 ( .A(n_549), .Y(n_728) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_559), .Y(n_549) );
OR2x2_ASAP7_75t_L g753 ( .A(n_550), .B(n_597), .Y(n_753) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_551), .B(n_560), .Y(n_619) );
AND2x2_ASAP7_75t_L g690 ( .A(n_551), .B(n_570), .Y(n_690) );
INVx1_ASAP7_75t_L g572 ( .A(n_552), .Y(n_572) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_552), .Y(n_581) );
INVx1_ASAP7_75t_L g614 ( .A(n_552), .Y(n_614) );
INVx2_ASAP7_75t_L g650 ( .A(n_552), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g580 ( .A(n_560), .B(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g640 ( .A(n_560), .Y(n_640) );
INVx2_ASAP7_75t_SL g716 ( .A(n_561), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_563), .A2(n_618), .B1(n_620), .B2(n_624), .Y(n_617) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g744 ( .A(n_564), .B(n_600), .Y(n_744) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_566), .B(n_610), .Y(n_689) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g655 ( .A(n_567), .B(n_603), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_568), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_569), .A2(n_713), .B1(n_717), .B2(n_719), .C(n_721), .Y(n_712) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g582 ( .A(n_570), .B(n_583), .Y(n_582) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_570), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_570), .B(n_613), .Y(n_668) );
INVx1_ASAP7_75t_SL g664 ( .A(n_571), .Y(n_664) );
AOI221xp5_ASAP7_75t_SL g692 ( .A1(n_571), .A2(n_582), .B1(n_693), .B2(n_694), .C(n_697), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g725 ( .A1(n_571), .A2(n_643), .A3(n_670), .B1(n_726), .B2(n_728), .C1(n_729), .C2(n_732), .Y(n_725) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx2_ASAP7_75t_L g592 ( .A(n_572), .Y(n_592) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_573), .Y(n_584) );
INVx2_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
AND2x2_ASAP7_75t_L g683 ( .A(n_573), .B(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OA21x2_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_582), .B(n_585), .Y(n_575) );
AOI211xp5_ASAP7_75t_L g745 ( .A1(n_576), .A2(n_746), .B(n_747), .C(n_751), .Y(n_745) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OR2x2_ASAP7_75t_L g634 ( .A(n_578), .B(n_596), .Y(n_634) );
OR2x2_ASAP7_75t_L g718 ( .A(n_578), .B(n_613), .Y(n_718) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g658 ( .A(n_580), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g736 ( .A(n_583), .Y(n_736) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g622 ( .A(n_584), .Y(n_622) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g591 ( .A(n_587), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g626 ( .A(n_589), .B(n_627), .Y(n_626) );
OAI322xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .A3(n_596), .B1(n_598), .B2(n_599), .C1(n_604), .C2(n_606), .Y(n_590) );
INVx1_ASAP7_75t_L g632 ( .A(n_591), .Y(n_632) );
OR2x2_ASAP7_75t_L g604 ( .A(n_593), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_593), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g615 ( .A(n_597), .B(n_616), .Y(n_615) );
OAI32xp33_ASAP7_75t_L g660 ( .A1(n_597), .A2(n_661), .A3(n_664), .B1(n_665), .B2(n_666), .Y(n_660) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx2_ASAP7_75t_L g605 ( .A(n_600), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_600), .B(n_663), .Y(n_662) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_600), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g726 ( .A(n_600), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g647 ( .A(n_601), .Y(n_647) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_605), .B(n_671), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_628), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B(n_617), .Y(n_608) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_SL g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g677 ( .A(n_616), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_619), .A2(n_639), .B1(n_741), .B2(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_621), .A2(n_668), .B(n_669), .C(n_672), .Y(n_667) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx3_ASAP7_75t_L g749 ( .A(n_623), .Y(n_749) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g630 ( .A(n_627), .Y(n_630) );
AO21x1_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_635), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g695 ( .A(n_630), .Y(n_695) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_636), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g651 ( .A(n_638), .Y(n_651) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g708 ( .A(n_641), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_667), .C(n_679), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_648), .A2(n_710), .B(n_711), .Y(n_709) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g684 ( .A(n_650), .Y(n_684) );
O2A1O1Ixp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_662), .Y(n_752) );
INVx2_ASAP7_75t_L g737 ( .A(n_665), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g751 ( .A1(n_666), .A2(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g731 ( .A(n_671), .Y(n_731) );
OAI31xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .A3(n_676), .B(n_677), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g750 ( .A(n_678), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_685), .B(n_688), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
BUFx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g700 ( .A(n_683), .Y(n_700) );
AOI21xp33_ASAP7_75t_SL g747 ( .A1(n_685), .A2(n_748), .B(n_750), .Y(n_747) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_L g715 ( .A(n_686), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_686), .B(n_706), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_686), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g696 ( .A(n_687), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NAND5xp2_ASAP7_75t_L g691 ( .A(n_692), .B(n_712), .C(n_725), .D(n_734), .E(n_745), .Y(n_691) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B1(n_704), .B2(n_707), .C(n_709), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_738), .B(n_740), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g762 ( .A(n_755), .Y(n_762) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
endmodule