module fake_jpeg_16528_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_25),
.Y(n_53)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_17),
.B1(n_28),
.B2(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_57),
.Y(n_86)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_54),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_30),
.B(n_21),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_73),
.B1(n_99),
.B2(n_101),
.Y(n_109)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_91),
.B1(n_29),
.B2(n_32),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_81),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_37),
.C(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_36),
.B1(n_38),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_55),
.B1(n_60),
.B2(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_19),
.B1(n_26),
.B2(n_22),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_38),
.B1(n_19),
.B2(n_42),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_92),
.A2(n_34),
.B1(n_18),
.B2(n_27),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_97),
.Y(n_119)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_38),
.B1(n_41),
.B2(n_36),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_41),
.B1(n_42),
.B2(n_21),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_55),
.B1(n_31),
.B2(n_51),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_48),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_98),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_129),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_27),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_112),
.B(n_81),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_86),
.B(n_67),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_116),
.B(n_108),
.Y(n_139)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_30),
.B(n_31),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_83),
.A2(n_41),
.B1(n_20),
.B2(n_18),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_20),
.B1(n_10),
.B2(n_15),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_20),
.B1(n_18),
.B2(n_34),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_72),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_69),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_137),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_120),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_99),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_141),
.C(n_157),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_94),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_78),
.B(n_99),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_34),
.B(n_18),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_144),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_118),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_89),
.C(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_76),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_76),
.B1(n_96),
.B2(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_74),
.B1(n_110),
.B2(n_105),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_80),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_104),
.C(n_125),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_34),
.B(n_18),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_160),
.B(n_0),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_0),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_161),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_157),
.A2(n_122),
.B1(n_117),
.B2(n_128),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_164),
.B1(n_174),
.B2(n_147),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_117),
.B1(n_75),
.B2(n_125),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_146),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_134),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_118),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_191),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_169),
.A2(n_177),
.B(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_117),
.B1(n_110),
.B2(n_131),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_105),
.B1(n_121),
.B2(n_74),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_11),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_183),
.A2(n_184),
.B(n_186),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_27),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_137),
.B(n_105),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_27),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_88),
.C(n_14),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_194),
.B(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_160),
.B1(n_154),
.B2(n_162),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_12),
.B(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_197),
.B(n_167),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_138),
.B(n_139),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_207),
.B(n_222),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_211),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_214),
.C(n_225),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_174),
.B1(n_164),
.B2(n_184),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_159),
.B(n_154),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_165),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_177),
.B1(n_183),
.B2(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_152),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_182),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_146),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_166),
.A2(n_160),
.B(n_132),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_161),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_231),
.C(n_234),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_201),
.B1(n_216),
.B2(n_208),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_180),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_180),
.C(n_191),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_186),
.C(n_163),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_237),
.C(n_198),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_179),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_244),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_197),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_199),
.A2(n_196),
.B1(n_173),
.B2(n_181),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_173),
.B1(n_216),
.B2(n_215),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_246),
.B(n_167),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_240),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_268),
.B1(n_269),
.B2(n_242),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_265),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_258),
.A2(n_245),
.B1(n_236),
.B2(n_247),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_219),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_239),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_209),
.C(n_207),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_222),
.C(n_215),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_217),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_195),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_217),
.B(n_205),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_212),
.B1(n_205),
.B2(n_200),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_234),
.C(n_235),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_231),
.C(n_237),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_226),
.C(n_239),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_244),
.CI(n_229),
.CON(n_275),
.SN(n_275)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_192),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_243),
.C(n_232),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_285),
.C(n_267),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_250),
.B1(n_256),
.B2(n_252),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_266),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_232),
.B1(n_229),
.B2(n_200),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_256),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_169),
.C(n_175),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_282),
.A2(n_268),
.B(n_252),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_295),
.B(n_280),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_291),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_275),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_297),
.C(n_299),
.Y(n_307)
);

NAND2x1_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_250),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_193),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_276),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_3),
.C(n_4),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_8),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_274),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_310),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_270),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_270),
.B(n_272),
.Y(n_309)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_290),
.B(n_6),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_273),
.B(n_10),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_297),
.A3(n_287),
.B1(n_290),
.B2(n_11),
.C1(n_12),
.C2(n_7),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_317),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_306),
.C(n_313),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_5),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_5),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_5),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_305),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_319),
.B(n_325),
.C(n_314),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_320),
.B(n_312),
.Y(n_327)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_6),
.A3(n_7),
.B1(n_300),
.B2(n_324),
.C(n_319),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);


endmodule