module fake_jpeg_30401_n_35 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_35);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_6),
.C(n_10),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_2),
.B(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_2),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.C(n_13),
.Y(n_30)
);

OAI322xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_14),
.A3(n_4),
.B1(n_5),
.B2(n_8),
.C1(n_9),
.C2(n_12),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_13),
.Y(n_32)
);

NAND4xp25_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_17),
.C(n_3),
.D(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);


endmodule