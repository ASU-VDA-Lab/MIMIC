module fake_ibex_2059_n_4039 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4039);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4039;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_3458;
wire n_3653;
wire n_2955;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_2979;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_3323;
wire n_2820;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3839;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3949;
wire n_3507;
wire n_3881;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3766;
wire n_2822;
wire n_4014;
wire n_3022;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_3030;
wire n_2906;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_3199;
wire n_1616;
wire n_2723;
wire n_3808;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3634;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3448;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_3614;
wire n_2339;
wire n_2888;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_3331;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_3578;
wire n_954;
wire n_2971;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3948;
wire n_3719;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_3398;
wire n_3718;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2923;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_3284;
wire n_2524;
wire n_3835;
wire n_1437;
wire n_2875;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_3902;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_961;
wire n_991;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3269;
wire n_3609;
wire n_3029;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3376;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2576;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_2658;
wire n_3236;
wire n_3576;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3343;
wire n_3163;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_980;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_3124;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2961;
wire n_2770;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3635;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_3180;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g846 ( 
.A(n_413),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_482),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_207),
.Y(n_848)
);

BUFx5_ASAP7_75t_L g849 ( 
.A(n_242),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_632),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_326),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_765),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_547),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_46),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_47),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_454),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_226),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_438),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_824),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_809),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_165),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_560),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_240),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_296),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_551),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_448),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_387),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_637),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_395),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_260),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_28),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_303),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_645),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_556),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_254),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_418),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_655),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_739),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_781),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_29),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_403),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_413),
.Y(n_882)
);

BUFx10_ASAP7_75t_L g883 ( 
.A(n_173),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_616),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_290),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_278),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_686),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_231),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_672),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_580),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_8),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_378),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_84),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_580),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_324),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_762),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_298),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_167),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_840),
.Y(n_899)
);

BUFx10_ASAP7_75t_L g900 ( 
.A(n_638),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_770),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_237),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_506),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_172),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_133),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_833),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_569),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_431),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_210),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_68),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_448),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_524),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_534),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_757),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_137),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_806),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_590),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_740),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_760),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_374),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_391),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_407),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_53),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_767),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_171),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_823),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_314),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_7),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_101),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_127),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_677),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_465),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_293),
.Y(n_933)
);

CKINVDCx16_ASAP7_75t_R g934 ( 
.A(n_820),
.Y(n_934)
);

BUFx10_ASAP7_75t_L g935 ( 
.A(n_213),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_12),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_721),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_810),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_442),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_301),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_547),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_611),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_659),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_154),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_108),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_287),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_195),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_302),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_170),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_627),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_802),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_298),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_21),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_249),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_700),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_800),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_205),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_643),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_454),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_649),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_278),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_84),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_61),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_48),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_550),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_262),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_579),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_288),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_830),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_181),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_369),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_94),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_544),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_465),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_670),
.Y(n_975)
);

CKINVDCx14_ASAP7_75t_R g976 ( 
.A(n_24),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_756),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_328),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_826),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_718),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_5),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_648),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_208),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_415),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_401),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_17),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_88),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_386),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_688),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_402),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_814),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_292),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_648),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_299),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_53),
.Y(n_995)
);

BUFx10_ASAP7_75t_L g996 ( 
.A(n_816),
.Y(n_996)
);

CKINVDCx16_ASAP7_75t_R g997 ( 
.A(n_682),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_459),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_444),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_321),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_549),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_822),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_314),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_115),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_593),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_652),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_45),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_482),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_308),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_158),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_21),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_829),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_807),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_0),
.Y(n_1014)
);

BUFx2_ASAP7_75t_SL g1015 ( 
.A(n_235),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_788),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_804),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_611),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_215),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_808),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_23),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_150),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_334),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_78),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_799),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_739),
.Y(n_1026)
);

BUFx8_ASAP7_75t_SL g1027 ( 
.A(n_455),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_474),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_60),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_165),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_155),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_819),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_168),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_172),
.Y(n_1034)
);

BUFx10_ASAP7_75t_L g1035 ( 
.A(n_36),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_468),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_511),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_167),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_402),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_11),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_59),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_319),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_11),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_456),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_825),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_840),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_241),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_393),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_180),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_405),
.Y(n_1050)
);

BUFx8_ASAP7_75t_SL g1051 ( 
.A(n_666),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_776),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_345),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_684),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_95),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_66),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_249),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_506),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_348),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_610),
.Y(n_1060)
);

BUFx5_ASAP7_75t_L g1061 ( 
.A(n_112),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_584),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_258),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_21),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_759),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_331),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_431),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_272),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_676),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_515),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_599),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_350),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_126),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_389),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_44),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_436),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_803),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_138),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_403),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_268),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_365),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_823),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_761),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_793),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_254),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_382),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_428),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_541),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_600),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_30),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_707),
.Y(n_1091)
);

BUFx10_ASAP7_75t_L g1092 ( 
.A(n_135),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_513),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_827),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_276),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_837),
.Y(n_1096)
);

INVxp33_ASAP7_75t_R g1097 ( 
.A(n_87),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_566),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_817),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_700),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_364),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_173),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_421),
.Y(n_1103)
);

CKINVDCx14_ASAP7_75t_R g1104 ( 
.A(n_407),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_361),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_812),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_322),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_594),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_160),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_520),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_418),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_831),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_286),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_213),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_505),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_754),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_706),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_762),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_31),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_69),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_280),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_133),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_261),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_441),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_634),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_522),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_822),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_590),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_815),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_142),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_42),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_349),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_529),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_295),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_432),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_607),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_585),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_816),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_689),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_350),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_297),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_231),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_470),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_201),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_832),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_828),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_568),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_714),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_811),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_362),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_22),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_161),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_809),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_523),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_488),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_669),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_577),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_477),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_279),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_819),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_633),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_151),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_359),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_175),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_667),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_633),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_679),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_352),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_359),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_398),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_46),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_566),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_100),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_157),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_131),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_457),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_773),
.Y(n_1177)
);

BUFx5_ASAP7_75t_L g1178 ( 
.A(n_646),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_698),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_460),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_228),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_221),
.Y(n_1182)
);

BUFx10_ASAP7_75t_L g1183 ( 
.A(n_735),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_839),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_99),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_422),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_282),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_229),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_293),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_765),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_257),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_195),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_546),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_484),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_172),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_835),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_832),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_677),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_576),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_642),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_326),
.Y(n_1201)
);

BUFx5_ASAP7_75t_L g1202 ( 
.A(n_556),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_489),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_585),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_94),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_838),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_154),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_199),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_280),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_647),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_332),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_391),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_9),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_470),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_821),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_755),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_541),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_579),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_304),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_813),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_443),
.Y(n_1221)
);

CKINVDCx14_ASAP7_75t_R g1222 ( 
.A(n_743),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_844),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_12),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_257),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_598),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_743),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_818),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_528),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_612),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_52),
.Y(n_1231)
);

BUFx8_ASAP7_75t_SL g1232 ( 
.A(n_805),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_834),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_461),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_353),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_635),
.Y(n_1236)
);

CKINVDCx16_ASAP7_75t_R g1237 ( 
.A(n_256),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_671),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_304),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_345),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_616),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_772),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_796),
.Y(n_1243)
);

BUFx8_ASAP7_75t_SL g1244 ( 
.A(n_440),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_340),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_769),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_347),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_306),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_15),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_191),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_602),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_169),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_401),
.Y(n_1253)
);

BUFx5_ASAP7_75t_L g1254 ( 
.A(n_605),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_275),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_98),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_90),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_358),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_654),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_346),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_344),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_682),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_167),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_360),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_569),
.Y(n_1265)
);

BUFx5_ASAP7_75t_L g1266 ( 
.A(n_795),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_583),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_419),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_194),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_699),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_678),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_331),
.Y(n_1272)
);

BUFx10_ASAP7_75t_L g1273 ( 
.A(n_351),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_85),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_272),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_267),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_609),
.Y(n_1277)
);

INVxp33_ASAP7_75t_SL g1278 ( 
.A(n_1024),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1252),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1056),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_849),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_976),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1056),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_976),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_865),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_865),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_L g1287 ( 
.A(n_899),
.B(n_0),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_957),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_957),
.Y(n_1289)
);

NOR2xp67_ASAP7_75t_L g1290 ( 
.A(n_899),
.B(n_0),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_986),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_948),
.Y(n_1292)
);

CKINVDCx16_ASAP7_75t_R g1293 ( 
.A(n_883),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_948),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1223),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1223),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1120),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_883),
.B(n_1),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_854),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1104),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1104),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_928),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_944),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_956),
.B(n_978),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_861),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_861),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1222),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1120),
.Y(n_1308)
);

CKINVDCx16_ASAP7_75t_R g1309 ( 
.A(n_883),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_953),
.Y(n_1310)
);

INVxp67_ASAP7_75t_SL g1311 ( 
.A(n_1055),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_963),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_R g1313 ( 
.A(n_1222),
.B(n_1),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1027),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_970),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_972),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_983),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1004),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1185),
.Y(n_1319)
);

XOR2xp5_ASAP7_75t_L g1320 ( 
.A(n_1256),
.B(n_2),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1027),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1051),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1051),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1256),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1032),
.B(n_3),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1232),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1232),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1244),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1031),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1244),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1038),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_869),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1043),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1055),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1070),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1142),
.B(n_3),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_847),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1090),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_848),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_855),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_871),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1162),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1122),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_934),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1130),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1131),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_959),
.B(n_3),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1152),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1175),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1042),
.B(n_4),
.Y(n_1351)
);

INVxp33_ASAP7_75t_L g1352 ( 
.A(n_1066),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1195),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1207),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1102),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1208),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1213),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_997),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1231),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1102),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_880),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1234),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_891),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1237),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1263),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_860),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_860),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1235),
.B(n_4),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1162),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_849),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_909),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_862),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_862),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_935),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_864),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_893),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_904),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1151),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1343),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1355),
.B(n_910),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1281),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1293),
.B(n_935),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1370),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1355),
.B(n_915),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1311),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1334),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1280),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1283),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1285),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1360),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1360),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1286),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1377),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1343),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1378),
.B(n_923),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1279),
.B(n_847),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1292),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1294),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1378),
.B(n_925),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1295),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1296),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1278),
.B(n_929),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1309),
.B(n_936),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1339),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1371),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1374),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1299),
.Y(n_1408)
);

BUFx8_ASAP7_75t_L g1409 ( 
.A(n_1298),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1302),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1340),
.Y(n_1411)
);

NOR2x1_ASAP7_75t_L g1412 ( 
.A(n_1304),
.B(n_852),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1303),
.A2(n_905),
.B(n_898),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1352),
.B(n_947),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1310),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1312),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1342),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1315),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1361),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1316),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1369),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1317),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1369),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1318),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1329),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1363),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1376),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1331),
.B(n_945),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1333),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1338),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1335),
.B(n_947),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1282),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1344),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1341),
.B(n_1035),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1346),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1347),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1320),
.A2(n_890),
.B1(n_894),
.B2(n_872),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1349),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1350),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1353),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1354),
.B(n_949),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1356),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1357),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1359),
.A2(n_905),
.B(n_898),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1365),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1287),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1314),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1290),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1348),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1336),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1325),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1351),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1368),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1321),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1300),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1301),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1313),
.Y(n_1458)
);

INVx5_ASAP7_75t_L g1459 ( 
.A(n_1307),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1284),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1322),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1323),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1332),
.B(n_962),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1326),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1327),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1328),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1330),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1345),
.B(n_964),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1358),
.B(n_1082),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1362),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1288),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1364),
.B(n_852),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1289),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1291),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1297),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1305),
.Y(n_1476)
);

CKINVDCx16_ASAP7_75t_R g1477 ( 
.A(n_1306),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1308),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1319),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1324),
.A2(n_981),
.B1(n_995),
.B2(n_987),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1366),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1367),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1372),
.B(n_1061),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1373),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1375),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1343),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1343),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1311),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1311),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1281),
.A2(n_1030),
.B(n_1022),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1311),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1343),
.Y(n_1492)
);

AND2x6_ASAP7_75t_L g1493 ( 
.A(n_1298),
.B(n_866),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1293),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1311),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1281),
.A2(n_1257),
.B(n_1182),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1377),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1311),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1311),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1337),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1311),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1311),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1337),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1279),
.B(n_866),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1311),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1311),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1337),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1311),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1311),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1293),
.B(n_1061),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1293),
.B(n_1035),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1343),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1279),
.B(n_967),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1311),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1377),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1311),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1355),
.B(n_1007),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1343),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1311),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1311),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1377),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1339),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1337),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1355),
.B(n_1010),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1311),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1311),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1311),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1293),
.B(n_1061),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1293),
.B(n_1092),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1311),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1279),
.B(n_967),
.Y(n_1531)
);

BUFx8_ASAP7_75t_L g1532 ( 
.A(n_1377),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1311),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1313),
.B(n_1011),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1281),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1355),
.B(n_1014),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1293),
.B(n_1092),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1293),
.B(n_1061),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1377),
.Y(n_1539)
);

INVx4_ASAP7_75t_L g1540 ( 
.A(n_1494),
.Y(n_1540)
);

AND2x6_ASAP7_75t_L g1541 ( 
.A(n_1382),
.B(n_1182),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1413),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1445),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1394),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1388),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1497),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1432),
.A2(n_1274),
.B1(n_1269),
.B2(n_1021),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1539),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1511),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1452),
.A2(n_1061),
.B1(n_1162),
.B2(n_1029),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1496),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1490),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1532),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1529),
.B(n_971),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1446),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1380),
.B(n_1019),
.Y(n_1556)
);

NOR2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1537),
.B(n_1097),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1452),
.B(n_1033),
.Y(n_1558)
);

AND2x6_ASAP7_75t_L g1559 ( 
.A(n_1538),
.B(n_1162),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1427),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1453),
.B(n_1040),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1496),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1532),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1456),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1385),
.B(n_1041),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1389),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1453),
.B(n_1049),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1390),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1446),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1405),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1477),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1414),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1401),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1425),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1446),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1456),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1507),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1440),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1515),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1406),
.B(n_1064),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1417),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1393),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1398),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1456),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1399),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1402),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1522),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1523),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1435),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1404),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1523),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1386),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1407),
.B(n_971),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1517),
.B(n_1073),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1464),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1493),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1407),
.B(n_1000),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1387),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1500),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1454),
.B(n_1075),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1503),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1524),
.B(n_1078),
.Y(n_1602)
);

AO22x2_ASAP7_75t_L g1603 ( 
.A1(n_1480),
.A2(n_1015),
.B1(n_1034),
.B2(n_930),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1536),
.B(n_1109),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1433),
.B(n_894),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1493),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1391),
.B(n_1392),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1493),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1521),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1403),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1411),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1420),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_R g1613 ( 
.A(n_1448),
.B(n_1455),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1459),
.B(n_1192),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1488),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1396),
.B(n_1114),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1461),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1489),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1491),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1495),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1459),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1454),
.B(n_1119),
.Y(n_1622)
);

INVx4_ASAP7_75t_SL g1623 ( 
.A(n_1472),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1475),
.Y(n_1624)
);

BUFx4f_ASAP7_75t_L g1625 ( 
.A(n_1472),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1428),
.Y(n_1627)
);

BUFx10_ASAP7_75t_L g1628 ( 
.A(n_1469),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1400),
.B(n_1457),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1397),
.Y(n_1630)
);

BUFx10_ASAP7_75t_L g1631 ( 
.A(n_1458),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1501),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1504),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1504),
.B(n_1000),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1513),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1502),
.Y(n_1636)
);

BUFx10_ASAP7_75t_L g1637 ( 
.A(n_1465),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1513),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1505),
.B(n_1144),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1409),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1506),
.B(n_1164),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1531),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1534),
.B(n_1509),
.C(n_1508),
.Y(n_1643)
);

AO22x2_ASAP7_75t_L g1644 ( 
.A1(n_1481),
.A2(n_1224),
.B1(n_921),
.B2(n_926),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1531),
.B(n_1006),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1408),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1514),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1409),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1516),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1419),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1421),
.Y(n_1651)
);

AO22x2_ASAP7_75t_L g1652 ( 
.A1(n_1481),
.A2(n_921),
.B1(n_926),
.B2(n_914),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1519),
.B(n_1171),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1429),
.B(n_1173),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1447),
.B(n_1006),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1520),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1442),
.B(n_1174),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1473),
.B(n_914),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1525),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1526),
.B(n_1205),
.Y(n_1660)
);

CKINVDCx11_ASAP7_75t_R g1661 ( 
.A(n_1473),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1527),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1449),
.B(n_1249),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1530),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1450),
.B(n_1079),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1533),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1463),
.B(n_1250),
.Y(n_1667)
);

AND2x6_ASAP7_75t_L g1668 ( 
.A(n_1451),
.B(n_1079),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1510),
.B(n_1138),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1410),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1471),
.A2(n_965),
.B1(n_985),
.B2(n_940),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1415),
.B(n_849),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1528),
.B(n_1138),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1438),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1468),
.B(n_850),
.Y(n_1675)
);

INVx4_ASAP7_75t_SL g1676 ( 
.A(n_1467),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1430),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1431),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1483),
.A2(n_1271),
.B1(n_1277),
.B2(n_1268),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1462),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1434),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1436),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1441),
.A2(n_1187),
.B1(n_1146),
.B2(n_846),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1416),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1466),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1423),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1426),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1412),
.B(n_1187),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1437),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1439),
.Y(n_1690)
);

CKINVDCx20_ASAP7_75t_R g1691 ( 
.A(n_1474),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1474),
.Y(n_1693)
);

AND2x6_ASAP7_75t_L g1694 ( 
.A(n_1381),
.B(n_853),
.Y(n_1694)
);

AND2x6_ASAP7_75t_L g1695 ( 
.A(n_1384),
.B(n_853),
.Y(n_1695)
);

BUFx10_ASAP7_75t_L g1696 ( 
.A(n_1470),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1535),
.B(n_879),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1470),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1460),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1518),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1479),
.B(n_1178),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1379),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1518),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1518),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1484),
.B(n_900),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1482),
.B(n_856),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1476),
.B(n_1178),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1478),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1485),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1383),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1383),
.B(n_1178),
.Y(n_1711)
);

INVx4_ASAP7_75t_L g1712 ( 
.A(n_1395),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1395),
.B(n_1178),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1395),
.Y(n_1714)
);

BUFx4f_ASAP7_75t_L g1715 ( 
.A(n_1418),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1418),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1418),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1422),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1422),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1422),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1512),
.Y(n_1721)
);

AND2x6_ASAP7_75t_L g1722 ( 
.A(n_1424),
.B(n_863),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1486),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1486),
.Y(n_1724)
);

BUFx10_ASAP7_75t_L g1725 ( 
.A(n_1487),
.Y(n_1725)
);

AND2x6_ASAP7_75t_L g1726 ( 
.A(n_1487),
.B(n_863),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1492),
.B(n_1178),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1492),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1382),
.B(n_900),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1388),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1413),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1382),
.B(n_979),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1382),
.B(n_870),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1413),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1394),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1382),
.B(n_940),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1413),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1382),
.B(n_979),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1413),
.Y(n_1739)
);

AND2x2_ASAP7_75t_SL g1740 ( 
.A(n_1627),
.B(n_965),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_SL g1741 ( 
.A(n_1553),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1649),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1605),
.B(n_875),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1560),
.B(n_985),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1547),
.A2(n_859),
.B1(n_902),
.B2(n_858),
.C(n_851),
.Y(n_1745)
);

AO22x2_ASAP7_75t_L g1746 ( 
.A1(n_1581),
.A2(n_1071),
.B1(n_1081),
.B2(n_1008),
.Y(n_1746)
);

AO22x2_ASAP7_75t_L g1747 ( 
.A1(n_1612),
.A2(n_1071),
.B1(n_1081),
.B2(n_1008),
.Y(n_1747)
);

AO22x2_ASAP7_75t_L g1748 ( 
.A1(n_1623),
.A2(n_1106),
.B1(n_1108),
.B2(n_1101),
.Y(n_1748)
);

BUFx8_ASAP7_75t_L g1749 ( 
.A(n_1648),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1733),
.A2(n_867),
.B1(n_868),
.B2(n_857),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1563),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1570),
.B(n_1111),
.Y(n_1752)
);

BUFx8_ASAP7_75t_L g1753 ( 
.A(n_1680),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1579),
.B(n_1111),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1656),
.Y(n_1755)
);

AO22x2_ASAP7_75t_L g1756 ( 
.A1(n_1652),
.A2(n_1128),
.B1(n_1134),
.B2(n_1117),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1579),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1656),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1609),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1733),
.A2(n_874),
.B1(n_876),
.B2(n_873),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1670),
.B(n_878),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1596),
.B(n_884),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1609),
.B(n_1117),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1662),
.Y(n_1764)
);

AO22x2_ASAP7_75t_L g1765 ( 
.A1(n_1652),
.A2(n_1134),
.B1(n_1143),
.B2(n_1128),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1605),
.B(n_875),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1587),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1627),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1662),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1664),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1558),
.B(n_886),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1564),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1590),
.A2(n_895),
.B1(n_901),
.B2(n_892),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1549),
.A2(n_1153),
.B1(n_1181),
.B2(n_1013),
.C(n_994),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1613),
.Y(n_1775)
);

AO22x2_ASAP7_75t_L g1776 ( 
.A1(n_1644),
.A2(n_1166),
.B1(n_1218),
.B2(n_1143),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1548),
.B(n_1166),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1610),
.A2(n_907),
.B1(n_908),
.B2(n_906),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1592),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1617),
.Y(n_1780)
);

NAND2x1p5_ASAP7_75t_L g1781 ( 
.A(n_1540),
.B(n_1196),
.Y(n_1781)
);

AO22x2_ASAP7_75t_L g1782 ( 
.A1(n_1644),
.A2(n_1241),
.B1(n_1265),
.B2(n_1218),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1735),
.B(n_1241),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1561),
.B(n_912),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1680),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1589),
.A2(n_916),
.B1(n_917),
.B2(n_913),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1611),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1659),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1572),
.A2(n_924),
.B1(n_927),
.B2(n_918),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1564),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1666),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1598),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1544),
.B(n_1265),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1595),
.B(n_1229),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1615),
.Y(n_1795)
);

AO22x2_ASAP7_75t_L g1796 ( 
.A1(n_1671),
.A2(n_1551),
.B1(n_1562),
.B2(n_1546),
.Y(n_1796)
);

AO22x2_ASAP7_75t_L g1797 ( 
.A1(n_1551),
.A2(n_1276),
.B1(n_1270),
.B2(n_1246),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1699),
.B(n_1270),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1618),
.Y(n_1799)
);

AO22x2_ASAP7_75t_L g1800 ( 
.A1(n_1562),
.A2(n_1276),
.B1(n_1247),
.B2(n_1272),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1619),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1620),
.Y(n_1802)
);

NAND2x1p5_ASAP7_75t_L g1803 ( 
.A(n_1693),
.B(n_1239),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1729),
.B(n_996),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1632),
.Y(n_1805)
);

AO22x2_ASAP7_75t_L g1806 ( 
.A1(n_1603),
.A2(n_882),
.B1(n_885),
.B2(n_877),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1596),
.B(n_931),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1736),
.B(n_932),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1636),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1567),
.A2(n_887),
.B(n_896),
.C(n_888),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1732),
.B(n_897),
.Y(n_1811)
);

AO22x2_ASAP7_75t_L g1812 ( 
.A1(n_1603),
.A2(n_903),
.B1(n_920),
.B2(n_919),
.Y(n_1812)
);

BUFx8_ASAP7_75t_L g1813 ( 
.A(n_1709),
.Y(n_1813)
);

AO22x2_ASAP7_75t_L g1814 ( 
.A1(n_1554),
.A2(n_938),
.B1(n_941),
.B2(n_933),
.Y(n_1814)
);

OR2x6_ASAP7_75t_SL g1815 ( 
.A(n_1640),
.B(n_937),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1616),
.B(n_939),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1629),
.B(n_942),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1647),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1582),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1580),
.B(n_943),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1738),
.B(n_946),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1583),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1571),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1585),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1586),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1684),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1686),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1667),
.B(n_996),
.Y(n_1828)
);

INVx4_ASAP7_75t_L g1829 ( 
.A(n_1576),
.Y(n_1829)
);

BUFx8_ASAP7_75t_L g1830 ( 
.A(n_1541),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1687),
.Y(n_1831)
);

AO22x2_ASAP7_75t_L g1832 ( 
.A1(n_1554),
.A2(n_955),
.B1(n_960),
.B2(n_950),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1658),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1689),
.Y(n_1834)
);

AO22x2_ASAP7_75t_L g1835 ( 
.A1(n_1706),
.A2(n_966),
.B1(n_968),
.B2(n_961),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1690),
.Y(n_1836)
);

OAI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1625),
.A2(n_954),
.B1(n_958),
.B2(n_952),
.C(n_951),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1706),
.A2(n_973),
.B1(n_974),
.B2(n_969),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1607),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1626),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1692),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1593),
.Y(n_1842)
);

AO22x2_ASAP7_75t_L g1843 ( 
.A1(n_1634),
.A2(n_977),
.B1(n_980),
.B2(n_975),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1736),
.B(n_1113),
.Y(n_1844)
);

BUFx8_ASAP7_75t_L g1845 ( 
.A(n_1584),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1658),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1593),
.Y(n_1847)
);

AO22x2_ASAP7_75t_L g1848 ( 
.A1(n_1634),
.A2(n_984),
.B1(n_988),
.B2(n_982),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1597),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1597),
.Y(n_1850)
);

NOR2xp67_ASAP7_75t_L g1851 ( 
.A(n_1624),
.B(n_6),
.Y(n_1851)
);

BUFx8_ASAP7_75t_L g1852 ( 
.A(n_1685),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1545),
.Y(n_1853)
);

AO22x2_ASAP7_75t_L g1854 ( 
.A1(n_1645),
.A2(n_999),
.B1(n_1003),
.B2(n_998),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1566),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1568),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1573),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1691),
.B(n_1009),
.Y(n_1858)
);

AO22x2_ASAP7_75t_L g1859 ( 
.A1(n_1645),
.A2(n_1016),
.B1(n_1017),
.B2(n_1012),
.Y(n_1859)
);

BUFx8_ASAP7_75t_L g1860 ( 
.A(n_1685),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1730),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1556),
.B(n_989),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1661),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1638),
.B(n_1675),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1628),
.B(n_1113),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1705),
.A2(n_991),
.B1(n_992),
.B2(n_990),
.Y(n_1866)
);

XNOR2xp5_ASAP7_75t_L g1867 ( 
.A(n_1557),
.B(n_6),
.Y(n_1867)
);

AO22x2_ASAP7_75t_L g1868 ( 
.A1(n_1633),
.A2(n_1039),
.B1(n_1046),
.B2(n_1036),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1677),
.Y(n_1869)
);

CKINVDCx11_ASAP7_75t_R g1870 ( 
.A(n_1696),
.Y(n_1870)
);

AO22x2_ASAP7_75t_L g1871 ( 
.A1(n_1606),
.A2(n_1050),
.B1(n_1060),
.B2(n_1047),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1698),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1646),
.Y(n_1873)
);

AND2x6_ASAP7_75t_L g1874 ( 
.A(n_1608),
.B(n_889),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1565),
.B(n_993),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1650),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1651),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1594),
.B(n_1602),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1604),
.B(n_1005),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1678),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1681),
.Y(n_1881)
);

AO22x2_ASAP7_75t_L g1882 ( 
.A1(n_1734),
.A2(n_1067),
.B1(n_1074),
.B2(n_1063),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1639),
.B(n_1641),
.Y(n_1883)
);

OAI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1614),
.A2(n_1020),
.B1(n_1023),
.B2(n_1018),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1628),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1682),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1694),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1621),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1574),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1694),
.Y(n_1890)
);

AO22x2_ASAP7_75t_L g1891 ( 
.A1(n_1734),
.A2(n_1083),
.B1(n_1084),
.B2(n_1077),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1578),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1676),
.B(n_1642),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1676),
.B(n_1085),
.Y(n_1894)
);

AO22x2_ASAP7_75t_L g1895 ( 
.A1(n_1643),
.A2(n_1087),
.B1(n_1088),
.B2(n_1086),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1696),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1708),
.B(n_1089),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1653),
.B(n_1026),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1672),
.Y(n_1899)
);

BUFx8_ASAP7_75t_L g1900 ( 
.A(n_1688),
.Y(n_1900)
);

AO22x2_ASAP7_75t_L g1901 ( 
.A1(n_1655),
.A2(n_1099),
.B1(n_1100),
.B2(n_1093),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1660),
.B(n_1028),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1543),
.Y(n_1903)
);

BUFx8_ASAP7_75t_L g1904 ( 
.A(n_1688),
.Y(n_1904)
);

INVxp33_ASAP7_75t_SL g1905 ( 
.A(n_1674),
.Y(n_1905)
);

BUFx8_ASAP7_75t_L g1906 ( 
.A(n_1668),
.Y(n_1906)
);

NAND2x1p5_ASAP7_75t_L g1907 ( 
.A(n_1630),
.B(n_1112),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1665),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1631),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1694),
.B(n_1037),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_1630),
.B(n_1115),
.Y(n_1911)
);

AO22x2_ASAP7_75t_L g1912 ( 
.A1(n_1669),
.A2(n_1673),
.B1(n_1701),
.B2(n_1731),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1695),
.B(n_1044),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1637),
.Y(n_1914)
);

OAI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1679),
.A2(n_1683),
.B1(n_1707),
.B2(n_1657),
.C(n_1654),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1695),
.B(n_1045),
.Y(n_1916)
);

AO22x2_ASAP7_75t_L g1917 ( 
.A1(n_1669),
.A2(n_1136),
.B1(n_1140),
.B2(n_1118),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1737),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1559),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1673),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1635),
.B(n_1141),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1599),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1739),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1631),
.B(n_1048),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1588),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1601),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1637),
.Y(n_1927)
);

NAND2x1p5_ASAP7_75t_L g1928 ( 
.A(n_1715),
.B(n_1145),
.Y(n_1928)
);

AO22x2_ASAP7_75t_L g1929 ( 
.A1(n_1600),
.A2(n_1148),
.B1(n_1156),
.B2(n_1147),
.Y(n_1929)
);

AO22x2_ASAP7_75t_L g1930 ( 
.A1(n_1622),
.A2(n_1168),
.B1(n_1170),
.B2(n_1158),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1552),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1550),
.B(n_1052),
.Y(n_1932)
);

AO22x2_ASAP7_75t_L g1933 ( 
.A1(n_1577),
.A2(n_1184),
.B1(n_1188),
.B2(n_1172),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1591),
.B(n_1154),
.Y(n_1934)
);

AO22x2_ASAP7_75t_L g1935 ( 
.A1(n_1663),
.A2(n_1200),
.B1(n_1204),
.B2(n_1191),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1668),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1668),
.Y(n_1937)
);

AO22x2_ASAP7_75t_L g1938 ( 
.A1(n_1559),
.A2(n_1220),
.B1(n_1221),
.B2(n_1216),
.Y(n_1938)
);

BUFx8_ASAP7_75t_L g1939 ( 
.A(n_1722),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1542),
.Y(n_1940)
);

AO22x2_ASAP7_75t_L g1941 ( 
.A1(n_1555),
.A2(n_1226),
.B1(n_1236),
.B2(n_1225),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1722),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1569),
.B(n_1248),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1722),
.Y(n_1944)
);

OAI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1697),
.A2(n_1057),
.B1(n_1058),
.B2(n_1054),
.C(n_1053),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1711),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1713),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1727),
.Y(n_1948)
);

AO22x2_ASAP7_75t_L g1949 ( 
.A1(n_1575),
.A2(n_1260),
.B1(n_1275),
.B2(n_1255),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1726),
.Y(n_1950)
);

AO22x2_ASAP7_75t_L g1951 ( 
.A1(n_1712),
.A2(n_911),
.B1(n_1001),
.B2(n_889),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1726),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1725),
.Y(n_1953)
);

OAI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1728),
.A2(n_1065),
.B1(n_1068),
.B2(n_1062),
.C(n_1059),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1719),
.B(n_1072),
.Y(n_1955)
);

OA22x2_ASAP7_75t_L g1956 ( 
.A1(n_1716),
.A2(n_1076),
.B1(n_1080),
.B2(n_1069),
.Y(n_1956)
);

AO22x2_ASAP7_75t_L g1957 ( 
.A1(n_1710),
.A2(n_1002),
.B1(n_1025),
.B2(n_1001),
.Y(n_1957)
);

AO22x2_ASAP7_75t_L g1958 ( 
.A1(n_1710),
.A2(n_1025),
.B1(n_1135),
.B2(n_1002),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1714),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1700),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1702),
.Y(n_1961)
);

BUFx8_ASAP7_75t_L g1962 ( 
.A(n_1703),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1704),
.A2(n_1094),
.B1(n_1095),
.B2(n_1091),
.Y(n_1963)
);

AO22x2_ASAP7_75t_L g1964 ( 
.A1(n_1718),
.A2(n_1150),
.B1(n_1253),
.B2(n_1149),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1717),
.B(n_1154),
.Y(n_1965)
);

AO22x2_ASAP7_75t_L g1966 ( 
.A1(n_1720),
.A2(n_1150),
.B1(n_1253),
.B2(n_1149),
.Y(n_1966)
);

BUFx8_ASAP7_75t_L g1967 ( 
.A(n_1721),
.Y(n_1967)
);

AO22x2_ASAP7_75t_L g1968 ( 
.A1(n_1724),
.A2(n_1262),
.B1(n_1267),
.B2(n_1261),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1841),
.B(n_1096),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1785),
.B(n_1098),
.Y(n_1970)
);

NAND2xp33_ASAP7_75t_SL g1971 ( 
.A(n_1890),
.B(n_1133),
.Y(n_1971)
);

NAND2xp33_ASAP7_75t_SL g1972 ( 
.A(n_1772),
.B(n_1133),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1757),
.B(n_1759),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1914),
.B(n_1103),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1927),
.B(n_1105),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1839),
.B(n_1840),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1768),
.B(n_1107),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1909),
.B(n_1261),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1787),
.B(n_1110),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1753),
.B(n_1872),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1767),
.B(n_1116),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1772),
.B(n_1121),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1790),
.B(n_1258),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1790),
.B(n_1259),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_SL g1985 ( 
.A(n_1887),
.B(n_1190),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1896),
.B(n_1123),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1744),
.B(n_1264),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1798),
.B(n_1124),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1781),
.B(n_1125),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1813),
.B(n_1126),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1819),
.B(n_1262),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1883),
.B(n_1127),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1878),
.B(n_1129),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1794),
.B(n_1132),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1740),
.B(n_1137),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1752),
.B(n_1139),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1754),
.B(n_1155),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1763),
.B(n_1157),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1792),
.B(n_1159),
.Y(n_1999)
);

NAND2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1742),
.B(n_881),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1795),
.B(n_1160),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1799),
.B(n_1161),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1822),
.B(n_1267),
.Y(n_2003)
);

NAND2xp33_ASAP7_75t_SL g2004 ( 
.A(n_1755),
.B(n_922),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1801),
.B(n_1163),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1884),
.B(n_1165),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1924),
.B(n_1167),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1788),
.B(n_1791),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1885),
.B(n_1169),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1803),
.B(n_1176),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1865),
.B(n_1177),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1780),
.B(n_1828),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1802),
.B(n_1179),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1830),
.B(n_1180),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1778),
.B(n_1238),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1928),
.B(n_1240),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1944),
.B(n_1186),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1793),
.B(n_1243),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1852),
.B(n_1245),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1860),
.B(n_1251),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1864),
.B(n_1189),
.Y(n_2021)
);

NAND2xp33_ASAP7_75t_SL g2022 ( 
.A(n_1775),
.B(n_1193),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1845),
.B(n_1194),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1805),
.B(n_1197),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1773),
.B(n_1198),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1955),
.B(n_1777),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1783),
.B(n_1199),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1919),
.B(n_1201),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1824),
.B(n_8),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1786),
.B(n_1206),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1789),
.B(n_1209),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1851),
.B(n_1228),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1835),
.B(n_1154),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_SL g2034 ( 
.A(n_1829),
.B(n_1210),
.Y(n_2034)
);

NAND2xp33_ASAP7_75t_SL g2035 ( 
.A(n_1953),
.B(n_1211),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1761),
.B(n_1212),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1963),
.B(n_1214),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1907),
.B(n_1215),
.Y(n_2038)
);

NAND2xp33_ASAP7_75t_SL g2039 ( 
.A(n_1952),
.B(n_1217),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1809),
.B(n_1219),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1911),
.B(n_1230),
.Y(n_2041)
);

NAND2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1942),
.B(n_1233),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1897),
.B(n_1750),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1825),
.B(n_8),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1760),
.B(n_1242),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1910),
.B(n_1183),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1826),
.B(n_1827),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1913),
.B(n_1183),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1808),
.B(n_1846),
.Y(n_2049)
);

NAND2xp33_ASAP7_75t_SL g2050 ( 
.A(n_1758),
.B(n_922),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1916),
.B(n_1183),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1925),
.B(n_1273),
.Y(n_2052)
);

NAND2xp33_ASAP7_75t_SL g2053 ( 
.A(n_1764),
.B(n_922),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1866),
.B(n_1804),
.Y(n_2054)
);

NAND2xp33_ASAP7_75t_SL g2055 ( 
.A(n_1769),
.B(n_1133),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1906),
.B(n_1202),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_SL g2057 ( 
.A(n_1770),
.B(n_1190),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1835),
.B(n_1254),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_SL g2059 ( 
.A(n_1831),
.B(n_1190),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1838),
.B(n_1266),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_SL g2061 ( 
.A(n_1834),
.B(n_1190),
.Y(n_2061)
);

NAND2xp33_ASAP7_75t_SL g2062 ( 
.A(n_1836),
.B(n_1227),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1743),
.B(n_1766),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1811),
.B(n_1821),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1818),
.B(n_9),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1817),
.B(n_1723),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1797),
.B(n_9),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1934),
.B(n_11),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1894),
.B(n_13),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_1833),
.B(n_13),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1797),
.B(n_10),
.Y(n_2071)
);

NAND2xp33_ASAP7_75t_SL g2072 ( 
.A(n_1779),
.B(n_10),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1810),
.B(n_10),
.Y(n_2073)
);

AND2x2_ASAP7_75t_SL g2074 ( 
.A(n_1938),
.B(n_14),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1868),
.B(n_1933),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1868),
.B(n_14),
.Y(n_2076)
);

NAND2xp33_ASAP7_75t_SL g2077 ( 
.A(n_1741),
.B(n_16),
.Y(n_2077)
);

NAND2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1862),
.B(n_18),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1933),
.B(n_19),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1776),
.B(n_19),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1920),
.B(n_19),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1899),
.B(n_22),
.Y(n_2082)
);

NAND2xp33_ASAP7_75t_SL g2083 ( 
.A(n_1875),
.B(n_20),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_SL g2084 ( 
.A(n_1879),
.B(n_20),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1853),
.B(n_23),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1855),
.B(n_24),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1856),
.B(n_25),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1956),
.B(n_26),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1893),
.B(n_26),
.Y(n_2089)
);

NAND2xp33_ASAP7_75t_SL g2090 ( 
.A(n_1903),
.B(n_25),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1857),
.B(n_27),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1861),
.B(n_27),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1820),
.B(n_28),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1898),
.B(n_1902),
.Y(n_2094)
);

NAND2xp33_ASAP7_75t_SL g2095 ( 
.A(n_1918),
.B(n_27),
.Y(n_2095)
);

NAND2xp33_ASAP7_75t_SL g2096 ( 
.A(n_1923),
.B(n_28),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_SL g2097 ( 
.A(n_1931),
.B(n_29),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1869),
.B(n_29),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1842),
.B(n_31),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1844),
.B(n_33),
.Y(n_2100)
);

NAND2xp33_ASAP7_75t_SL g2101 ( 
.A(n_1959),
.B(n_32),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1921),
.B(n_35),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1816),
.B(n_35),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1847),
.B(n_34),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1849),
.B(n_34),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1900),
.B(n_35),
.Y(n_2106)
);

NAND2xp33_ASAP7_75t_SL g2107 ( 
.A(n_1936),
.B(n_34),
.Y(n_2107)
);

NAND2xp33_ASAP7_75t_SL g2108 ( 
.A(n_1937),
.B(n_36),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1850),
.B(n_36),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1904),
.B(n_1771),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1917),
.B(n_37),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1784),
.B(n_38),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1888),
.B(n_38),
.Y(n_2113)
);

NAND2xp33_ASAP7_75t_SL g2114 ( 
.A(n_1873),
.B(n_37),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1743),
.B(n_1766),
.Y(n_2115)
);

NAND2xp33_ASAP7_75t_SL g2116 ( 
.A(n_1876),
.B(n_37),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1965),
.B(n_40),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1917),
.B(n_39),
.Y(n_2118)
);

NAND2xp33_ASAP7_75t_SL g2119 ( 
.A(n_1877),
.B(n_41),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1880),
.B(n_42),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1881),
.B(n_42),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1886),
.B(n_43),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1751),
.B(n_43),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1932),
.B(n_1939),
.Y(n_2124)
);

NAND2xp33_ASAP7_75t_SL g2125 ( 
.A(n_1940),
.B(n_41),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1882),
.B(n_46),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_SL g2127 ( 
.A(n_1863),
.B(n_48),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1922),
.B(n_49),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1889),
.B(n_48),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1926),
.B(n_50),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1776),
.B(n_49),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1882),
.B(n_49),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1943),
.B(n_51),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1858),
.B(n_51),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1962),
.B(n_51),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1967),
.B(n_52),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1908),
.B(n_52),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1891),
.B(n_53),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1782),
.B(n_1747),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1905),
.B(n_55),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1946),
.B(n_56),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1947),
.B(n_56),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1814),
.B(n_54),
.Y(n_2143)
);

NAND2xp33_ASAP7_75t_SL g2144 ( 
.A(n_1950),
.B(n_54),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1948),
.B(n_56),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1782),
.B(n_54),
.Y(n_2146)
);

NAND2xp33_ASAP7_75t_SL g2147 ( 
.A(n_1870),
.B(n_57),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1892),
.B(n_57),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1814),
.B(n_57),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1832),
.B(n_58),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1749),
.B(n_59),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1832),
.B(n_1935),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1762),
.B(n_1807),
.Y(n_2153)
);

NAND2xp33_ASAP7_75t_SL g2154 ( 
.A(n_1823),
.B(n_60),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1960),
.B(n_62),
.Y(n_2155)
);

XNOR2xp5_ASAP7_75t_L g2156 ( 
.A(n_1756),
.B(n_61),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1961),
.B(n_62),
.Y(n_2157)
);

NAND2xp33_ASAP7_75t_SL g2158 ( 
.A(n_1938),
.B(n_1867),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_SL g2159 ( 
.A(n_1796),
.B(n_61),
.Y(n_2159)
);

NAND2xp33_ASAP7_75t_SL g2160 ( 
.A(n_1796),
.B(n_1748),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1929),
.B(n_63),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1929),
.B(n_64),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1815),
.B(n_1941),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1941),
.B(n_65),
.Y(n_2164)
);

NAND2xp33_ASAP7_75t_SL g2165 ( 
.A(n_1748),
.B(n_64),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1949),
.B(n_66),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1930),
.B(n_64),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_SL g2168 ( 
.A(n_1949),
.B(n_67),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1837),
.B(n_67),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1871),
.B(n_67),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1871),
.B(n_68),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1800),
.B(n_69),
.Y(n_2172)
);

NAND2xp33_ASAP7_75t_SL g2173 ( 
.A(n_1800),
.B(n_66),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1874),
.B(n_71),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1874),
.B(n_71),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1954),
.B(n_72),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1930),
.B(n_72),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1843),
.B(n_72),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1843),
.B(n_73),
.Y(n_2179)
);

NAND2xp33_ASAP7_75t_SL g2180 ( 
.A(n_1806),
.B(n_70),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1848),
.B(n_73),
.Y(n_2181)
);

NAND2xp33_ASAP7_75t_SL g2182 ( 
.A(n_1806),
.B(n_1812),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1848),
.B(n_70),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_1854),
.B(n_73),
.Y(n_2184)
);

NAND2xp33_ASAP7_75t_SL g2185 ( 
.A(n_1812),
.B(n_70),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1854),
.B(n_75),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1859),
.B(n_74),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1859),
.B(n_75),
.Y(n_2188)
);

NAND2xp33_ASAP7_75t_SL g2189 ( 
.A(n_1957),
.B(n_1958),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1912),
.B(n_74),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1951),
.B(n_75),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_1912),
.B(n_74),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1957),
.B(n_77),
.Y(n_2193)
);

NAND2xp33_ASAP7_75t_SL g2194 ( 
.A(n_1901),
.B(n_76),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1901),
.B(n_79),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1895),
.B(n_78),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1895),
.B(n_79),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1964),
.B(n_79),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1964),
.B(n_80),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1747),
.B(n_80),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1966),
.B(n_81),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1746),
.B(n_80),
.Y(n_2202)
);

NAND2xp33_ASAP7_75t_SL g2203 ( 
.A(n_1968),
.B(n_81),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1915),
.B(n_82),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_1774),
.B(n_83),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1945),
.B(n_83),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1745),
.B(n_84),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1746),
.B(n_82),
.Y(n_2208)
);

NAND2xp33_ASAP7_75t_SL g2209 ( 
.A(n_1756),
.B(n_1765),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1785),
.B(n_86),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1841),
.B(n_85),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_1785),
.B(n_85),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1785),
.B(n_87),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1785),
.B(n_88),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1841),
.B(n_86),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_1785),
.B(n_88),
.Y(n_2216)
);

NAND2xp33_ASAP7_75t_SL g2217 ( 
.A(n_1890),
.B(n_86),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1841),
.B(n_89),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1785),
.B(n_90),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1785),
.B(n_89),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_1785),
.B(n_90),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1785),
.B(n_91),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1785),
.B(n_92),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_1785),
.B(n_92),
.Y(n_2224)
);

NAND2xp33_ASAP7_75t_SL g2225 ( 
.A(n_1914),
.B(n_89),
.Y(n_2225)
);

NAND2xp33_ASAP7_75t_SL g2226 ( 
.A(n_1914),
.B(n_92),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1785),
.B(n_95),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1785),
.B(n_95),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_1785),
.B(n_96),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_1785),
.B(n_93),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1841),
.B(n_93),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1785),
.B(n_97),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1785),
.B(n_97),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_1785),
.B(n_97),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1785),
.B(n_98),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1785),
.B(n_98),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1785),
.B(n_99),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_SL g2238 ( 
.A(n_1785),
.B(n_99),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1841),
.B(n_96),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_1785),
.B(n_100),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1785),
.B(n_100),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1785),
.B(n_101),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1785),
.B(n_102),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1785),
.B(n_96),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_1785),
.B(n_103),
.Y(n_2245)
);

NAND2xp33_ASAP7_75t_SL g2246 ( 
.A(n_1914),
.B(n_102),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_1785),
.B(n_104),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1785),
.B(n_104),
.Y(n_2248)
);

NAND2xp33_ASAP7_75t_SL g2249 ( 
.A(n_1914),
.B(n_103),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_1785),
.B(n_105),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1785),
.B(n_106),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1785),
.B(n_106),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1785),
.B(n_106),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_1785),
.B(n_107),
.Y(n_2254)
);

NAND2xp33_ASAP7_75t_SL g2255 ( 
.A(n_1914),
.B(n_104),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1841),
.B(n_107),
.Y(n_2256)
);

NAND2xp33_ASAP7_75t_SL g2257 ( 
.A(n_1914),
.B(n_107),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_1785),
.B(n_108),
.Y(n_2258)
);

NAND2xp33_ASAP7_75t_SL g2259 ( 
.A(n_1914),
.B(n_108),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_1785),
.B(n_110),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_1785),
.B(n_110),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_1785),
.B(n_111),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_1785),
.B(n_111),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1841),
.B(n_109),
.Y(n_2264)
);

NAND2xp33_ASAP7_75t_SL g2265 ( 
.A(n_1914),
.B(n_109),
.Y(n_2265)
);

NAND2xp33_ASAP7_75t_SL g2266 ( 
.A(n_1914),
.B(n_109),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_1785),
.B(n_113),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_1785),
.B(n_113),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_SL g2269 ( 
.A(n_1914),
.B(n_112),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_1785),
.B(n_114),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_1785),
.B(n_114),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_1785),
.B(n_115),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1841),
.B(n_113),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_1785),
.B(n_117),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1785),
.B(n_117),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_1785),
.B(n_117),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_1785),
.B(n_118),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_1785),
.B(n_119),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_1785),
.B(n_119),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_1785),
.B(n_119),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1785),
.B(n_120),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1785),
.B(n_120),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_1785),
.B(n_121),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1785),
.B(n_121),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_1785),
.B(n_121),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_1841),
.B(n_116),
.Y(n_2286)
);

NAND2xp33_ASAP7_75t_SL g2287 ( 
.A(n_1914),
.B(n_116),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_1785),
.B(n_116),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1841),
.B(n_122),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_1785),
.B(n_123),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_1785),
.B(n_123),
.Y(n_2291)
);

NAND2xp33_ASAP7_75t_SL g2292 ( 
.A(n_1914),
.B(n_122),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_1785),
.B(n_124),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_1785),
.B(n_124),
.Y(n_2294)
);

NAND2xp33_ASAP7_75t_SL g2295 ( 
.A(n_1914),
.B(n_122),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_1785),
.B(n_125),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_SL g2297 ( 
.A(n_1914),
.B(n_124),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_1785),
.B(n_126),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_1785),
.B(n_126),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_1785),
.B(n_127),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_1785),
.B(n_127),
.Y(n_2301)
);

NAND2xp33_ASAP7_75t_SL g2302 ( 
.A(n_1914),
.B(n_125),
.Y(n_2302)
);

NAND2xp33_ASAP7_75t_SL g2303 ( 
.A(n_1914),
.B(n_128),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_1785),
.B(n_129),
.Y(n_2304)
);

NAND2xp33_ASAP7_75t_SL g2305 ( 
.A(n_1914),
.B(n_128),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1785),
.B(n_128),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_SL g2307 ( 
.A(n_1914),
.B(n_129),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_1785),
.B(n_130),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_1785),
.B(n_129),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1841),
.B(n_130),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1785),
.B(n_131),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1841),
.B(n_130),
.Y(n_2312)
);

NAND2xp33_ASAP7_75t_SL g2313 ( 
.A(n_1890),
.B(n_131),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1841),
.B(n_132),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_1841),
.B(n_132),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1841),
.B(n_132),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_1841),
.B(n_134),
.Y(n_2317)
);

NAND2xp33_ASAP7_75t_SL g2318 ( 
.A(n_1890),
.B(n_134),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_1785),
.B(n_134),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_1785),
.B(n_137),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1785),
.B(n_137),
.Y(n_2321)
);

NAND2xp33_ASAP7_75t_SL g2322 ( 
.A(n_1890),
.B(n_136),
.Y(n_2322)
);

XNOR2xp5_ASAP7_75t_L g2323 ( 
.A(n_1756),
.B(n_136),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1785),
.B(n_139),
.Y(n_2324)
);

NAND2xp33_ASAP7_75t_SL g2325 ( 
.A(n_1890),
.B(n_138),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1841),
.B(n_138),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_1785),
.B(n_141),
.Y(n_2327)
);

AND3x1_ASAP7_75t_L g2328 ( 
.A(n_1754),
.B(n_140),
.C(n_141),
.Y(n_2328)
);

NAND2xp33_ASAP7_75t_SL g2329 ( 
.A(n_1890),
.B(n_141),
.Y(n_2329)
);

NAND2xp33_ASAP7_75t_SL g2330 ( 
.A(n_1890),
.B(n_143),
.Y(n_2330)
);

NAND2xp33_ASAP7_75t_SL g2331 ( 
.A(n_1890),
.B(n_143),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_1785),
.B(n_144),
.Y(n_2332)
);

NAND2xp33_ASAP7_75t_SL g2333 ( 
.A(n_1890),
.B(n_143),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_1785),
.B(n_146),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_1785),
.B(n_146),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_1785),
.B(n_147),
.Y(n_2336)
);

NAND2xp33_ASAP7_75t_SL g2337 ( 
.A(n_1890),
.B(n_145),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_SL g2338 ( 
.A(n_1785),
.B(n_147),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_1785),
.B(n_147),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1785),
.B(n_148),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_1841),
.B(n_145),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1841),
.B(n_145),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1785),
.B(n_149),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_1785),
.B(n_149),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_SL g2345 ( 
.A(n_1890),
.B(n_148),
.Y(n_2345)
);

NAND2xp33_ASAP7_75t_SL g2346 ( 
.A(n_1890),
.B(n_148),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_1785),
.B(n_149),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_1785),
.B(n_151),
.Y(n_2348)
);

NAND2xp33_ASAP7_75t_SL g2349 ( 
.A(n_1890),
.B(n_150),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_1785),
.B(n_151),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_1785),
.B(n_152),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_1890),
.B(n_150),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_1785),
.B(n_153),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1841),
.B(n_152),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_1785),
.B(n_152),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_1785),
.B(n_155),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1785),
.B(n_155),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_1785),
.B(n_156),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1841),
.B(n_154),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_1785),
.B(n_157),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_1785),
.B(n_158),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1785),
.B(n_158),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1841),
.B(n_156),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_1785),
.B(n_159),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_1785),
.B(n_159),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_1785),
.B(n_159),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_1785),
.B(n_160),
.Y(n_2367)
);

NAND2xp33_ASAP7_75t_SL g2368 ( 
.A(n_1890),
.B(n_156),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_1785),
.B(n_161),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_1785),
.B(n_161),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_1785),
.B(n_162),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1976),
.B(n_160),
.Y(n_2372)
);

OAI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2204),
.A2(n_163),
.B(n_164),
.Y(n_2373)
);

INVxp67_ASAP7_75t_SL g2374 ( 
.A(n_2273),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2047),
.Y(n_2375)
);

OAI22x1_ASAP7_75t_L g2376 ( 
.A1(n_2156),
.A2(n_2323),
.B1(n_2163),
.B2(n_2172),
.Y(n_2376)
);

OAI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_1993),
.A2(n_166),
.B(n_169),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2047),
.B(n_2054),
.Y(n_2378)
);

BUFx10_ASAP7_75t_L g2379 ( 
.A(n_2273),
.Y(n_2379)
);

NOR2x1_ASAP7_75t_SL g2380 ( 
.A(n_2164),
.B(n_166),
.Y(n_2380)
);

OAI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_1992),
.A2(n_166),
.B(n_169),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2047),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2029),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_1995),
.B(n_174),
.Y(n_2384)
);

AOI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2000),
.A2(n_175),
.B(n_176),
.Y(n_2385)
);

OAI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2094),
.A2(n_176),
.B(n_177),
.Y(n_2386)
);

OAI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_1969),
.A2(n_177),
.B(n_178),
.Y(n_2387)
);

BUFx2_ASAP7_75t_L g2388 ( 
.A(n_2273),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2152),
.B(n_177),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2309),
.B(n_178),
.Y(n_2390)
);

OAI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2211),
.A2(n_178),
.B(n_179),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2059),
.B(n_222),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2286),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2029),
.Y(n_2394)
);

BUFx4_ASAP7_75t_SL g2395 ( 
.A(n_2063),
.Y(n_2395)
);

OR2x6_ASAP7_75t_SL g2396 ( 
.A(n_2075),
.B(n_179),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2000),
.A2(n_179),
.B(n_180),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2043),
.B(n_181),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2029),
.Y(n_2399)
);

BUFx10_ASAP7_75t_L g2400 ( 
.A(n_2286),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2044),
.Y(n_2401)
);

AO31x2_ASAP7_75t_L g2402 ( 
.A1(n_2198),
.A2(n_184),
.A3(n_182),
.B(n_183),
.Y(n_2402)
);

AOI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_2209),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2044),
.Y(n_2404)
);

NAND3x1_ASAP7_75t_L g2405 ( 
.A(n_2139),
.B(n_185),
.C(n_186),
.Y(n_2405)
);

AO21x2_ASAP7_75t_L g2406 ( 
.A1(n_2190),
.A2(n_186),
.B(n_187),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_2061),
.B(n_223),
.Y(n_2407)
);

AOI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2004),
.A2(n_186),
.B(n_187),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2200),
.B(n_187),
.Y(n_2409)
);

BUFx4_ASAP7_75t_SL g2410 ( 
.A(n_2127),
.Y(n_2410)
);

AO32x2_ASAP7_75t_L g2411 ( 
.A1(n_2173),
.A2(n_190),
.A3(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_2411)
);

A2O1A1Ixp33_ASAP7_75t_L g2412 ( 
.A1(n_2061),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2004),
.A2(n_190),
.B(n_192),
.Y(n_2413)
);

BUFx12f_ASAP7_75t_L g2414 ( 
.A(n_2202),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2044),
.Y(n_2415)
);

NOR2xp67_ASAP7_75t_L g2416 ( 
.A(n_1989),
.B(n_192),
.Y(n_2416)
);

A2O1A1Ixp33_ASAP7_75t_L g2417 ( 
.A1(n_2062),
.A2(n_196),
.B(n_193),
.C(n_195),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2085),
.Y(n_2418)
);

A2O1A1Ixp33_ASAP7_75t_L g2419 ( 
.A1(n_2062),
.A2(n_197),
.B(n_193),
.C(n_196),
.Y(n_2419)
);

INVxp67_ASAP7_75t_L g2420 ( 
.A(n_1973),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_SL g2421 ( 
.A1(n_2192),
.A2(n_2317),
.B(n_2286),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2317),
.B(n_196),
.Y(n_2422)
);

BUFx4f_ASAP7_75t_SL g2423 ( 
.A(n_1980),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2317),
.Y(n_2424)
);

AOI21xp5_ASAP7_75t_L g2425 ( 
.A1(n_2057),
.A2(n_2053),
.B(n_2050),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2215),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2085),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2218),
.B(n_2363),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2085),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2231),
.B(n_197),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2091),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2055),
.A2(n_198),
.B(n_199),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2026),
.B(n_198),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2074),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2012),
.B(n_200),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2239),
.B(n_201),
.Y(n_2436)
);

BUFx8_ASAP7_75t_L g2437 ( 
.A(n_2208),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2192),
.Y(n_2438)
);

NOR2xp67_ASAP7_75t_SL g2439 ( 
.A(n_2023),
.B(n_202),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_2091),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2256),
.B(n_2264),
.Y(n_2441)
);

AOI211x1_ASAP7_75t_L g2442 ( 
.A1(n_2170),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_2442)
);

INVxp67_ASAP7_75t_L g2443 ( 
.A(n_2230),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2091),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2289),
.B(n_205),
.Y(n_2445)
);

AO31x2_ASAP7_75t_L g2446 ( 
.A1(n_2199),
.A2(n_2079),
.A3(n_2197),
.B(n_2196),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_SL g2447 ( 
.A1(n_2129),
.A2(n_206),
.B(n_207),
.Y(n_2447)
);

NAND2xp33_ASAP7_75t_R g2448 ( 
.A(n_2033),
.B(n_206),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2310),
.B(n_206),
.Y(n_2449)
);

OAI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2312),
.A2(n_208),
.B(n_209),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2314),
.B(n_209),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2258),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2315),
.B(n_210),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2316),
.B(n_211),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2129),
.Y(n_2455)
);

AOI22xp5_ASAP7_75t_L g2456 ( 
.A1(n_2182),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2129),
.B(n_212),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2326),
.B(n_214),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2341),
.B(n_215),
.Y(n_2459)
);

BUFx3_ASAP7_75t_L g2460 ( 
.A(n_2148),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2342),
.B(n_216),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2148),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2189),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2463)
);

NOR2xp67_ASAP7_75t_SL g2464 ( 
.A(n_2019),
.B(n_217),
.Y(n_2464)
);

AO32x2_ASAP7_75t_L g2465 ( 
.A1(n_2173),
.A2(n_220),
.A3(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_2465)
);

AOI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2066),
.A2(n_218),
.B(n_219),
.Y(n_2466)
);

OAI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2354),
.A2(n_219),
.B(n_220),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2080),
.B(n_2131),
.Y(n_2468)
);

AO31x2_ASAP7_75t_L g2469 ( 
.A1(n_2076),
.A2(n_2161),
.A3(n_2167),
.B(n_2162),
.Y(n_2469)
);

BUFx12f_ASAP7_75t_L g2470 ( 
.A(n_2146),
.Y(n_2470)
);

AOI221x1_ASAP7_75t_L g2471 ( 
.A1(n_2182),
.A2(n_221),
.B1(n_225),
.B2(n_224),
.C(n_226),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_R g2472 ( 
.A(n_2147),
.B(n_227),
.Y(n_2472)
);

AOI211x1_ASAP7_75t_L g2473 ( 
.A1(n_2171),
.A2(n_233),
.B(n_230),
.C(n_232),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2212),
.B(n_233),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2359),
.B(n_234),
.Y(n_2475)
);

AO32x2_ASAP7_75t_L g2476 ( 
.A1(n_2160),
.A2(n_238),
.A3(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_2476)
);

INVx6_ASAP7_75t_SL g2477 ( 
.A(n_1978),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2086),
.Y(n_2478)
);

NOR2x1_ASAP7_75t_SL g2479 ( 
.A(n_2166),
.B(n_238),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_1978),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2220),
.B(n_241),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2074),
.A2(n_2168),
.B1(n_2328),
.B2(n_2177),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_1991),
.B(n_243),
.Y(n_2483)
);

AO32x2_ASAP7_75t_L g2484 ( 
.A1(n_2159),
.A2(n_246),
.A3(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_2484)
);

OR2x6_ASAP7_75t_L g2485 ( 
.A(n_2020),
.B(n_248),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_1971),
.B(n_250),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_1991),
.B(n_250),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_1991),
.B(n_251),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2110),
.B(n_2124),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2087),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_1978),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2003),
.B(n_252),
.Y(n_2492)
);

AOI221xp5_ASAP7_75t_L g2493 ( 
.A1(n_2165),
.A2(n_256),
.B1(n_259),
.B2(n_255),
.C(n_258),
.Y(n_2493)
);

BUFx3_ASAP7_75t_L g2494 ( 
.A(n_2115),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2038),
.B(n_253),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2003),
.B(n_259),
.Y(n_2496)
);

CKINVDCx14_ASAP7_75t_R g2497 ( 
.A(n_2154),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2158),
.A2(n_2194),
.B1(n_2049),
.B2(n_2064),
.Y(n_2498)
);

A2O1A1Ixp33_ASAP7_75t_L g2499 ( 
.A1(n_2114),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_2499)
);

AND2x4_ASAP7_75t_L g2500 ( 
.A(n_2041),
.B(n_2008),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2003),
.B(n_266),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2207),
.B(n_268),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2092),
.Y(n_2503)
);

A2O1A1Ixp33_ASAP7_75t_L g2504 ( 
.A1(n_2114),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2098),
.Y(n_2505)
);

BUFx4f_ASAP7_75t_L g2506 ( 
.A(n_2067),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2068),
.B(n_273),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2244),
.B(n_273),
.Y(n_2508)
);

INVxp67_ASAP7_75t_SL g2509 ( 
.A(n_2288),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2034),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_1971),
.B(n_274),
.Y(n_2511)
);

AOI21xp5_ASAP7_75t_SL g2512 ( 
.A1(n_2201),
.A2(n_275),
.B(n_276),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2193),
.A2(n_281),
.B1(n_277),
.B2(n_279),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2065),
.Y(n_2514)
);

INVx1_ASAP7_75t_SL g2515 ( 
.A(n_2306),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2319),
.B(n_283),
.Y(n_2516)
);

BUFx12f_ASAP7_75t_L g2517 ( 
.A(n_2071),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2347),
.B(n_284),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2081),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2099),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2355),
.B(n_285),
.Y(n_2521)
);

BUFx2_ASAP7_75t_L g2522 ( 
.A(n_2035),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_1985),
.B(n_286),
.Y(n_2523)
);

HB1xp67_ASAP7_75t_L g2524 ( 
.A(n_2191),
.Y(n_2524)
);

BUFx3_ASAP7_75t_L g2525 ( 
.A(n_2058),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2117),
.B(n_289),
.Y(n_2526)
);

AND2x4_ASAP7_75t_L g2527 ( 
.A(n_2153),
.B(n_291),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_2217),
.B(n_294),
.Y(n_2528)
);

BUFx2_ASAP7_75t_R g2529 ( 
.A(n_1990),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2104),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2073),
.B(n_2100),
.Y(n_2531)
);

OAI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2112),
.Y(n_2532)
);

CKINVDCx11_ASAP7_75t_R g2533 ( 
.A(n_2151),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2060),
.B(n_300),
.Y(n_2534)
);

CKINVDCx6p67_ASAP7_75t_R g2535 ( 
.A(n_2135),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2018),
.B(n_301),
.Y(n_2536)
);

O2A1O1Ixp5_ASAP7_75t_SL g2537 ( 
.A1(n_2088),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_2537)
);

A2O1A1Ixp33_ASAP7_75t_L g2538 ( 
.A1(n_2116),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_2538)
);

OAI22x1_ASAP7_75t_L g2539 ( 
.A1(n_2195),
.A2(n_312),
.B1(n_313),
.B2(n_311),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_R g2540 ( 
.A(n_2194),
.B(n_837),
.Y(n_2540)
);

AND3x2_ASAP7_75t_L g2541 ( 
.A(n_1988),
.B(n_319),
.C(n_309),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_1999),
.B(n_315),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2101),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2105),
.Y(n_2544)
);

BUFx2_ASAP7_75t_SL g2545 ( 
.A(n_2014),
.Y(n_2545)
);

AO21x1_ASAP7_75t_L g2546 ( 
.A1(n_2203),
.A2(n_315),
.B(n_316),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2001),
.B(n_2002),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2178),
.B(n_2179),
.Y(n_2548)
);

OAI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2126),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2109),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2078),
.A2(n_320),
.B1(n_317),
.B2(n_318),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2005),
.B(n_2013),
.Y(n_2552)
);

INVx2_ASAP7_75t_SL g2553 ( 
.A(n_1994),
.Y(n_2553)
);

INVx4_ASAP7_75t_L g2554 ( 
.A(n_2180),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2111),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_R g2556 ( 
.A(n_2217),
.B(n_836),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2118),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2313),
.B(n_323),
.Y(n_2558)
);

BUFx2_ASAP7_75t_L g2559 ( 
.A(n_2101),
.Y(n_2559)
);

INVx4_ASAP7_75t_L g2560 ( 
.A(n_2185),
.Y(n_2560)
);

OAI21x1_ASAP7_75t_L g2561 ( 
.A1(n_2120),
.A2(n_2122),
.B(n_2121),
.Y(n_2561)
);

AO21x2_ASAP7_75t_L g2562 ( 
.A1(n_2128),
.A2(n_325),
.B(n_327),
.Y(n_2562)
);

NOR4xp25_ASAP7_75t_L g2563 ( 
.A(n_2181),
.B(n_330),
.C(n_328),
.D(n_329),
.Y(n_2563)
);

NAND2x1_ASAP7_75t_L g2564 ( 
.A(n_2132),
.B(n_329),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2313),
.B(n_330),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2072),
.Y(n_2566)
);

NAND3x1_ASAP7_75t_L g2567 ( 
.A(n_2143),
.B(n_2150),
.C(n_2149),
.Y(n_2567)
);

OAI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2082),
.A2(n_332),
.B(n_333),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2010),
.B(n_333),
.Y(n_2569)
);

AO21x2_ASAP7_75t_L g2570 ( 
.A1(n_2130),
.A2(n_334),
.B(n_335),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2024),
.B(n_335),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2083),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_2572)
);

OAI22x1_ASAP7_75t_L g2573 ( 
.A1(n_2184),
.A2(n_341),
.B1(n_342),
.B2(n_340),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2040),
.B(n_339),
.Y(n_2574)
);

BUFx2_ASAP7_75t_R g2575 ( 
.A(n_2106),
.Y(n_2575)
);

AO32x2_ASAP7_75t_L g2576 ( 
.A1(n_2203),
.A2(n_343),
.A3(n_341),
.B1(n_342),
.B2(n_344),
.Y(n_2576)
);

OAI21x1_ASAP7_75t_L g2577 ( 
.A1(n_2141),
.A2(n_2145),
.B(n_2142),
.Y(n_2577)
);

NOR4xp25_ASAP7_75t_L g2578 ( 
.A(n_2186),
.B(n_356),
.C(n_354),
.D(n_355),
.Y(n_2578)
);

OAI22xp5_ASAP7_75t_L g2579 ( 
.A1(n_2138),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2133),
.B(n_357),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2084),
.A2(n_357),
.B(n_358),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2188),
.B(n_360),
.Y(n_2582)
);

NAND2x1_ASAP7_75t_L g2583 ( 
.A(n_2183),
.B(n_363),
.Y(n_2583)
);

CKINVDCx5p33_ASAP7_75t_R g2584 ( 
.A(n_2022),
.Y(n_2584)
);

OR2x6_ASAP7_75t_L g2585 ( 
.A(n_2136),
.B(n_366),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2134),
.B(n_366),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2102),
.Y(n_2587)
);

AND3x4_ASAP7_75t_L g2588 ( 
.A(n_2077),
.B(n_367),
.C(n_368),
.Y(n_2588)
);

AO21x2_ASAP7_75t_L g2589 ( 
.A1(n_2155),
.A2(n_369),
.B(n_370),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2187),
.Y(n_2590)
);

OAI21xp33_ASAP7_75t_L g2591 ( 
.A1(n_2205),
.A2(n_370),
.B(n_371),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2157),
.Y(n_2592)
);

NOR4xp25_ASAP7_75t_L g2593 ( 
.A(n_2371),
.B(n_2210),
.C(n_2214),
.D(n_2213),
.Y(n_2593)
);

AO31x2_ASAP7_75t_L g2594 ( 
.A1(n_2119),
.A2(n_373),
.A3(n_371),
.B(n_372),
.Y(n_2594)
);

NAND3xp33_ASAP7_75t_L g2595 ( 
.A(n_2072),
.B(n_372),
.C(n_373),
.Y(n_2595)
);

AO31x2_ASAP7_75t_L g2596 ( 
.A1(n_2090),
.A2(n_2095),
.A3(n_2097),
.B(n_2096),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_1997),
.B(n_1998),
.Y(n_2597)
);

INVxp67_ASAP7_75t_L g2598 ( 
.A(n_1979),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2185),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2216),
.Y(n_2600)
);

NAND2xp33_ASAP7_75t_L g2601 ( 
.A(n_2318),
.B(n_377),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2206),
.A2(n_379),
.B(n_380),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_SL g2603 ( 
.A(n_2225),
.B(n_381),
.C(n_382),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2169),
.A2(n_384),
.B1(n_381),
.B2(n_383),
.Y(n_2604)
);

INVx2_ASAP7_75t_SL g2605 ( 
.A(n_1986),
.Y(n_2605)
);

AOI21xp5_ASAP7_75t_SL g2606 ( 
.A1(n_2174),
.A2(n_383),
.B(n_384),
.Y(n_2606)
);

AOI211x1_ASAP7_75t_L g2607 ( 
.A1(n_2176),
.A2(n_387),
.B(n_385),
.C(n_386),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2219),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_SL g2609 ( 
.A(n_2318),
.B(n_385),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2027),
.B(n_388),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2045),
.B(n_390),
.Y(n_2611)
);

INVx1_ASAP7_75t_SL g2612 ( 
.A(n_1970),
.Y(n_2612)
);

NAND2x1p5_ASAP7_75t_L g2613 ( 
.A(n_2016),
.B(n_392),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_1987),
.B(n_392),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2322),
.B(n_393),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2140),
.B(n_394),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_1982),
.Y(n_2617)
);

BUFx3_ASAP7_75t_L g2618 ( 
.A(n_1996),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2322),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2069),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2123),
.B(n_396),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2015),
.B(n_397),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2221),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2090),
.A2(n_399),
.B(n_400),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2222),
.Y(n_2625)
);

AO22x2_ASAP7_75t_L g2626 ( 
.A1(n_2175),
.A2(n_408),
.B1(n_404),
.B2(n_406),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2021),
.B(n_409),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2223),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2030),
.B(n_409),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2325),
.B(n_410),
.Y(n_2630)
);

BUFx12f_ASAP7_75t_L g2631 ( 
.A(n_2226),
.Y(n_2631)
);

OAI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2224),
.A2(n_414),
.B1(n_411),
.B2(n_412),
.Y(n_2632)
);

CKINVDCx20_ASAP7_75t_R g2633 ( 
.A(n_2017),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2325),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2227),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2144),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2329),
.B(n_419),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2228),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2125),
.A2(n_420),
.B(n_421),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2031),
.B(n_420),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2229),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2144),
.Y(n_2642)
);

O2A1O1Ixp33_ASAP7_75t_L g2643 ( 
.A1(n_2232),
.A2(n_424),
.B(n_422),
.C(n_423),
.Y(n_2643)
);

AOI21xp33_ASAP7_75t_L g2644 ( 
.A1(n_2032),
.A2(n_2007),
.B(n_2006),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2246),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2137),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2233),
.B(n_423),
.Y(n_2647)
);

NOR2xp67_ASAP7_75t_L g2648 ( 
.A(n_1974),
.B(n_424),
.Y(n_2648)
);

NOR2xp67_ASAP7_75t_L g2649 ( 
.A(n_1975),
.B(n_425),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2234),
.Y(n_2650)
);

AO32x2_ASAP7_75t_L g2651 ( 
.A1(n_2107),
.A2(n_428),
.A3(n_426),
.B1(n_427),
.B2(n_429),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2235),
.B(n_429),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_1983),
.Y(n_2653)
);

INVxp67_ASAP7_75t_SL g2654 ( 
.A(n_2236),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2070),
.B(n_430),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_1972),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2028),
.B(n_433),
.Y(n_2657)
);

BUFx3_ASAP7_75t_L g2658 ( 
.A(n_2009),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2237),
.B(n_434),
.Y(n_2659)
);

O2A1O1Ixp33_ASAP7_75t_L g2660 ( 
.A1(n_2238),
.A2(n_438),
.B(n_435),
.C(n_437),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2036),
.A2(n_437),
.B(n_439),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2240),
.Y(n_2662)
);

INVx5_ASAP7_75t_L g2663 ( 
.A(n_2329),
.Y(n_2663)
);

OR2x2_ASAP7_75t_L g2664 ( 
.A(n_1977),
.B(n_2370),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2241),
.Y(n_2665)
);

INVx1_ASAP7_75t_SL g2666 ( 
.A(n_2249),
.Y(n_2666)
);

CKINVDCx20_ASAP7_75t_R g2667 ( 
.A(n_2255),
.Y(n_2667)
);

OR2x2_ASAP7_75t_L g2668 ( 
.A(n_2369),
.B(n_444),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2242),
.B(n_445),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2257),
.Y(n_2670)
);

AO32x2_ASAP7_75t_L g2671 ( 
.A1(n_2107),
.A2(n_449),
.A3(n_446),
.B1(n_447),
.B2(n_450),
.Y(n_2671)
);

A2O1A1Ixp33_ASAP7_75t_L g2672 ( 
.A1(n_2330),
.A2(n_450),
.B(n_446),
.C(n_447),
.Y(n_2672)
);

BUFx5_ASAP7_75t_L g2673 ( 
.A(n_2330),
.Y(n_2673)
);

OAI21x1_ASAP7_75t_L g2674 ( 
.A1(n_1984),
.A2(n_451),
.B(n_452),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2243),
.Y(n_2675)
);

OAI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2037),
.A2(n_453),
.B(n_456),
.Y(n_2676)
);

O2A1O1Ixp33_ASAP7_75t_L g2677 ( 
.A1(n_2245),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_2677)
);

A2O1A1Ixp33_ASAP7_75t_L g2678 ( 
.A1(n_2331),
.A2(n_463),
.B(n_461),
.C(n_462),
.Y(n_2678)
);

BUFx12f_ASAP7_75t_L g2679 ( 
.A(n_2259),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2247),
.B(n_462),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2331),
.A2(n_467),
.B1(n_464),
.B2(n_466),
.Y(n_2681)
);

AOI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_2108),
.A2(n_467),
.B(n_468),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2113),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_SL g2684 ( 
.A(n_2333),
.B(n_469),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2248),
.Y(n_2685)
);

NOR2x1_ASAP7_75t_L g2686 ( 
.A(n_2250),
.B(n_471),
.Y(n_2686)
);

AOI21xp33_ASAP7_75t_L g2687 ( 
.A1(n_2046),
.A2(n_472),
.B(n_473),
.Y(n_2687)
);

OAI22x1_ASAP7_75t_L g2688 ( 
.A1(n_2251),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2108),
.A2(n_475),
.B(n_477),
.Y(n_2689)
);

BUFx10_ASAP7_75t_L g2690 ( 
.A(n_2265),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_L g2691 ( 
.A(n_2056),
.Y(n_2691)
);

AOI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2333),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2252),
.B(n_478),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2253),
.Y(n_2694)
);

A2O1A1Ixp33_ASAP7_75t_L g2695 ( 
.A1(n_2337),
.A2(n_481),
.B(n_479),
.C(n_480),
.Y(n_2695)
);

OAI21x1_ASAP7_75t_SL g2696 ( 
.A1(n_2337),
.A2(n_483),
.B(n_485),
.Y(n_2696)
);

NOR3xp33_ASAP7_75t_L g2697 ( 
.A(n_2266),
.B(n_486),
.C(n_487),
.Y(n_2697)
);

AOI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_2048),
.A2(n_2051),
.B(n_2025),
.Y(n_2698)
);

INVxp67_ASAP7_75t_SL g2699 ( 
.A(n_2254),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2345),
.Y(n_2700)
);

NAND2xp33_ASAP7_75t_L g2701 ( 
.A(n_2345),
.B(n_2346),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2260),
.B(n_490),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2261),
.B(n_2262),
.Y(n_2703)
);

A2O1A1Ixp33_ASAP7_75t_L g2704 ( 
.A1(n_2346),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_2704)
);

NAND3xp33_ASAP7_75t_L g2705 ( 
.A(n_2269),
.B(n_491),
.C(n_492),
.Y(n_2705)
);

CKINVDCx14_ASAP7_75t_R g2706 ( 
.A(n_2287),
.Y(n_2706)
);

BUFx3_ASAP7_75t_L g2707 ( 
.A(n_2292),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2263),
.B(n_493),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2042),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2267),
.B(n_493),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2268),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2089),
.B(n_494),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2349),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2270),
.B(n_495),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2295),
.Y(n_2715)
);

AOI21xp33_ASAP7_75t_L g2716 ( 
.A1(n_2011),
.A2(n_496),
.B(n_497),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2271),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2272),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2274),
.Y(n_2719)
);

INVx1_ASAP7_75t_SL g2720 ( 
.A(n_2297),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2352),
.A2(n_498),
.B(n_499),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2275),
.B(n_499),
.Y(n_2722)
);

OAI21x1_ASAP7_75t_L g2723 ( 
.A1(n_2425),
.A2(n_2277),
.B(n_2276),
.Y(n_2723)
);

AO21x2_ASAP7_75t_L g2724 ( 
.A1(n_2566),
.A2(n_2279),
.B(n_2278),
.Y(n_2724)
);

CKINVDCx16_ASAP7_75t_R g2725 ( 
.A(n_2472),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2457),
.Y(n_2726)
);

AO31x2_ASAP7_75t_L g2727 ( 
.A1(n_2566),
.A2(n_2368),
.A3(n_2352),
.B(n_2280),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2468),
.B(n_2281),
.Y(n_2728)
);

O2A1O1Ixp33_ASAP7_75t_SL g2729 ( 
.A1(n_2412),
.A2(n_2282),
.B(n_2284),
.C(n_2283),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2457),
.Y(n_2730)
);

AO31x2_ASAP7_75t_L g2731 ( 
.A1(n_2636),
.A2(n_2368),
.A3(n_2285),
.B(n_2291),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2554),
.B(n_2290),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2515),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2482),
.A2(n_2303),
.B1(n_2305),
.B2(n_2302),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2554),
.A2(n_2307),
.B1(n_2293),
.B2(n_2294),
.Y(n_2735)
);

INVx6_ASAP7_75t_L g2736 ( 
.A(n_2489),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2560),
.B(n_2296),
.Y(n_2737)
);

HB1xp67_ASAP7_75t_L g2738 ( 
.A(n_2393),
.Y(n_2738)
);

AO21x2_ASAP7_75t_L g2739 ( 
.A1(n_2636),
.A2(n_2299),
.B(n_2298),
.Y(n_2739)
);

AO31x2_ASAP7_75t_L g2740 ( 
.A1(n_2642),
.A2(n_2300),
.A3(n_2304),
.B(n_2301),
.Y(n_2740)
);

AO21x2_ASAP7_75t_L g2741 ( 
.A1(n_2642),
.A2(n_2311),
.B(n_2308),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2375),
.Y(n_2742)
);

INVxp67_ASAP7_75t_SL g2743 ( 
.A(n_2374),
.Y(n_2743)
);

INVx3_ASAP7_75t_L g2744 ( 
.A(n_2379),
.Y(n_2744)
);

INVx2_ASAP7_75t_SL g2745 ( 
.A(n_2395),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2389),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2402),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2375),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2382),
.Y(n_2749)
);

BUFx2_ASAP7_75t_SL g2750 ( 
.A(n_2633),
.Y(n_2750)
);

HB1xp67_ASAP7_75t_L g2751 ( 
.A(n_2480),
.Y(n_2751)
);

AOI21x1_ASAP7_75t_L g2752 ( 
.A1(n_2543),
.A2(n_2321),
.B(n_2320),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2560),
.B(n_2324),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2426),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_2410),
.Y(n_2755)
);

NOR2xp67_ASAP7_75t_L g2756 ( 
.A(n_2663),
.B(n_2327),
.Y(n_2756)
);

OAI21x1_ASAP7_75t_L g2757 ( 
.A1(n_2561),
.A2(n_2334),
.B(n_2332),
.Y(n_2757)
);

OAI221xp5_ASAP7_75t_L g2758 ( 
.A1(n_2498),
.A2(n_2448),
.B1(n_2684),
.B2(n_2552),
.C(n_2547),
.Y(n_2758)
);

OAI21x1_ASAP7_75t_L g2759 ( 
.A1(n_2567),
.A2(n_2336),
.B(n_2335),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2426),
.Y(n_2760)
);

AOI221xp5_ASAP7_75t_L g2761 ( 
.A1(n_2376),
.A2(n_2340),
.B1(n_2343),
.B2(n_2339),
.C(n_2338),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_2533),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2555),
.B(n_2344),
.Y(n_2763)
);

O2A1O1Ixp33_ASAP7_75t_SL g2764 ( 
.A1(n_2417),
.A2(n_2348),
.B(n_2351),
.C(n_2350),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2557),
.B(n_2353),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2402),
.Y(n_2766)
);

AO21x2_ASAP7_75t_L g2767 ( 
.A1(n_2700),
.A2(n_2357),
.B(n_2356),
.Y(n_2767)
);

AOI21xp33_ASAP7_75t_SL g2768 ( 
.A1(n_2588),
.A2(n_2360),
.B(n_2358),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2421),
.A2(n_2362),
.B(n_2361),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2440),
.Y(n_2770)
);

OAI21x1_ASAP7_75t_L g2771 ( 
.A1(n_2713),
.A2(n_2365),
.B(n_2364),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2590),
.B(n_2366),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2440),
.Y(n_2773)
);

OAI21x1_ASAP7_75t_L g2774 ( 
.A1(n_2577),
.A2(n_2367),
.B(n_2052),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2402),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_2701),
.A2(n_2039),
.B1(n_1981),
.B2(n_502),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2379),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2460),
.B(n_500),
.Y(n_2778)
);

INVx4_ASAP7_75t_L g2779 ( 
.A(n_2440),
.Y(n_2779)
);

HB1xp67_ASAP7_75t_L g2780 ( 
.A(n_2444),
.Y(n_2780)
);

OAI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2373),
.A2(n_501),
.B(n_502),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2372),
.Y(n_2782)
);

OA21x2_ASAP7_75t_L g2783 ( 
.A1(n_2471),
.A2(n_503),
.B(n_504),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2590),
.B(n_503),
.Y(n_2784)
);

CKINVDCx11_ASAP7_75t_R g2785 ( 
.A(n_2535),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2601),
.A2(n_2523),
.B(n_2407),
.Y(n_2786)
);

BUFx12f_ASAP7_75t_L g2787 ( 
.A(n_2489),
.Y(n_2787)
);

O2A1O1Ixp33_ASAP7_75t_L g2788 ( 
.A1(n_2443),
.A2(n_507),
.B(n_504),
.C(n_505),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2383),
.B(n_507),
.Y(n_2789)
);

INVx3_ASAP7_75t_L g2790 ( 
.A(n_2400),
.Y(n_2790)
);

OR2x6_ASAP7_75t_L g2791 ( 
.A(n_2388),
.B(n_508),
.Y(n_2791)
);

AO21x2_ASAP7_75t_L g2792 ( 
.A1(n_2696),
.A2(n_508),
.B(n_509),
.Y(n_2792)
);

NAND3xp33_ASAP7_75t_L g2793 ( 
.A(n_2607),
.B(n_509),
.C(n_510),
.Y(n_2793)
);

INVx2_ASAP7_75t_SL g2794 ( 
.A(n_2423),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2399),
.B(n_510),
.Y(n_2795)
);

OAI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2428),
.A2(n_512),
.B(n_514),
.Y(n_2796)
);

BUFx3_ASAP7_75t_L g2797 ( 
.A(n_2494),
.Y(n_2797)
);

O2A1O1Ixp33_ASAP7_75t_SL g2798 ( 
.A1(n_2419),
.A2(n_518),
.B(n_516),
.C(n_517),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2506),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_2799)
);

INVxp33_ASAP7_75t_L g2800 ( 
.A(n_2506),
.Y(n_2800)
);

BUFx2_ASAP7_75t_SL g2801 ( 
.A(n_2667),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2478),
.Y(n_2802)
);

AND2x2_ASAP7_75t_SL g2803 ( 
.A(n_2424),
.B(n_521),
.Y(n_2803)
);

INVx4_ASAP7_75t_L g2804 ( 
.A(n_2444),
.Y(n_2804)
);

NAND3xp33_ASAP7_75t_L g2805 ( 
.A(n_2493),
.B(n_525),
.C(n_526),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_SL g2806 ( 
.A1(n_2540),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_2806)
);

CKINVDCx12_ASAP7_75t_R g2807 ( 
.A(n_2485),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2444),
.Y(n_2808)
);

CKINVDCx20_ASAP7_75t_R g2809 ( 
.A(n_2437),
.Y(n_2809)
);

OR2x2_ASAP7_75t_L g2810 ( 
.A(n_2390),
.B(n_527),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2490),
.Y(n_2811)
);

NAND3xp33_ASAP7_75t_L g2812 ( 
.A(n_2473),
.B(n_530),
.C(n_531),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_SL g2813 ( 
.A(n_2663),
.B(n_531),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_2529),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2548),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2524),
.A2(n_535),
.B1(n_532),
.B2(n_533),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2582),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2668),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2404),
.B(n_535),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2697),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2503),
.Y(n_2821)
);

AO21x2_ASAP7_75t_L g2822 ( 
.A1(n_2546),
.A2(n_539),
.B(n_540),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2505),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2409),
.B(n_539),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2707),
.A2(n_543),
.B1(n_540),
.B2(n_542),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2415),
.B(n_544),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2514),
.Y(n_2827)
);

BUFx2_ASAP7_75t_SL g2828 ( 
.A(n_2416),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_2437),
.Y(n_2829)
);

NAND2x1p5_ASAP7_75t_L g2830 ( 
.A(n_2510),
.B(n_545),
.Y(n_2830)
);

OR2x2_ASAP7_75t_L g2831 ( 
.A(n_2509),
.B(n_548),
.Y(n_2831)
);

OAI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2441),
.A2(n_2381),
.B(n_2377),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2474),
.B(n_548),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2400),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_2477),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2714),
.Y(n_2836)
);

BUFx12f_ASAP7_75t_L g2837 ( 
.A(n_2485),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2452),
.B(n_2497),
.Y(n_2838)
);

AO21x2_ASAP7_75t_L g2839 ( 
.A1(n_2391),
.A2(n_552),
.B(n_553),
.Y(n_2839)
);

OAI21x1_ASAP7_75t_SL g2840 ( 
.A1(n_2380),
.A2(n_552),
.B(n_553),
.Y(n_2840)
);

OAI221xp5_ASAP7_75t_L g2841 ( 
.A1(n_2456),
.A2(n_557),
.B1(n_554),
.B2(n_555),
.C(n_558),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2594),
.Y(n_2842)
);

O2A1O1Ixp33_ASAP7_75t_SL g2843 ( 
.A1(n_2634),
.A2(n_557),
.B(n_554),
.C(n_555),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2455),
.Y(n_2844)
);

AOI22x1_ASAP7_75t_L g2845 ( 
.A1(n_2688),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2586),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2527),
.Y(n_2847)
);

INVx3_ASAP7_75t_L g2848 ( 
.A(n_2455),
.Y(n_2848)
);

INVx3_ASAP7_75t_L g2849 ( 
.A(n_2455),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2418),
.B(n_561),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2462),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2527),
.Y(n_2852)
);

BUFx2_ASAP7_75t_L g2853 ( 
.A(n_2477),
.Y(n_2853)
);

INVx4_ASAP7_75t_L g2854 ( 
.A(n_2462),
.Y(n_2854)
);

AO21x1_ASAP7_75t_L g2855 ( 
.A1(n_2528),
.A2(n_562),
.B(n_563),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2491),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2618),
.B(n_563),
.Y(n_2857)
);

AOI221xp5_ASAP7_75t_L g2858 ( 
.A1(n_2434),
.A2(n_567),
.B1(n_564),
.B2(n_565),
.C(n_568),
.Y(n_2858)
);

BUFx12f_ASAP7_75t_L g2859 ( 
.A(n_2584),
.Y(n_2859)
);

INVx6_ASAP7_75t_L g2860 ( 
.A(n_2631),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2663),
.B(n_567),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2545),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2715),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_2863)
);

AOI22xp33_ASAP7_75t_L g2864 ( 
.A1(n_2712),
.A2(n_2556),
.B1(n_2703),
.B2(n_2603),
.Y(n_2864)
);

INVxp67_ASAP7_75t_L g2865 ( 
.A(n_2396),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2427),
.B(n_573),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2598),
.B(n_574),
.Y(n_2867)
);

OR2x2_ASAP7_75t_L g2868 ( 
.A(n_2481),
.B(n_575),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2656),
.Y(n_2869)
);

NAND3xp33_ASAP7_75t_SL g2870 ( 
.A(n_2670),
.B(n_577),
.C(n_578),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2442),
.Y(n_2871)
);

INVx2_ASAP7_75t_SL g2872 ( 
.A(n_2690),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2517),
.B(n_578),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2398),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2392),
.A2(n_581),
.B(n_582),
.Y(n_2875)
);

INVx3_ASAP7_75t_L g2876 ( 
.A(n_2438),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2626),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2626),
.Y(n_2878)
);

INVx1_ASAP7_75t_SL g2879 ( 
.A(n_2491),
.Y(n_2879)
);

AOI22xp33_ASAP7_75t_L g2880 ( 
.A1(n_2712),
.A2(n_586),
.B1(n_583),
.B2(n_584),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2429),
.B(n_586),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2679),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2612),
.B(n_587),
.Y(n_2883)
);

OAI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2559),
.A2(n_591),
.B1(n_588),
.B2(n_589),
.Y(n_2884)
);

BUFx2_ASAP7_75t_L g2885 ( 
.A(n_2709),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2394),
.B(n_592),
.Y(n_2886)
);

NAND2x1p5_ASAP7_75t_L g2887 ( 
.A(n_2522),
.B(n_595),
.Y(n_2887)
);

A2O1A1Ixp33_ASAP7_75t_L g2888 ( 
.A1(n_2385),
.A2(n_598),
.B(n_596),
.C(n_597),
.Y(n_2888)
);

INVxp67_ASAP7_75t_SL g2889 ( 
.A(n_2401),
.Y(n_2889)
);

INVx1_ASAP7_75t_SL g2890 ( 
.A(n_2438),
.Y(n_2890)
);

OAI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2387),
.A2(n_596),
.B(n_597),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_SL g2892 ( 
.A1(n_2479),
.A2(n_599),
.B(n_600),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2536),
.Y(n_2893)
);

OAI22xp5_ASAP7_75t_L g2894 ( 
.A1(n_2438),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2610),
.Y(n_2895)
);

AOI22xp33_ASAP7_75t_SL g2896 ( 
.A1(n_2706),
.A2(n_604),
.B1(n_601),
.B2(n_603),
.Y(n_2896)
);

AOI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_2587),
.A2(n_609),
.B1(n_606),
.B2(n_608),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2596),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2614),
.Y(n_2899)
);

OAI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2463),
.A2(n_610),
.B1(n_606),
.B2(n_608),
.Y(n_2900)
);

A2O1A1Ixp33_ASAP7_75t_L g2901 ( 
.A1(n_2397),
.A2(n_614),
.B(n_612),
.C(n_613),
.Y(n_2901)
);

HB1xp67_ASAP7_75t_L g2902 ( 
.A(n_2508),
.Y(n_2902)
);

NAND3xp33_ASAP7_75t_L g2903 ( 
.A(n_2537),
.B(n_613),
.C(n_614),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2518),
.B(n_615),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2575),
.B(n_615),
.Y(n_2905)
);

AOI22x1_ASAP7_75t_L g2906 ( 
.A1(n_2539),
.A2(n_619),
.B1(n_617),
.B2(n_618),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2674),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_2422),
.B(n_2525),
.Y(n_2908)
);

BUFx3_ASAP7_75t_L g2909 ( 
.A(n_2414),
.Y(n_2909)
);

AOI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2486),
.A2(n_617),
.B(n_618),
.Y(n_2910)
);

INVx3_ASAP7_75t_SL g2911 ( 
.A(n_2585),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2431),
.B(n_620),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2544),
.A2(n_2620),
.B1(n_2495),
.B2(n_2470),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2519),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2406),
.Y(n_2915)
);

OAI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2450),
.A2(n_621),
.B(n_622),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2605),
.B(n_623),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_2495),
.Y(n_2918)
);

NOR2xp67_ASAP7_75t_L g2919 ( 
.A(n_2595),
.B(n_624),
.Y(n_2919)
);

AO31x2_ASAP7_75t_L g2920 ( 
.A1(n_2499),
.A2(n_627),
.A3(n_625),
.B(n_626),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2469),
.B(n_626),
.Y(n_2921)
);

O2A1O1Ixp33_ASAP7_75t_SL g2922 ( 
.A1(n_2672),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_2922)
);

OAI21x1_ASAP7_75t_SL g2923 ( 
.A1(n_2721),
.A2(n_628),
.B(n_629),
.Y(n_2923)
);

INVxp33_ASAP7_75t_L g2924 ( 
.A(n_2439),
.Y(n_2924)
);

OR2x6_ASAP7_75t_L g2925 ( 
.A(n_2447),
.B(n_630),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2406),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2469),
.B(n_631),
.Y(n_2927)
);

BUFx2_ASAP7_75t_SL g2928 ( 
.A(n_2648),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2585),
.B(n_632),
.Y(n_2929)
);

NAND2x1p5_ASAP7_75t_L g2930 ( 
.A(n_2464),
.B(n_845),
.Y(n_2930)
);

BUFx3_ASAP7_75t_L g2931 ( 
.A(n_2658),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2511),
.A2(n_636),
.B(n_637),
.Y(n_2932)
);

AO21x2_ASAP7_75t_L g2933 ( 
.A1(n_2467),
.A2(n_639),
.B(n_640),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2520),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2616),
.Y(n_2935)
);

INVx2_ASAP7_75t_SL g2936 ( 
.A(n_2690),
.Y(n_2936)
);

BUFx3_ASAP7_75t_L g2937 ( 
.A(n_2553),
.Y(n_2937)
);

INVxp67_ASAP7_75t_SL g2938 ( 
.A(n_2673),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2569),
.Y(n_2939)
);

NAND2x1p5_ASAP7_75t_L g2940 ( 
.A(n_2645),
.B(n_641),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2573),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2530),
.Y(n_2942)
);

CKINVDCx20_ASAP7_75t_R g2943 ( 
.A(n_2420),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2433),
.Y(n_2944)
);

AO21x2_ASAP7_75t_L g2945 ( 
.A1(n_2408),
.A2(n_845),
.B(n_644),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2550),
.Y(n_2946)
);

CKINVDCx16_ASAP7_75t_R g2947 ( 
.A(n_2569),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2710),
.Y(n_2948)
);

AOI21xp33_ASAP7_75t_L g2949 ( 
.A1(n_2583),
.A2(n_650),
.B(n_651),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2657),
.Y(n_2950)
);

AOI21x1_ASAP7_75t_L g2951 ( 
.A1(n_2558),
.A2(n_650),
.B(n_651),
.Y(n_2951)
);

AOI21x1_ASAP7_75t_L g2952 ( 
.A1(n_2565),
.A2(n_652),
.B(n_653),
.Y(n_2952)
);

AO21x2_ASAP7_75t_L g2953 ( 
.A1(n_2413),
.A2(n_844),
.B(n_653),
.Y(n_2953)
);

INVxp67_ASAP7_75t_SL g2954 ( 
.A(n_2673),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2544),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_2955)
);

AOI22xp5_ASAP7_75t_L g2956 ( 
.A1(n_2531),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_2956)
);

BUFx3_ASAP7_75t_L g2957 ( 
.A(n_2617),
.Y(n_2957)
);

A2O1A1Ixp33_ASAP7_75t_SL g2958 ( 
.A1(n_2384),
.A2(n_2386),
.B(n_2435),
.C(n_2676),
.Y(n_2958)
);

CKINVDCx11_ASAP7_75t_R g2959 ( 
.A(n_2666),
.Y(n_2959)
);

OAI21x1_ASAP7_75t_SL g2960 ( 
.A1(n_2682),
.A2(n_660),
.B(n_661),
.Y(n_2960)
);

INVx3_ASAP7_75t_SL g2961 ( 
.A(n_2653),
.Y(n_2961)
);

INVx1_ASAP7_75t_SL g2962 ( 
.A(n_2673),
.Y(n_2962)
);

HB1xp67_ASAP7_75t_L g2963 ( 
.A(n_2483),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2657),
.Y(n_2964)
);

NAND3xp33_ASAP7_75t_L g2965 ( 
.A(n_2705),
.B(n_662),
.C(n_663),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2596),
.Y(n_2966)
);

O2A1O1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2716),
.A2(n_665),
.B(n_663),
.C(n_664),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2534),
.B(n_667),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2686),
.A2(n_671),
.B1(n_668),
.B2(n_670),
.Y(n_2969)
);

OAI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2602),
.A2(n_673),
.B(n_674),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_L g2971 ( 
.A1(n_2564),
.A2(n_673),
.B(n_675),
.Y(n_2971)
);

OR2x2_ASAP7_75t_L g2972 ( 
.A(n_2516),
.B(n_680),
.Y(n_2972)
);

INVx4_ASAP7_75t_L g2973 ( 
.A(n_2673),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2720),
.A2(n_683),
.B1(n_680),
.B2(n_681),
.Y(n_2974)
);

AOI221xp5_ASAP7_75t_SL g2975 ( 
.A1(n_2504),
.A2(n_681),
.B1(n_683),
.B2(n_685),
.C(n_687),
.Y(n_2975)
);

A2O1A1Ixp33_ASAP7_75t_L g2976 ( 
.A1(n_2624),
.A2(n_688),
.B(n_685),
.C(n_687),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2487),
.Y(n_2977)
);

BUFx3_ASAP7_75t_L g2978 ( 
.A(n_2500),
.Y(n_2978)
);

AO32x2_ASAP7_75t_L g2979 ( 
.A1(n_2549),
.A2(n_689),
.A3(n_690),
.B1(n_691),
.B2(n_692),
.Y(n_2979)
);

AO21x2_ASAP7_75t_L g2980 ( 
.A1(n_2689),
.A2(n_690),
.B(n_691),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2446),
.B(n_692),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2655),
.Y(n_2982)
);

NAND2x1p5_ASAP7_75t_L g2983 ( 
.A(n_2609),
.B(n_843),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2378),
.B(n_693),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2600),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_2985)
);

BUFx12f_ASAP7_75t_L g2986 ( 
.A(n_2500),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2673),
.B(n_695),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2621),
.Y(n_2988)
);

AOI22xp33_ASAP7_75t_L g2989 ( 
.A1(n_2608),
.A2(n_701),
.B1(n_697),
.B2(n_699),
.Y(n_2989)
);

AOI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2403),
.A2(n_703),
.B1(n_701),
.B2(n_702),
.Y(n_2990)
);

HB1xp67_ASAP7_75t_L g2991 ( 
.A(n_2488),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2492),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2623),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_2993)
);

AOI22xp33_ASAP7_75t_L g2994 ( 
.A1(n_2625),
.A2(n_704),
.B1(n_705),
.B2(n_706),
.Y(n_2994)
);

O2A1O1Ixp33_ASAP7_75t_SL g2995 ( 
.A1(n_2678),
.A2(n_707),
.B(n_708),
.C(n_709),
.Y(n_2995)
);

OAI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2619),
.A2(n_708),
.B1(n_709),
.B2(n_710),
.Y(n_2996)
);

BUFx3_ASAP7_75t_L g2997 ( 
.A(n_2613),
.Y(n_2997)
);

BUFx6f_ASAP7_75t_L g2998 ( 
.A(n_2691),
.Y(n_2998)
);

INVxp67_ASAP7_75t_L g2999 ( 
.A(n_2597),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2649),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2580),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2532),
.A2(n_711),
.B(n_712),
.Y(n_3002)
);

AOI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2615),
.A2(n_712),
.B(n_713),
.Y(n_3003)
);

OAI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2466),
.A2(n_713),
.B(n_714),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2521),
.B(n_715),
.Y(n_3005)
);

OR2x2_ASAP7_75t_L g3006 ( 
.A(n_2496),
.B(n_715),
.Y(n_3006)
);

NOR2x1_ASAP7_75t_SL g3007 ( 
.A(n_2630),
.B(n_716),
.Y(n_3007)
);

AOI21xp33_ASAP7_75t_SL g3008 ( 
.A1(n_2637),
.A2(n_716),
.B(n_717),
.Y(n_3008)
);

NOR3xp33_ASAP7_75t_L g3009 ( 
.A(n_2644),
.B(n_717),
.C(n_718),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2592),
.B(n_719),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2432),
.A2(n_720),
.B(n_721),
.Y(n_3011)
);

OAI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2692),
.A2(n_2599),
.B1(n_2681),
.B2(n_2695),
.Y(n_3012)
);

INVx3_ASAP7_75t_SL g3013 ( 
.A(n_2664),
.Y(n_3013)
);

AOI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2579),
.A2(n_2513),
.B1(n_2502),
.B2(n_2405),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2691),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_2512),
.Y(n_3016)
);

AOI21x1_ASAP7_75t_L g3017 ( 
.A1(n_2475),
.A2(n_720),
.B(n_722),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2628),
.B(n_722),
.Y(n_3018)
);

INVxp67_ASAP7_75t_L g3019 ( 
.A(n_2501),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2704),
.A2(n_723),
.B1(n_724),
.B2(n_725),
.Y(n_3020)
);

CKINVDCx14_ASAP7_75t_R g3021 ( 
.A(n_2551),
.Y(n_3021)
);

AO32x2_ASAP7_75t_L g3022 ( 
.A1(n_2604),
.A2(n_723),
.A3(n_724),
.B1(n_725),
.B2(n_726),
.Y(n_3022)
);

BUFx12f_ASAP7_75t_L g3023 ( 
.A(n_2691),
.Y(n_3023)
);

AO21x2_ASAP7_75t_L g3024 ( 
.A1(n_2568),
.A2(n_843),
.B(n_727),
.Y(n_3024)
);

BUFx3_ASAP7_75t_L g3025 ( 
.A(n_2635),
.Y(n_3025)
);

CKINVDCx11_ASAP7_75t_R g3026 ( 
.A(n_2694),
.Y(n_3026)
);

OAI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2430),
.A2(n_728),
.B(n_729),
.Y(n_3027)
);

AO21x1_ASAP7_75t_L g3028 ( 
.A1(n_2639),
.A2(n_729),
.B(n_730),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2638),
.A2(n_730),
.B1(n_731),
.B2(n_732),
.Y(n_3029)
);

INVx4_ASAP7_75t_SL g3030 ( 
.A(n_2641),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2646),
.B(n_731),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2650),
.B(n_732),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2662),
.B(n_733),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2665),
.A2(n_733),
.B1(n_734),
.B2(n_735),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2675),
.B(n_2685),
.Y(n_3035)
);

HB1xp67_ASAP7_75t_L g3036 ( 
.A(n_2507),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2717),
.A2(n_734),
.B1(n_736),
.B2(n_737),
.Y(n_3037)
);

AO31x2_ASAP7_75t_L g3038 ( 
.A1(n_2538),
.A2(n_736),
.A3(n_737),
.B(n_738),
.Y(n_3038)
);

INVxp67_ASAP7_75t_L g3039 ( 
.A(n_2622),
.Y(n_3039)
);

BUFx2_ASAP7_75t_L g3040 ( 
.A(n_2654),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2647),
.Y(n_3041)
);

A2O1A1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_2581),
.A2(n_741),
.B(n_742),
.C(n_744),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2652),
.Y(n_3043)
);

OAI221xp5_ASAP7_75t_L g3044 ( 
.A1(n_2593),
.A2(n_842),
.B1(n_745),
.B2(n_746),
.C(n_747),
.Y(n_3044)
);

OA21x2_ASAP7_75t_L g3045 ( 
.A1(n_2591),
.A2(n_744),
.B(n_745),
.Y(n_3045)
);

CKINVDCx9p33_ASAP7_75t_R g3046 ( 
.A(n_2882),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2754),
.Y(n_3047)
);

INVx3_ASAP7_75t_L g3048 ( 
.A(n_2973),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2747),
.Y(n_3049)
);

AND2x4_ASAP7_75t_L g3050 ( 
.A(n_3030),
.B(n_2779),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2760),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2973),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2766),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2775),
.Y(n_3054)
);

HB1xp67_ASAP7_75t_L g3055 ( 
.A(n_2733),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2842),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2824),
.B(n_2476),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2802),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2811),
.Y(n_3059)
);

INVx3_ASAP7_75t_L g3060 ( 
.A(n_2744),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2898),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2898),
.Y(n_3062)
);

INVx2_ASAP7_75t_SL g3063 ( 
.A(n_2745),
.Y(n_3063)
);

HB1xp67_ASAP7_75t_L g3064 ( 
.A(n_2902),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2966),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2821),
.Y(n_3066)
);

INVx5_ASAP7_75t_L g3067 ( 
.A(n_2791),
.Y(n_3067)
);

INVx1_ASAP7_75t_SL g3068 ( 
.A(n_2862),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2823),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2827),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2966),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2915),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2833),
.B(n_2476),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2914),
.Y(n_3074)
);

OAI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2758),
.A2(n_2947),
.B1(n_2925),
.B2(n_2734),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2758),
.A2(n_2699),
.B1(n_2719),
.B2(n_2718),
.Y(n_3076)
);

INVx2_ASAP7_75t_SL g3077 ( 
.A(n_2829),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2934),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2942),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2746),
.B(n_2563),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2946),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2846),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2742),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_2911),
.B(n_2541),
.Y(n_3084)
);

NOR2x1_ASAP7_75t_R g3085 ( 
.A(n_2785),
.B(n_2659),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2871),
.Y(n_3086)
);

INVx4_ASAP7_75t_L g3087 ( 
.A(n_2797),
.Y(n_3087)
);

INVx3_ASAP7_75t_L g3088 ( 
.A(n_2744),
.Y(n_3088)
);

INVx2_ASAP7_75t_SL g3089 ( 
.A(n_2909),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2818),
.Y(n_3090)
);

INVx3_ASAP7_75t_L g3091 ( 
.A(n_2777),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2782),
.B(n_2578),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2836),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2748),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2749),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_3021),
.A2(n_2711),
.B1(n_2632),
.B2(n_2683),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2869),
.Y(n_3097)
);

OR2x2_ASAP7_75t_L g3098 ( 
.A(n_3013),
.B(n_2810),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2784),
.Y(n_3099)
);

CKINVDCx8_ASAP7_75t_R g3100 ( 
.A(n_2725),
.Y(n_3100)
);

INVx3_ASAP7_75t_L g3101 ( 
.A(n_2777),
.Y(n_3101)
);

AOI211xp5_ASAP7_75t_L g3102 ( 
.A1(n_2865),
.A2(n_2687),
.B(n_2698),
.C(n_2606),
.Y(n_3102)
);

BUFx3_ASAP7_75t_L g3103 ( 
.A(n_2809),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2738),
.Y(n_3104)
);

OR2x2_ASAP7_75t_L g3105 ( 
.A(n_2868),
.B(n_2436),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2790),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_2904),
.B(n_2476),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2944),
.B(n_2445),
.Y(n_3108)
);

BUFx6f_ASAP7_75t_L g3109 ( 
.A(n_2869),
.Y(n_3109)
);

CKINVDCx20_ASAP7_75t_R g3110 ( 
.A(n_2755),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2784),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2831),
.Y(n_3112)
);

HB1xp67_ASAP7_75t_L g3113 ( 
.A(n_2751),
.Y(n_3113)
);

HB1xp67_ASAP7_75t_L g3114 ( 
.A(n_2885),
.Y(n_3114)
);

BUFx6f_ASAP7_75t_L g3115 ( 
.A(n_2869),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2817),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_2743),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2988),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2941),
.Y(n_3119)
);

CKINVDCx5p33_ASAP7_75t_R g3120 ( 
.A(n_2762),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2877),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2878),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2728),
.B(n_2411),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2837),
.B(n_2627),
.Y(n_3124)
);

OR2x2_ASAP7_75t_L g3125 ( 
.A(n_2918),
.B(n_2449),
.Y(n_3125)
);

BUFx2_ASAP7_75t_L g3126 ( 
.A(n_3023),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2935),
.Y(n_3127)
);

HB1xp67_ASAP7_75t_L g3128 ( 
.A(n_2791),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2982),
.Y(n_3129)
);

BUFx2_ASAP7_75t_L g3130 ( 
.A(n_2787),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2790),
.Y(n_3131)
);

INVx4_ASAP7_75t_L g3132 ( 
.A(n_2834),
.Y(n_3132)
);

HB1xp67_ASAP7_75t_L g3133 ( 
.A(n_2791),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_2859),
.Y(n_3134)
);

HB1xp67_ASAP7_75t_L g3135 ( 
.A(n_3040),
.Y(n_3135)
);

A2O1A1Ixp33_ASAP7_75t_L g3136 ( 
.A1(n_2768),
.A2(n_2677),
.B(n_2643),
.C(n_2660),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2803),
.A2(n_2572),
.B1(n_2722),
.B2(n_2702),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2834),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2948),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3010),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3010),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2999),
.B(n_2874),
.Y(n_3142)
);

BUFx2_ASAP7_75t_L g3143 ( 
.A(n_2986),
.Y(n_3143)
);

INVx3_ASAP7_75t_L g3144 ( 
.A(n_2779),
.Y(n_3144)
);

CKINVDCx20_ASAP7_75t_R g3145 ( 
.A(n_2807),
.Y(n_3145)
);

INVx2_ASAP7_75t_SL g3146 ( 
.A(n_2794),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3031),
.Y(n_3147)
);

CKINVDCx5p33_ASAP7_75t_R g3148 ( 
.A(n_2814),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3031),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2968),
.B(n_2411),
.Y(n_3150)
);

INVx2_ASAP7_75t_SL g3151 ( 
.A(n_2860),
.Y(n_3151)
);

INVx3_ASAP7_75t_L g3152 ( 
.A(n_2804),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2886),
.Y(n_3153)
);

AOI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_2786),
.A2(n_2453),
.B(n_2451),
.Y(n_3154)
);

BUFx2_ASAP7_75t_L g3155 ( 
.A(n_2931),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2929),
.B(n_2411),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2789),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2950),
.B(n_2454),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_2726),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2789),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2939),
.B(n_2458),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2795),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2795),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2819),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_2730),
.Y(n_3165)
);

BUFx3_ASAP7_75t_L g3166 ( 
.A(n_2961),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2819),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2826),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2826),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_2804),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_2801),
.B(n_2465),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_SL g3172 ( 
.A1(n_2813),
.A2(n_2589),
.B1(n_2570),
.B2(n_2562),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2926),
.Y(n_3173)
);

HB1xp67_ASAP7_75t_L g3174 ( 
.A(n_2770),
.Y(n_3174)
);

BUFx3_ASAP7_75t_L g3175 ( 
.A(n_2937),
.Y(n_3175)
);

BUFx6f_ASAP7_75t_L g3176 ( 
.A(n_2773),
.Y(n_3176)
);

OAI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_2925),
.A2(n_2708),
.B1(n_2693),
.B2(n_2680),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3005),
.B(n_2465),
.Y(n_3178)
);

NAND2xp33_ASAP7_75t_SL g3179 ( 
.A(n_2800),
.B(n_2864),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2850),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2964),
.B(n_2459),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_2854),
.Y(n_3182)
);

OR2x2_ASAP7_75t_L g3183 ( 
.A(n_2908),
.B(n_2461),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2921),
.Y(n_3184)
);

HB1xp67_ASAP7_75t_L g3185 ( 
.A(n_2780),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2927),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2927),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2850),
.Y(n_3188)
);

BUFx2_ASAP7_75t_L g3189 ( 
.A(n_2854),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_2750),
.B(n_2669),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2866),
.Y(n_3191)
);

CKINVDCx5p33_ASAP7_75t_R g3192 ( 
.A(n_2860),
.Y(n_3192)
);

INVx2_ASAP7_75t_SL g3193 ( 
.A(n_2957),
.Y(n_3193)
);

INVxp67_ASAP7_75t_L g3194 ( 
.A(n_2838),
.Y(n_3194)
);

INVx3_ASAP7_75t_L g3195 ( 
.A(n_2773),
.Y(n_3195)
);

INVx1_ASAP7_75t_SL g3196 ( 
.A(n_2959),
.Y(n_3196)
);

BUFx2_ASAP7_75t_L g3197 ( 
.A(n_3015),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2866),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2778),
.B(n_2465),
.Y(n_3199)
);

A2O1A1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_2768),
.A2(n_2769),
.B(n_2916),
.C(n_2781),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_2773),
.Y(n_3201)
);

INVx3_ASAP7_75t_L g3202 ( 
.A(n_2732),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2881),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2881),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2912),
.Y(n_3205)
);

CKINVDCx14_ASAP7_75t_R g3206 ( 
.A(n_2943),
.Y(n_3206)
);

AO221x2_ASAP7_75t_L g3207 ( 
.A1(n_2884),
.A2(n_2576),
.B1(n_2671),
.B2(n_2651),
.C(n_2484),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2912),
.Y(n_3208)
);

HB1xp67_ASAP7_75t_L g3209 ( 
.A(n_2808),
.Y(n_3209)
);

BUFx12f_ASAP7_75t_L g3210 ( 
.A(n_3026),
.Y(n_3210)
);

BUFx6f_ASAP7_75t_L g3211 ( 
.A(n_2998),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_3001),
.B(n_2526),
.Y(n_3212)
);

OAI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2805),
.A2(n_2661),
.B(n_2571),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3025),
.Y(n_3214)
);

INVxp67_ASAP7_75t_L g3215 ( 
.A(n_2828),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2981),
.Y(n_3216)
);

CKINVDCx11_ASAP7_75t_R g3217 ( 
.A(n_2835),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2893),
.B(n_2542),
.Y(n_3218)
);

INVx3_ASAP7_75t_L g3219 ( 
.A(n_2732),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2981),
.Y(n_3220)
);

OR2x2_ASAP7_75t_L g3221 ( 
.A(n_2978),
.B(n_2574),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3035),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3000),
.Y(n_3223)
);

AO21x2_ASAP7_75t_L g3224 ( 
.A1(n_2987),
.A2(n_2611),
.B(n_2629),
.Y(n_3224)
);

OR2x6_ASAP7_75t_L g3225 ( 
.A(n_2925),
.B(n_2640),
.Y(n_3225)
);

INVx3_ASAP7_75t_L g3226 ( 
.A(n_2737),
.Y(n_3226)
);

BUFx2_ASAP7_75t_SL g3227 ( 
.A(n_2872),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3036),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3033),
.Y(n_3229)
);

NAND3xp33_ASAP7_75t_L g3230 ( 
.A(n_2761),
.B(n_2484),
.C(n_2576),
.Y(n_3230)
);

INVxp67_ASAP7_75t_L g3231 ( 
.A(n_2857),
.Y(n_3231)
);

BUFx3_ASAP7_75t_L g3232 ( 
.A(n_2853),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3041),
.Y(n_3233)
);

AOI21x1_ASAP7_75t_L g3234 ( 
.A1(n_2919),
.A2(n_2671),
.B(n_2651),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3043),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_2778),
.B(n_2651),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2763),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2763),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2765),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2765),
.Y(n_3240)
);

INVx1_ASAP7_75t_SL g3241 ( 
.A(n_2736),
.Y(n_3241)
);

OAI21x1_ASAP7_75t_SL g3242 ( 
.A1(n_3007),
.A2(n_2671),
.B(n_748),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2737),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2812),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2895),
.B(n_748),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2844),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2812),
.Y(n_3247)
);

O2A1O1Ixp5_ASAP7_75t_L g3248 ( 
.A1(n_2861),
.A2(n_749),
.B(n_750),
.C(n_751),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2772),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_2883),
.B(n_749),
.Y(n_3250)
);

BUFx2_ASAP7_75t_L g3251 ( 
.A(n_2936),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2772),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3017),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2899),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2847),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2852),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_2736),
.Y(n_3257)
);

OR2x6_ASAP7_75t_L g3258 ( 
.A(n_2928),
.B(n_750),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2851),
.Y(n_3259)
);

INVxp67_ASAP7_75t_L g3260 ( 
.A(n_2917),
.Y(n_3260)
);

BUFx3_ASAP7_75t_L g3261 ( 
.A(n_2876),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2867),
.B(n_751),
.Y(n_3262)
);

OA21x2_ASAP7_75t_L g3263 ( 
.A1(n_2907),
.A2(n_752),
.B(n_753),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2793),
.Y(n_3264)
);

CKINVDCx5p33_ASAP7_75t_R g3265 ( 
.A(n_2873),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_2963),
.B(n_2977),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2793),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2984),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2984),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_2997),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2920),
.Y(n_3271)
);

BUFx6f_ASAP7_75t_L g3272 ( 
.A(n_2848),
.Y(n_3272)
);

OR2x2_ASAP7_75t_L g3273 ( 
.A(n_2991),
.B(n_752),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2920),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2920),
.Y(n_3275)
);

INVx3_ASAP7_75t_L g3276 ( 
.A(n_2753),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_2761),
.A2(n_755),
.B1(n_756),
.B2(n_757),
.Y(n_3277)
);

HB1xp67_ASAP7_75t_L g3278 ( 
.A(n_2856),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3038),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3038),
.Y(n_3280)
);

BUFx2_ASAP7_75t_SL g3281 ( 
.A(n_2756),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_2890),
.Y(n_3282)
);

OAI21xp33_ASAP7_75t_L g3283 ( 
.A1(n_2813),
.A2(n_758),
.B(n_760),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3038),
.Y(n_3284)
);

BUFx2_ASAP7_75t_L g3285 ( 
.A(n_3030),
.Y(n_3285)
);

INVx2_ASAP7_75t_SL g3286 ( 
.A(n_2887),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2884),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3019),
.B(n_763),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2945),
.Y(n_3289)
);

BUFx6f_ASAP7_75t_L g3290 ( 
.A(n_2848),
.Y(n_3290)
);

BUFx2_ASAP7_75t_L g3291 ( 
.A(n_2876),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2945),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2992),
.B(n_842),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_2890),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2938),
.Y(n_3295)
);

INVx3_ASAP7_75t_L g3296 ( 
.A(n_2753),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2954),
.Y(n_3297)
);

BUFx2_ASAP7_75t_L g3298 ( 
.A(n_2849),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2962),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2962),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2822),
.Y(n_3301)
);

BUFx4f_ASAP7_75t_SL g3302 ( 
.A(n_2849),
.Y(n_3302)
);

OAI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2805),
.A2(n_764),
.B(n_766),
.Y(n_3303)
);

OR2x2_ASAP7_75t_L g3304 ( 
.A(n_2879),
.B(n_764),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2792),
.Y(n_3305)
);

INVxp67_ASAP7_75t_SL g3306 ( 
.A(n_2889),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2792),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_2806),
.B(n_841),
.Y(n_3308)
);

HB1xp67_ASAP7_75t_L g3309 ( 
.A(n_2879),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3039),
.B(n_2972),
.Y(n_3310)
);

HB1xp67_ASAP7_75t_L g3311 ( 
.A(n_3117),
.Y(n_3311)
);

NAND2xp33_ASAP7_75t_SL g3312 ( 
.A(n_3285),
.B(n_2913),
.Y(n_3312)
);

INVx1_ASAP7_75t_SL g3313 ( 
.A(n_3046),
.Y(n_3313)
);

INVxp67_ASAP7_75t_L g3314 ( 
.A(n_3113),
.Y(n_3314)
);

OR2x6_ASAP7_75t_L g3315 ( 
.A(n_3281),
.B(n_3087),
.Y(n_3315)
);

NAND2xp33_ASAP7_75t_R g3316 ( 
.A(n_3192),
.B(n_2905),
.Y(n_3316)
);

CKINVDCx5p33_ASAP7_75t_R g3317 ( 
.A(n_3110),
.Y(n_3317)
);

INVxp67_ASAP7_75t_L g3318 ( 
.A(n_3227),
.Y(n_3318)
);

INVxp67_ASAP7_75t_L g3319 ( 
.A(n_3114),
.Y(n_3319)
);

OR2x6_ASAP7_75t_L g3320 ( 
.A(n_3087),
.B(n_2830),
.Y(n_3320)
);

INVx8_ASAP7_75t_L g3321 ( 
.A(n_3210),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3058),
.Y(n_3322)
);

AND2x4_ASAP7_75t_L g3323 ( 
.A(n_3132),
.B(n_2756),
.Y(n_3323)
);

NAND2xp33_ASAP7_75t_R g3324 ( 
.A(n_3258),
.B(n_3016),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_R g3325 ( 
.A(n_3206),
.B(n_2870),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_R g3326 ( 
.A(n_3145),
.B(n_2752),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_R g3327 ( 
.A(n_3100),
.B(n_2951),
.Y(n_3327)
);

NOR2xp33_ASAP7_75t_R g3328 ( 
.A(n_3120),
.B(n_2952),
.Y(n_3328)
);

NAND2xp33_ASAP7_75t_R g3329 ( 
.A(n_3258),
.B(n_2783),
.Y(n_3329)
);

AND2x4_ASAP7_75t_L g3330 ( 
.A(n_3132),
.B(n_3067),
.Y(n_3330)
);

XNOR2xp5_ASAP7_75t_L g3331 ( 
.A(n_3148),
.B(n_2896),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3266),
.B(n_2767),
.Y(n_3332)
);

AND2x6_ASAP7_75t_L g3333 ( 
.A(n_3050),
.B(n_2956),
.Y(n_3333)
);

AND2x4_ASAP7_75t_L g3334 ( 
.A(n_3067),
.B(n_2796),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3082),
.Y(n_3335)
);

CKINVDCx5p33_ASAP7_75t_R g3336 ( 
.A(n_3103),
.Y(n_3336)
);

CKINVDCx20_ASAP7_75t_R g3337 ( 
.A(n_3217),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3059),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3118),
.B(n_2832),
.Y(n_3339)
);

BUFx3_ASAP7_75t_L g3340 ( 
.A(n_3166),
.Y(n_3340)
);

BUFx10_ASAP7_75t_L g3341 ( 
.A(n_3089),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3127),
.B(n_3129),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3090),
.Y(n_3343)
);

INVxp67_ASAP7_75t_L g3344 ( 
.A(n_3064),
.Y(n_3344)
);

INVxp67_ASAP7_75t_L g3345 ( 
.A(n_3098),
.Y(n_3345)
);

NAND2xp33_ASAP7_75t_R g3346 ( 
.A(n_3126),
.B(n_2783),
.Y(n_3346)
);

BUFx10_ASAP7_75t_L g3347 ( 
.A(n_3077),
.Y(n_3347)
);

AND2x4_ASAP7_75t_L g3348 ( 
.A(n_3067),
.B(n_2796),
.Y(n_3348)
);

CKINVDCx8_ASAP7_75t_R g3349 ( 
.A(n_3130),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3093),
.Y(n_3350)
);

XOR2x2_ASAP7_75t_SL g3351 ( 
.A(n_3075),
.B(n_2940),
.Y(n_3351)
);

OR2x6_ASAP7_75t_L g3352 ( 
.A(n_3050),
.B(n_3143),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_R g3353 ( 
.A(n_3134),
.B(n_3003),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3222),
.B(n_2767),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3310),
.B(n_2724),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3066),
.Y(n_3356)
);

XNOR2xp5_ASAP7_75t_L g3357 ( 
.A(n_3196),
.B(n_2924),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_R g3358 ( 
.A(n_3063),
.B(n_768),
.Y(n_3358)
);

XNOR2xp5_ASAP7_75t_L g3359 ( 
.A(n_3265),
.B(n_2894),
.Y(n_3359)
);

BUFx3_ASAP7_75t_L g3360 ( 
.A(n_3175),
.Y(n_3360)
);

AND2x4_ASAP7_75t_L g3361 ( 
.A(n_3189),
.B(n_3197),
.Y(n_3361)
);

INVxp67_ASAP7_75t_L g3362 ( 
.A(n_3155),
.Y(n_3362)
);

NOR2xp33_ASAP7_75t_R g3363 ( 
.A(n_3151),
.B(n_768),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3139),
.B(n_2724),
.Y(n_3364)
);

INVxp67_ASAP7_75t_L g3365 ( 
.A(n_3104),
.Y(n_3365)
);

NAND2xp33_ASAP7_75t_R g3366 ( 
.A(n_3251),
.B(n_3045),
.Y(n_3366)
);

XNOR2xp5_ASAP7_75t_L g3367 ( 
.A(n_3068),
.B(n_2894),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3144),
.B(n_2975),
.Y(n_3368)
);

CKINVDCx5p33_ASAP7_75t_R g3369 ( 
.A(n_3146),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_3194),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3112),
.B(n_3079),
.Y(n_3371)
);

AND2x4_ASAP7_75t_L g3372 ( 
.A(n_3144),
.B(n_2727),
.Y(n_3372)
);

XOR2xp5_ASAP7_75t_L g3373 ( 
.A(n_3190),
.B(n_3105),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3116),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_3152),
.B(n_2975),
.Y(n_3375)
);

NAND2xp33_ASAP7_75t_R g3376 ( 
.A(n_3084),
.B(n_769),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3233),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_R g3378 ( 
.A(n_3179),
.B(n_771),
.Y(n_3378)
);

NAND2xp33_ASAP7_75t_R g3379 ( 
.A(n_3308),
.B(n_771),
.Y(n_3379)
);

INVxp67_ASAP7_75t_L g3380 ( 
.A(n_3135),
.Y(n_3380)
);

INVx8_ASAP7_75t_L g3381 ( 
.A(n_3152),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_R g3382 ( 
.A(n_3270),
.B(n_773),
.Y(n_3382)
);

OR2x6_ASAP7_75t_L g3383 ( 
.A(n_3286),
.B(n_2840),
.Y(n_3383)
);

INVxp67_ASAP7_75t_L g3384 ( 
.A(n_3055),
.Y(n_3384)
);

NAND2xp33_ASAP7_75t_R g3385 ( 
.A(n_3170),
.B(n_774),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_R g3386 ( 
.A(n_3193),
.B(n_774),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3235),
.Y(n_3387)
);

CKINVDCx11_ASAP7_75t_R g3388 ( 
.A(n_3232),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3254),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3081),
.B(n_2832),
.Y(n_3390)
);

NAND2xp33_ASAP7_75t_R g3391 ( 
.A(n_3170),
.B(n_775),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_R g3392 ( 
.A(n_3182),
.B(n_775),
.Y(n_3392)
);

AND2x4_ASAP7_75t_L g3393 ( 
.A(n_3182),
.B(n_2727),
.Y(n_3393)
);

XNOR2xp5_ASAP7_75t_L g3394 ( 
.A(n_3250),
.B(n_2956),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3069),
.B(n_3018),
.Y(n_3395)
);

XNOR2xp5_ASAP7_75t_L g3396 ( 
.A(n_3128),
.B(n_2930),
.Y(n_3396)
);

AND2x4_ASAP7_75t_L g3397 ( 
.A(n_3060),
.B(n_3088),
.Y(n_3397)
);

AND2x4_ASAP7_75t_L g3398 ( 
.A(n_3060),
.B(n_3088),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3070),
.B(n_3032),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3074),
.B(n_2739),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3078),
.Y(n_3401)
);

INVxp67_ASAP7_75t_L g3402 ( 
.A(n_3174),
.Y(n_3402)
);

XNOR2xp5_ASAP7_75t_L g3403 ( 
.A(n_3133),
.B(n_3231),
.Y(n_3403)
);

OR2x6_ASAP7_75t_L g3404 ( 
.A(n_3225),
.B(n_2769),
.Y(n_3404)
);

XOR2xp5_ASAP7_75t_L g3405 ( 
.A(n_3183),
.B(n_3006),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_R g3406 ( 
.A(n_3302),
.B(n_776),
.Y(n_3406)
);

NOR2xp33_ASAP7_75t_R g3407 ( 
.A(n_3048),
.B(n_777),
.Y(n_3407)
);

OR2x6_ASAP7_75t_L g3408 ( 
.A(n_3225),
.B(n_2892),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_R g3409 ( 
.A(n_3048),
.B(n_777),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_R g3410 ( 
.A(n_3052),
.B(n_778),
.Y(n_3410)
);

HB1xp67_ASAP7_75t_L g3411 ( 
.A(n_3278),
.Y(n_3411)
);

AND2x4_ASAP7_75t_L g3412 ( 
.A(n_3091),
.B(n_3101),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_3047),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3228),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3171),
.B(n_2739),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_R g3416 ( 
.A(n_3052),
.B(n_778),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3142),
.Y(n_3417)
);

HB1xp67_ASAP7_75t_L g3418 ( 
.A(n_3185),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3156),
.B(n_2741),
.Y(n_3419)
);

NAND2xp33_ASAP7_75t_R g3420 ( 
.A(n_3091),
.B(n_779),
.Y(n_3420)
);

NAND2xp33_ASAP7_75t_R g3421 ( 
.A(n_3101),
.B(n_779),
.Y(n_3421)
);

NAND2xp33_ASAP7_75t_R g3422 ( 
.A(n_3106),
.B(n_780),
.Y(n_3422)
);

BUFx10_ASAP7_75t_L g3423 ( 
.A(n_3124),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3051),
.Y(n_3424)
);

AND2x4_ASAP7_75t_L g3425 ( 
.A(n_3106),
.B(n_2741),
.Y(n_3425)
);

NAND2xp33_ASAP7_75t_R g3426 ( 
.A(n_3131),
.B(n_780),
.Y(n_3426)
);

OR2x6_ASAP7_75t_L g3427 ( 
.A(n_3215),
.B(n_2916),
.Y(n_3427)
);

NAND2xp33_ASAP7_75t_R g3428 ( 
.A(n_3131),
.B(n_781),
.Y(n_3428)
);

NOR2xp33_ASAP7_75t_R g3429 ( 
.A(n_3138),
.B(n_782),
.Y(n_3429)
);

XNOR2xp5_ASAP7_75t_L g3430 ( 
.A(n_3262),
.B(n_2906),
.Y(n_3430)
);

AND2x4_ASAP7_75t_L g3431 ( 
.A(n_3138),
.B(n_2759),
.Y(n_3431)
);

OR2x6_ASAP7_75t_L g3432 ( 
.A(n_3283),
.B(n_2983),
.Y(n_3432)
);

INVx8_ASAP7_75t_L g3433 ( 
.A(n_3097),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3086),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3083),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_R g3436 ( 
.A(n_3109),
.B(n_782),
.Y(n_3436)
);

BUFx10_ASAP7_75t_L g3437 ( 
.A(n_3115),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_3214),
.B(n_2731),
.Y(n_3438)
);

NAND2xp33_ASAP7_75t_SL g3439 ( 
.A(n_3236),
.B(n_2839),
.Y(n_3439)
);

XNOR2xp5_ASAP7_75t_L g3440 ( 
.A(n_3293),
.B(n_2845),
.Y(n_3440)
);

NAND2xp33_ASAP7_75t_R g3441 ( 
.A(n_3199),
.B(n_783),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_R g3442 ( 
.A(n_3115),
.B(n_783),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3119),
.B(n_3223),
.Y(n_3443)
);

CKINVDCx5p33_ASAP7_75t_R g3444 ( 
.A(n_3257),
.Y(n_3444)
);

CKINVDCx5p33_ASAP7_75t_R g3445 ( 
.A(n_3241),
.Y(n_3445)
);

OR2x4_ASAP7_75t_L g3446 ( 
.A(n_3085),
.B(n_3044),
.Y(n_3446)
);

XOR2xp5_ASAP7_75t_L g3447 ( 
.A(n_3273),
.B(n_2990),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3237),
.B(n_3027),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_3123),
.B(n_2731),
.Y(n_3449)
);

NOR2xp33_ASAP7_75t_R g3450 ( 
.A(n_3115),
.B(n_784),
.Y(n_3450)
);

NAND2xp33_ASAP7_75t_R g3451 ( 
.A(n_3263),
.B(n_784),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_SL g3452 ( 
.A(n_3306),
.B(n_2841),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3209),
.B(n_2731),
.Y(n_3453)
);

AND2x4_ASAP7_75t_L g3454 ( 
.A(n_3261),
.B(n_3027),
.Y(n_3454)
);

XNOR2xp5_ASAP7_75t_L g3455 ( 
.A(n_3260),
.B(n_3096),
.Y(n_3455)
);

OR2x6_ASAP7_75t_L g3456 ( 
.A(n_3304),
.B(n_2781),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3200),
.B(n_2786),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3238),
.B(n_2990),
.Y(n_3458)
);

NAND2xp33_ASAP7_75t_R g3459 ( 
.A(n_3263),
.B(n_785),
.Y(n_3459)
);

INVxp67_ASAP7_75t_L g3460 ( 
.A(n_3288),
.Y(n_3460)
);

NAND2xp33_ASAP7_75t_R g3461 ( 
.A(n_3150),
.B(n_786),
.Y(n_3461)
);

AND2x4_ASAP7_75t_L g3462 ( 
.A(n_3202),
.B(n_2771),
.Y(n_3462)
);

CKINVDCx11_ASAP7_75t_R g3463 ( 
.A(n_3176),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3255),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3230),
.B(n_3008),
.Y(n_3465)
);

XNOR2xp5_ASAP7_75t_L g3466 ( 
.A(n_3102),
.B(n_3229),
.Y(n_3466)
);

BUFx3_ASAP7_75t_L g3467 ( 
.A(n_3291),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3256),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3121),
.Y(n_3469)
);

XNOR2xp5_ASAP7_75t_L g3470 ( 
.A(n_3178),
.B(n_3137),
.Y(n_3470)
);

BUFx2_ASAP7_75t_L g3471 ( 
.A(n_3282),
.Y(n_3471)
);

AND2x4_ASAP7_75t_L g3472 ( 
.A(n_3202),
.B(n_2774),
.Y(n_3472)
);

AND2x4_ASAP7_75t_L g3473 ( 
.A(n_3219),
.B(n_3226),
.Y(n_3473)
);

AND2x4_ASAP7_75t_L g3474 ( 
.A(n_3219),
.B(n_2723),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3095),
.B(n_2980),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_3294),
.Y(n_3476)
);

AND2x4_ASAP7_75t_L g3477 ( 
.A(n_3226),
.B(n_2757),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3073),
.B(n_3107),
.Y(n_3478)
);

XOR2xp5_ASAP7_75t_L g3479 ( 
.A(n_3125),
.B(n_2996),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3094),
.Y(n_3480)
);

CKINVDCx5p33_ASAP7_75t_R g3481 ( 
.A(n_3298),
.Y(n_3481)
);

NAND2xp33_ASAP7_75t_R g3482 ( 
.A(n_3057),
.B(n_786),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3239),
.B(n_2858),
.Y(n_3483)
);

AND2x4_ASAP7_75t_L g3484 ( 
.A(n_3243),
.B(n_2740),
.Y(n_3484)
);

NAND2xp33_ASAP7_75t_R g3485 ( 
.A(n_3243),
.B(n_787),
.Y(n_3485)
);

CKINVDCx5p33_ASAP7_75t_R g3486 ( 
.A(n_3276),
.Y(n_3486)
);

NAND2xp33_ASAP7_75t_R g3487 ( 
.A(n_3276),
.B(n_787),
.Y(n_3487)
);

OR2x6_ASAP7_75t_L g3488 ( 
.A(n_3303),
.B(n_2891),
.Y(n_3488)
);

CKINVDCx11_ASAP7_75t_R g3489 ( 
.A(n_3176),
.Y(n_3489)
);

INVxp33_ASAP7_75t_L g3490 ( 
.A(n_3272),
.Y(n_3490)
);

NAND2xp33_ASAP7_75t_R g3491 ( 
.A(n_3296),
.B(n_788),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3122),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3159),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3240),
.B(n_2858),
.Y(n_3494)
);

INVxp67_ASAP7_75t_L g3495 ( 
.A(n_3108),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3249),
.B(n_3014),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3252),
.B(n_3014),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3099),
.B(n_2839),
.Y(n_3498)
);

BUFx6f_ASAP7_75t_L g3499 ( 
.A(n_3211),
.Y(n_3499)
);

XNOR2xp5_ASAP7_75t_L g3500 ( 
.A(n_3177),
.B(n_2996),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_R g3501 ( 
.A(n_3296),
.B(n_789),
.Y(n_3501)
);

XNOR2xp5_ASAP7_75t_L g3502 ( 
.A(n_3165),
.B(n_3076),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3268),
.B(n_2980),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3269),
.B(n_2740),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3049),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3111),
.B(n_2933),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_R g3507 ( 
.A(n_3195),
.B(n_790),
.Y(n_3507)
);

NAND2xp33_ASAP7_75t_R g3508 ( 
.A(n_3287),
.B(n_790),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3246),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_R g3510 ( 
.A(n_3201),
.B(n_791),
.Y(n_3510)
);

INVxp67_ASAP7_75t_L g3511 ( 
.A(n_3245),
.Y(n_3511)
);

INVxp33_ASAP7_75t_SL g3512 ( 
.A(n_3309),
.Y(n_3512)
);

HB1xp67_ASAP7_75t_L g3513 ( 
.A(n_3295),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_R g3514 ( 
.A(n_3234),
.B(n_791),
.Y(n_3514)
);

OR2x6_ASAP7_75t_L g3515 ( 
.A(n_3242),
.B(n_2891),
.Y(n_3515)
);

NAND2xp33_ASAP7_75t_R g3516 ( 
.A(n_3221),
.B(n_792),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3259),
.B(n_2953),
.Y(n_3517)
);

HB1xp67_ASAP7_75t_L g3518 ( 
.A(n_3295),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_3290),
.Y(n_3519)
);

NAND2xp33_ASAP7_75t_R g3520 ( 
.A(n_3080),
.B(n_792),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3049),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3157),
.B(n_2933),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3053),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3160),
.B(n_2880),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3162),
.B(n_2958),
.Y(n_3525)
);

NAND2xp33_ASAP7_75t_SL g3526 ( 
.A(n_3244),
.B(n_2735),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_3290),
.Y(n_3527)
);

XOR2xp5_ASAP7_75t_L g3528 ( 
.A(n_3158),
.B(n_2799),
.Y(n_3528)
);

BUFx3_ASAP7_75t_L g3529 ( 
.A(n_3211),
.Y(n_3529)
);

AND2x4_ASAP7_75t_L g3530 ( 
.A(n_3153),
.B(n_2740),
.Y(n_3530)
);

INVxp67_ASAP7_75t_L g3531 ( 
.A(n_3161),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3505),
.Y(n_3532)
);

OR2x2_ASAP7_75t_L g3533 ( 
.A(n_3311),
.B(n_3072),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3478),
.B(n_3443),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3417),
.B(n_3470),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3521),
.Y(n_3536)
);

NAND3xp33_ASAP7_75t_L g3537 ( 
.A(n_3525),
.B(n_3092),
.C(n_3044),
.Y(n_3537)
);

AND2x4_ASAP7_75t_L g3538 ( 
.A(n_3372),
.B(n_3061),
.Y(n_3538)
);

AND2x4_ASAP7_75t_L g3539 ( 
.A(n_3393),
.B(n_3061),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3523),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3374),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3495),
.B(n_3355),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3513),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3471),
.B(n_3297),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3411),
.B(n_3297),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3380),
.B(n_3299),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3518),
.Y(n_3547)
);

BUFx3_ASAP7_75t_L g3548 ( 
.A(n_3360),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3332),
.B(n_3299),
.Y(n_3549)
);

AOI22xp5_ASAP7_75t_SL g3550 ( 
.A1(n_3313),
.A2(n_3247),
.B1(n_3267),
.B2(n_3264),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3413),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3377),
.Y(n_3552)
);

HB1xp67_ASAP7_75t_L g3553 ( 
.A(n_3418),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3318),
.B(n_3218),
.Y(n_3554)
);

NOR2x1p5_ASAP7_75t_L g3555 ( 
.A(n_3340),
.B(n_3330),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3414),
.B(n_3140),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3476),
.B(n_3300),
.Y(n_3557)
);

AOI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3500),
.A2(n_3009),
.B1(n_3277),
.B2(n_3207),
.Y(n_3558)
);

HB1xp67_ASAP7_75t_L g3559 ( 
.A(n_3402),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3319),
.B(n_3300),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3387),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3424),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3361),
.B(n_3184),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3435),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3531),
.B(n_3141),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3389),
.Y(n_3566)
);

OAI22xp5_ASAP7_75t_L g3567 ( 
.A1(n_3446),
.A2(n_2841),
.B1(n_3172),
.B2(n_2974),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3434),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3493),
.B(n_3147),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3335),
.Y(n_3570)
);

BUFx2_ASAP7_75t_L g3571 ( 
.A(n_3315),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3314),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3480),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3345),
.B(n_3184),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3344),
.B(n_3186),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3322),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3365),
.B(n_3149),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_L g3578 ( 
.A(n_3357),
.B(n_3212),
.Y(n_3578)
);

HB1xp67_ASAP7_75t_L g3579 ( 
.A(n_3467),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_3333),
.A2(n_3207),
.B1(n_3012),
.B2(n_3213),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_3499),
.Y(n_3581)
);

OAI221xp5_ASAP7_75t_L g3582 ( 
.A1(n_3520),
.A2(n_3136),
.B1(n_3181),
.B2(n_2776),
.C(n_3164),
.Y(n_3582)
);

HB1xp67_ASAP7_75t_L g3583 ( 
.A(n_3384),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3338),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3343),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3350),
.Y(n_3586)
);

INVx2_ASAP7_75t_SL g3587 ( 
.A(n_3341),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3342),
.Y(n_3588)
);

AND2x4_ASAP7_75t_L g3589 ( 
.A(n_3530),
.B(n_3062),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3333),
.A2(n_2900),
.B1(n_3020),
.B2(n_3012),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3371),
.Y(n_3591)
);

AND2x4_ASAP7_75t_L g3592 ( 
.A(n_3504),
.B(n_3062),
.Y(n_3592)
);

OR2x2_ASAP7_75t_L g3593 ( 
.A(n_3356),
.B(n_3072),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3496),
.B(n_3163),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3315),
.A2(n_3427),
.B1(n_3432),
.B2(n_3320),
.Y(n_3595)
);

OR2x2_ASAP7_75t_L g3596 ( 
.A(n_3401),
.B(n_3173),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3362),
.B(n_3186),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3469),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3354),
.B(n_3187),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3333),
.A2(n_3028),
.B1(n_2900),
.B2(n_3020),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3509),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3497),
.B(n_3167),
.Y(n_3602)
);

OR2x2_ASAP7_75t_L g3603 ( 
.A(n_3492),
.B(n_3173),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3464),
.Y(n_3604)
);

OR2x2_ASAP7_75t_L g3605 ( 
.A(n_3419),
.B(n_3053),
.Y(n_3605)
);

AND2x4_ASAP7_75t_L g3606 ( 
.A(n_3438),
.B(n_3065),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3468),
.Y(n_3607)
);

OAI21xp5_ASAP7_75t_SL g3608 ( 
.A1(n_3396),
.A2(n_3008),
.B(n_2949),
.Y(n_3608)
);

OR2x2_ASAP7_75t_L g3609 ( 
.A(n_3390),
.B(n_3449),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3400),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3364),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3397),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3339),
.B(n_3168),
.Y(n_3613)
);

INVxp67_ASAP7_75t_L g3614 ( 
.A(n_3385),
.Y(n_3614)
);

OR2x2_ASAP7_75t_L g3615 ( 
.A(n_3352),
.B(n_3054),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3398),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3522),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3403),
.B(n_3473),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3453),
.B(n_3187),
.Y(n_3619)
);

INVx1_ASAP7_75t_SL g3620 ( 
.A(n_3388),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3415),
.B(n_3373),
.Y(n_3621)
);

NAND3xp33_ASAP7_75t_SL g3622 ( 
.A(n_3386),
.B(n_3248),
.C(n_2855),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_3349),
.B(n_3423),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3481),
.B(n_3352),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3475),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3503),
.B(n_3216),
.Y(n_3626)
);

OR2x2_ASAP7_75t_L g3627 ( 
.A(n_3498),
.B(n_3054),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3512),
.B(n_3169),
.Y(n_3628)
);

INVxp67_ASAP7_75t_L g3629 ( 
.A(n_3391),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3460),
.B(n_3220),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3412),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3517),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3506),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3381),
.Y(n_3634)
);

AOI22xp5_ASAP7_75t_L g3635 ( 
.A1(n_3508),
.A2(n_3180),
.B1(n_3191),
.B2(n_3188),
.Y(n_3635)
);

INVxp67_ASAP7_75t_SL g3636 ( 
.A(n_3368),
.Y(n_3636)
);

AND2x6_ASAP7_75t_L g3637 ( 
.A(n_3334),
.B(n_3305),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_3484),
.B(n_3065),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3425),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3458),
.B(n_3198),
.Y(n_3640)
);

AOI221xp5_ASAP7_75t_L g3641 ( 
.A1(n_3582),
.A2(n_3479),
.B1(n_3382),
.B2(n_3511),
.C(n_3466),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3534),
.B(n_3404),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3595),
.A2(n_3375),
.B(n_3452),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3532),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_R g3645 ( 
.A(n_3571),
.B(n_3324),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3607),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_L g3647 ( 
.A(n_3614),
.B(n_3455),
.Y(n_3647)
);

BUFx2_ASAP7_75t_L g3648 ( 
.A(n_3555),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3617),
.B(n_3289),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3607),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3629),
.B(n_3427),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3532),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3536),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3541),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3548),
.Y(n_3655)
);

INVx4_ASAP7_75t_L g3656 ( 
.A(n_3587),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3536),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3621),
.B(n_3553),
.Y(n_3658)
);

BUFx2_ASAP7_75t_L g3659 ( 
.A(n_3579),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3617),
.B(n_3292),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3563),
.B(n_3404),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3552),
.Y(n_3662)
);

AOI31xp33_ASAP7_75t_L g3663 ( 
.A1(n_3620),
.A2(n_3421),
.A3(n_3422),
.B(n_3420),
.Y(n_3663)
);

INVxp67_ASAP7_75t_SL g3664 ( 
.A(n_3636),
.Y(n_3664)
);

OR2x2_ASAP7_75t_L g3665 ( 
.A(n_3542),
.B(n_3056),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_3612),
.B(n_3474),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3616),
.B(n_3462),
.Y(n_3667)
);

NOR2x1_ASAP7_75t_L g3668 ( 
.A(n_3624),
.B(n_3337),
.Y(n_3668)
);

AO21x2_ASAP7_75t_L g3669 ( 
.A1(n_3635),
.A2(n_3465),
.B(n_3457),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3609),
.B(n_3056),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3551),
.Y(n_3671)
);

OAI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3567),
.A2(n_3394),
.B(n_3447),
.Y(n_3672)
);

INVx4_ASAP7_75t_L g3673 ( 
.A(n_3634),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3562),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3564),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3573),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3631),
.B(n_3477),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3549),
.B(n_3472),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3561),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3566),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3576),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3633),
.B(n_3271),
.Y(n_3682)
);

AND2x2_ASAP7_75t_L g3683 ( 
.A(n_3559),
.B(n_3431),
.Y(n_3683)
);

INVx1_ASAP7_75t_SL g3684 ( 
.A(n_3623),
.Y(n_3684)
);

INVx2_ASAP7_75t_SL g3685 ( 
.A(n_3618),
.Y(n_3685)
);

HB1xp67_ASAP7_75t_L g3686 ( 
.A(n_3543),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3572),
.B(n_3445),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3584),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3583),
.B(n_3574),
.Y(n_3689)
);

INVx2_ASAP7_75t_SL g3690 ( 
.A(n_3545),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3601),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3540),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3630),
.B(n_3370),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3544),
.B(n_3486),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3547),
.Y(n_3695)
);

OR2x2_ASAP7_75t_L g3696 ( 
.A(n_3605),
.B(n_3305),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3633),
.B(n_3274),
.Y(n_3697)
);

AND2x4_ASAP7_75t_L g3698 ( 
.A(n_3538),
.B(n_3071),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3540),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3568),
.Y(n_3700)
);

INVx5_ASAP7_75t_SL g3701 ( 
.A(n_3581),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3546),
.B(n_3348),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3610),
.B(n_3275),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3570),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3585),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3586),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3598),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3632),
.Y(n_3708)
);

OAI21xp33_ASAP7_75t_L g3709 ( 
.A1(n_3580),
.A2(n_3358),
.B(n_3363),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3610),
.B(n_3279),
.Y(n_3710)
);

OAI21xp33_ASAP7_75t_L g3711 ( 
.A1(n_3535),
.A2(n_3378),
.B(n_3328),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3560),
.B(n_3454),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3604),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3533),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3588),
.B(n_3280),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3603),
.Y(n_3716)
);

AND2x4_ASAP7_75t_SL g3717 ( 
.A(n_3581),
.B(n_3323),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3619),
.B(n_3347),
.Y(n_3718)
);

AOI33xp33_ASAP7_75t_L g3719 ( 
.A1(n_3558),
.A2(n_2815),
.A3(n_2816),
.B1(n_2820),
.B2(n_2863),
.B3(n_2825),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3557),
.B(n_3490),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3625),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3569),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_SL g3723 ( 
.A(n_3554),
.B(n_3321),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3625),
.Y(n_3724)
);

BUFx6f_ASAP7_75t_SL g3725 ( 
.A(n_3655),
.Y(n_3725)
);

OR2x2_ASAP7_75t_L g3726 ( 
.A(n_3670),
.B(n_3611),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3656),
.B(n_3578),
.Y(n_3727)
);

AND2x4_ASAP7_75t_SL g3728 ( 
.A(n_3656),
.B(n_3320),
.Y(n_3728)
);

AOI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_3641),
.A2(n_3428),
.B1(n_3426),
.B2(n_3485),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3659),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3683),
.B(n_3639),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_SL g3732 ( 
.A(n_3673),
.B(n_3381),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3648),
.B(n_3639),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3658),
.B(n_3597),
.Y(n_3734)
);

OR2x2_ASAP7_75t_L g3735 ( 
.A(n_3696),
.B(n_3577),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3713),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3722),
.B(n_3575),
.Y(n_3737)
);

O2A1O1Ixp33_ASAP7_75t_L g3738 ( 
.A1(n_3672),
.A2(n_3608),
.B(n_3622),
.C(n_3565),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3642),
.B(n_3591),
.Y(n_3739)
);

INVx4_ASAP7_75t_L g3740 ( 
.A(n_3655),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3712),
.B(n_3606),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3721),
.B(n_3599),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3686),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3721),
.B(n_3626),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3689),
.B(n_3606),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3678),
.B(n_3538),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3702),
.B(n_3539),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3646),
.Y(n_3748)
);

OR2x2_ASAP7_75t_L g3749 ( 
.A(n_3714),
.B(n_3627),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3724),
.B(n_3613),
.Y(n_3750)
);

OR2x2_ASAP7_75t_L g3751 ( 
.A(n_3665),
.B(n_3593),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3661),
.B(n_3539),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3690),
.B(n_3638),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3724),
.B(n_3594),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3686),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3650),
.Y(n_3756)
);

OR2x2_ASAP7_75t_L g3757 ( 
.A(n_3716),
.B(n_3596),
.Y(n_3757)
);

AND2x4_ASAP7_75t_SL g3758 ( 
.A(n_3673),
.B(n_3437),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3644),
.B(n_3602),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3654),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3662),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3679),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3680),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3720),
.B(n_3638),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3667),
.B(n_3589),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3664),
.B(n_3640),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3644),
.B(n_3556),
.Y(n_3767)
);

NOR2x1_ASAP7_75t_L g3768 ( 
.A(n_3668),
.B(n_3432),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3700),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3704),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3705),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3706),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3652),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3652),
.B(n_3284),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3653),
.Y(n_3775)
);

XNOR2xp5_ASAP7_75t_L g3776 ( 
.A(n_3641),
.B(n_3317),
.Y(n_3776)
);

BUFx2_ASAP7_75t_L g3777 ( 
.A(n_3645),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3666),
.B(n_3589),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3677),
.B(n_3718),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3651),
.B(n_3592),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3653),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3651),
.B(n_3592),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3694),
.B(n_3615),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3707),
.Y(n_3784)
);

AOI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3672),
.A2(n_3537),
.B1(n_3526),
.B2(n_3590),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3657),
.B(n_3550),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3664),
.B(n_3628),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3685),
.B(n_3637),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3657),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3695),
.B(n_3307),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3692),
.B(n_3301),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3692),
.B(n_3301),
.Y(n_3792)
);

OR2x2_ASAP7_75t_L g3793 ( 
.A(n_3708),
.B(n_3307),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3687),
.B(n_3637),
.Y(n_3794)
);

OR2x2_ASAP7_75t_L g3795 ( 
.A(n_3708),
.B(n_3671),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3693),
.B(n_3637),
.Y(n_3796)
);

NAND2xp33_ASAP7_75t_SL g3797 ( 
.A(n_3740),
.B(n_3645),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3766),
.B(n_3669),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3754),
.B(n_3669),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3754),
.B(n_3643),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3759),
.B(n_3643),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_L g3802 ( 
.A(n_3777),
.B(n_3723),
.Y(n_3802)
);

NOR2xp67_ASAP7_75t_L g3803 ( 
.A(n_3740),
.B(n_3709),
.Y(n_3803)
);

AO221x2_ASAP7_75t_L g3804 ( 
.A1(n_3728),
.A2(n_3405),
.B1(n_3663),
.B2(n_3321),
.C(n_3316),
.Y(n_3804)
);

OAI22xp33_ASAP7_75t_L g3805 ( 
.A1(n_3732),
.A2(n_3441),
.B1(n_3461),
.B2(n_3487),
.Y(n_3805)
);

NAND2xp33_ASAP7_75t_R g3806 ( 
.A(n_3732),
.B(n_3406),
.Y(n_3806)
);

NOR2xp67_ASAP7_75t_L g3807 ( 
.A(n_3729),
.B(n_3711),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_SL g3808 ( 
.A(n_3725),
.B(n_3369),
.Y(n_3808)
);

OAI221xp5_ASAP7_75t_L g3809 ( 
.A1(n_3785),
.A2(n_3647),
.B1(n_3376),
.B2(n_3684),
.C(n_3516),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3759),
.B(n_3715),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3750),
.B(n_3715),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3795),
.Y(n_3812)
);

AO221x2_ASAP7_75t_L g3813 ( 
.A1(n_3725),
.A2(n_3379),
.B1(n_3351),
.B2(n_3491),
.C(n_3528),
.Y(n_3813)
);

AOI22xp5_ASAP7_75t_SL g3814 ( 
.A1(n_3727),
.A2(n_3647),
.B1(n_3336),
.B2(n_3359),
.Y(n_3814)
);

NOR2x1_ASAP7_75t_L g3815 ( 
.A(n_3768),
.B(n_3408),
.Y(n_3815)
);

OAI22xp33_ASAP7_75t_L g3816 ( 
.A1(n_3729),
.A2(n_3482),
.B1(n_3366),
.B2(n_3329),
.Y(n_3816)
);

OR2x2_ASAP7_75t_L g3817 ( 
.A(n_3751),
.B(n_3674),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3750),
.B(n_3649),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3736),
.B(n_3649),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3743),
.B(n_3660),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3755),
.B(n_3660),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3767),
.B(n_3682),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3758),
.B(n_3717),
.Y(n_3823)
);

OAI22xp33_ASAP7_75t_L g3824 ( 
.A1(n_3787),
.A2(n_3408),
.B1(n_3346),
.B2(n_3515),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3767),
.B(n_3682),
.Y(n_3825)
);

AOI22xp33_ASAP7_75t_L g3826 ( 
.A1(n_3733),
.A2(n_3776),
.B1(n_3788),
.B2(n_3730),
.Y(n_3826)
);

INVxp33_ASAP7_75t_SL g3827 ( 
.A(n_3796),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_R g3828 ( 
.A(n_3794),
.B(n_3444),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3735),
.B(n_3697),
.Y(n_3829)
);

OAI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_3786),
.A2(n_3515),
.B1(n_3488),
.B2(n_3451),
.Y(n_3830)
);

OAI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3786),
.A2(n_3488),
.B1(n_3459),
.B2(n_3456),
.Y(n_3831)
);

NAND2xp33_ASAP7_75t_R g3832 ( 
.A(n_3733),
.B(n_3407),
.Y(n_3832)
);

NOR2xp33_ASAP7_75t_L g3833 ( 
.A(n_3738),
.B(n_3331),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_L g3834 ( 
.A(n_3780),
.B(n_3717),
.Y(n_3834)
);

NAND2xp33_ASAP7_75t_SL g3835 ( 
.A(n_3753),
.B(n_3409),
.Y(n_3835)
);

NAND2xp33_ASAP7_75t_SL g3836 ( 
.A(n_3782),
.B(n_3410),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3760),
.B(n_3697),
.Y(n_3837)
);

AO221x2_ASAP7_75t_L g3838 ( 
.A1(n_3744),
.A2(n_3416),
.B1(n_3392),
.B2(n_3325),
.C(n_3429),
.Y(n_3838)
);

NAND2xp33_ASAP7_75t_SL g3839 ( 
.A(n_3779),
.B(n_3501),
.Y(n_3839)
);

AO221x2_ASAP7_75t_L g3840 ( 
.A1(n_3744),
.A2(n_3510),
.B1(n_3507),
.B2(n_3450),
.C(n_3442),
.Y(n_3840)
);

BUFx2_ASAP7_75t_L g3841 ( 
.A(n_3765),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_SL g3842 ( 
.A(n_3783),
.B(n_3519),
.Y(n_3842)
);

NAND2xp33_ASAP7_75t_SL g3843 ( 
.A(n_3745),
.B(n_3326),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3819),
.Y(n_3844)
);

INVx2_ASAP7_75t_SL g3845 ( 
.A(n_3804),
.Y(n_3845)
);

AOI222xp33_ASAP7_75t_L g3846 ( 
.A1(n_3807),
.A2(n_3312),
.B1(n_3367),
.B2(n_3600),
.C1(n_3430),
.C2(n_3761),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3818),
.B(n_3762),
.Y(n_3847)
);

INVx1_ASAP7_75t_SL g3848 ( 
.A(n_3797),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3817),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3810),
.B(n_3763),
.Y(n_3850)
);

OR2x2_ASAP7_75t_L g3851 ( 
.A(n_3811),
.B(n_3742),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3800),
.B(n_3769),
.Y(n_3852)
);

INVx1_ASAP7_75t_SL g3853 ( 
.A(n_3839),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3837),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3829),
.Y(n_3855)
);

OR2x2_ASAP7_75t_L g3856 ( 
.A(n_3822),
.B(n_3742),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3825),
.B(n_3801),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3804),
.A2(n_3637),
.B1(n_3327),
.B2(n_3353),
.Y(n_3858)
);

HB1xp67_ASAP7_75t_L g3859 ( 
.A(n_3803),
.Y(n_3859)
);

INVx2_ASAP7_75t_SL g3860 ( 
.A(n_3823),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3802),
.B(n_3752),
.Y(n_3861)
);

AOI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3813),
.A2(n_3737),
.B1(n_3439),
.B2(n_3739),
.Y(n_3862)
);

OAI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3832),
.A2(n_3726),
.B1(n_3749),
.B2(n_3757),
.Y(n_3863)
);

AND2x4_ASAP7_75t_L g3864 ( 
.A(n_3815),
.B(n_3741),
.Y(n_3864)
);

HB1xp67_ASAP7_75t_L g3865 ( 
.A(n_3820),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3812),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3826),
.B(n_3778),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3841),
.B(n_3834),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3821),
.Y(n_3869)
);

HB1xp67_ASAP7_75t_L g3870 ( 
.A(n_3799),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3798),
.B(n_3793),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3827),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3828),
.B(n_3764),
.Y(n_3873)
);

AOI222xp33_ASAP7_75t_L g3874 ( 
.A1(n_3833),
.A2(n_3770),
.B1(n_3771),
.B2(n_3784),
.C1(n_3772),
.C2(n_3440),
.Y(n_3874)
);

INVx2_ASAP7_75t_SL g3875 ( 
.A(n_3838),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3831),
.B(n_3748),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3842),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3814),
.B(n_3747),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3830),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3806),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3816),
.B(n_3790),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3813),
.B(n_3756),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3838),
.B(n_3746),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3840),
.B(n_3731),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3843),
.B(n_3773),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3835),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3840),
.B(n_3734),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3836),
.Y(n_3888)
);

INVxp67_ASAP7_75t_L g3889 ( 
.A(n_3809),
.Y(n_3889)
);

OR2x2_ASAP7_75t_L g3890 ( 
.A(n_3824),
.B(n_3775),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3808),
.Y(n_3891)
);

NAND3xp33_ASAP7_75t_SL g3892 ( 
.A(n_3805),
.B(n_3436),
.C(n_3514),
.Y(n_3892)
);

OAI21x1_ASAP7_75t_L g3893 ( 
.A1(n_3815),
.A2(n_3792),
.B(n_3791),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3802),
.B(n_3698),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3817),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3849),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3845),
.A2(n_3502),
.B1(n_3456),
.B2(n_3698),
.Y(n_3897)
);

OR2x2_ASAP7_75t_L g3898 ( 
.A(n_3857),
.B(n_3774),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3872),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3895),
.Y(n_3900)
);

OAI221xp5_ASAP7_75t_L g3901 ( 
.A1(n_3846),
.A2(n_3383),
.B1(n_3710),
.B2(n_3703),
.C(n_3792),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3880),
.A2(n_3791),
.B(n_3383),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3846),
.B(n_3855),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3891),
.B(n_3789),
.Y(n_3904)
);

AND2x4_ASAP7_75t_L g3905 ( 
.A(n_3860),
.B(n_3781),
.Y(n_3905)
);

AOI22xp33_ASAP7_75t_L g3906 ( 
.A1(n_3879),
.A2(n_3489),
.B1(n_3463),
.B2(n_3703),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3865),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3844),
.B(n_3854),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3852),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3850),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3875),
.A2(n_3399),
.B1(n_3395),
.B2(n_3524),
.Y(n_3911)
);

INVx1_ASAP7_75t_SL g3912 ( 
.A(n_3848),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3866),
.Y(n_3913)
);

OR2x2_ASAP7_75t_L g3914 ( 
.A(n_3856),
.B(n_3774),
.Y(n_3914)
);

AOI22xp5_ASAP7_75t_L g3915 ( 
.A1(n_3853),
.A2(n_3494),
.B1(n_3483),
.B2(n_3204),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3883),
.B(n_3699),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3850),
.Y(n_3917)
);

AOI221xp5_ASAP7_75t_L g3918 ( 
.A1(n_3889),
.A2(n_3710),
.B1(n_2788),
.B2(n_3699),
.C(n_2764),
.Y(n_3918)
);

OAI22xp5_ASAP7_75t_L g3919 ( 
.A1(n_3862),
.A2(n_3527),
.B1(n_3701),
.B2(n_3676),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3868),
.B(n_3853),
.Y(n_3920)
);

AOI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3848),
.A2(n_3154),
.B(n_2798),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3874),
.B(n_3675),
.Y(n_3922)
);

AOI221xp5_ASAP7_75t_L g3923 ( 
.A1(n_3882),
.A2(n_2729),
.B1(n_3688),
.B2(n_3691),
.C(n_3681),
.Y(n_3923)
);

BUFx2_ASAP7_75t_L g3924 ( 
.A(n_3859),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3847),
.Y(n_3925)
);

AOI221xp5_ASAP7_75t_L g3926 ( 
.A1(n_3882),
.A2(n_2949),
.B1(n_3203),
.B2(n_3208),
.C(n_3205),
.Y(n_3926)
);

INVxp67_ASAP7_75t_SL g3927 ( 
.A(n_3876),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3847),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_3877),
.B(n_3581),
.Y(n_3929)
);

HB1xp67_ASAP7_75t_L g3930 ( 
.A(n_3870),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3910),
.B(n_3869),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3899),
.Y(n_3932)
);

INVxp67_ASAP7_75t_L g3933 ( 
.A(n_3924),
.Y(n_3933)
);

HB1xp67_ASAP7_75t_L g3934 ( 
.A(n_3930),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3907),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3927),
.B(n_3874),
.Y(n_3936)
);

INVx2_ASAP7_75t_SL g3937 ( 
.A(n_3905),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3920),
.B(n_3884),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3896),
.Y(n_3939)
);

INVx2_ASAP7_75t_SL g3940 ( 
.A(n_3905),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3912),
.B(n_3867),
.Y(n_3941)
);

INVx2_ASAP7_75t_SL g3942 ( 
.A(n_3900),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3903),
.B(n_3878),
.Y(n_3943)
);

INVx1_ASAP7_75t_SL g3944 ( 
.A(n_3908),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3915),
.B(n_3887),
.Y(n_3945)
);

NAND2x1p5_ASAP7_75t_L g3946 ( 
.A(n_3913),
.B(n_3864),
.Y(n_3946)
);

OR2x2_ASAP7_75t_L g3947 ( 
.A(n_3898),
.B(n_3914),
.Y(n_3947)
);

AND2x2_ASAP7_75t_L g3948 ( 
.A(n_3906),
.B(n_3864),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3904),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3916),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3909),
.Y(n_3951)
);

HB1xp67_ASAP7_75t_L g3952 ( 
.A(n_3917),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3929),
.B(n_3888),
.Y(n_3953)
);

OAI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3901),
.A2(n_3886),
.B(n_3876),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3925),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3928),
.B(n_3851),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3915),
.B(n_3926),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3934),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3933),
.Y(n_3959)
);

BUFx6f_ASAP7_75t_L g3960 ( 
.A(n_3937),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3942),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3939),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3940),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3947),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3949),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3948),
.B(n_3861),
.Y(n_3966)
);

INVx1_ASAP7_75t_SL g3967 ( 
.A(n_3953),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3952),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3935),
.Y(n_3969)
);

INVxp67_ASAP7_75t_L g3970 ( 
.A(n_3941),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3931),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3931),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3944),
.B(n_3911),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3956),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3956),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3932),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3951),
.Y(n_3977)
);

OR2x2_ASAP7_75t_L g3978 ( 
.A(n_3944),
.B(n_3881),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3955),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3938),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3946),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3946),
.Y(n_3982)
);

NOR3xp33_ASAP7_75t_L g3983 ( 
.A(n_3959),
.B(n_3936),
.C(n_3943),
.Y(n_3983)
);

NAND3xp33_ASAP7_75t_L g3984 ( 
.A(n_3960),
.B(n_3954),
.C(n_3923),
.Y(n_3984)
);

NAND3xp33_ASAP7_75t_SL g3985 ( 
.A(n_3967),
.B(n_3954),
.C(n_3957),
.Y(n_3985)
);

AOI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3973),
.A2(n_3945),
.B(n_3957),
.Y(n_3986)
);

NAND4xp25_ASAP7_75t_L g3987 ( 
.A(n_3963),
.B(n_3858),
.C(n_3918),
.D(n_3892),
.Y(n_3987)
);

NAND3x1_ASAP7_75t_L g3988 ( 
.A(n_3981),
.B(n_3922),
.C(n_3902),
.Y(n_3988)
);

NOR2xp33_ASAP7_75t_SL g3989 ( 
.A(n_3961),
.B(n_3863),
.Y(n_3989)
);

NOR3xp33_ASAP7_75t_L g3990 ( 
.A(n_3958),
.B(n_3897),
.C(n_3919),
.Y(n_3990)
);

NAND4xp25_ASAP7_75t_L g3991 ( 
.A(n_3970),
.B(n_3982),
.C(n_3964),
.D(n_3978),
.Y(n_3991)
);

NAND4xp25_ASAP7_75t_SL g3992 ( 
.A(n_3980),
.B(n_3911),
.C(n_3921),
.D(n_3873),
.Y(n_3992)
);

OAI32xp33_ASAP7_75t_L g3993 ( 
.A1(n_3974),
.A2(n_3950),
.A3(n_3885),
.B1(n_3890),
.B2(n_3871),
.Y(n_3993)
);

NAND4xp25_ASAP7_75t_L g3994 ( 
.A(n_3975),
.B(n_3719),
.C(n_3894),
.D(n_2897),
.Y(n_3994)
);

NOR2x1_ASAP7_75t_L g3995 ( 
.A(n_3958),
.B(n_3960),
.Y(n_3995)
);

NAND4xp25_ASAP7_75t_L g3996 ( 
.A(n_3968),
.B(n_3719),
.C(n_2969),
.D(n_2955),
.Y(n_3996)
);

NOR3xp33_ASAP7_75t_L g3997 ( 
.A(n_3962),
.B(n_3893),
.C(n_2967),
.Y(n_3997)
);

NOR3x1_ASAP7_75t_L g3998 ( 
.A(n_3971),
.B(n_3004),
.C(n_2970),
.Y(n_3998)
);

NAND3xp33_ASAP7_75t_L g3999 ( 
.A(n_3960),
.B(n_2989),
.C(n_2985),
.Y(n_3999)
);

NAND3xp33_ASAP7_75t_SL g4000 ( 
.A(n_3983),
.B(n_3972),
.C(n_3965),
.Y(n_4000)
);

AOI211xp5_ASAP7_75t_L g4001 ( 
.A1(n_3985),
.A2(n_3969),
.B(n_3977),
.C(n_3979),
.Y(n_4001)
);

AOI221x1_ASAP7_75t_L g4002 ( 
.A1(n_3991),
.A2(n_3976),
.B1(n_3966),
.B2(n_2875),
.C(n_2932),
.Y(n_4002)
);

INVx1_ASAP7_75t_SL g4003 ( 
.A(n_3995),
.Y(n_4003)
);

AOI221xp5_ASAP7_75t_L g4004 ( 
.A1(n_3986),
.A2(n_2995),
.B1(n_2922),
.B2(n_2843),
.C(n_3002),
.Y(n_4004)
);

OAI222xp33_ASAP7_75t_L g4005 ( 
.A1(n_3992),
.A2(n_3988),
.B1(n_3987),
.B2(n_3990),
.C1(n_3984),
.C2(n_3989),
.Y(n_4005)
);

AOI211xp5_ASAP7_75t_L g4006 ( 
.A1(n_3993),
.A2(n_3004),
.B(n_2970),
.C(n_2976),
.Y(n_4006)
);

AOI221xp5_ASAP7_75t_L g4007 ( 
.A1(n_3997),
.A2(n_3994),
.B1(n_3996),
.B2(n_3999),
.C(n_3998),
.Y(n_4007)
);

AOI221xp5_ASAP7_75t_SL g4008 ( 
.A1(n_3986),
.A2(n_2910),
.B1(n_2932),
.B2(n_2875),
.C(n_3042),
.Y(n_4008)
);

XNOR2xp5_ASAP7_75t_L g4009 ( 
.A(n_3985),
.B(n_793),
.Y(n_4009)
);

OAI221xp5_ASAP7_75t_L g4010 ( 
.A1(n_3987),
.A2(n_2993),
.B1(n_3037),
.B2(n_3034),
.C(n_3029),
.Y(n_4010)
);

AOI211x1_ASAP7_75t_SL g4011 ( 
.A1(n_3985),
.A2(n_2888),
.B(n_2901),
.C(n_2910),
.Y(n_4011)
);

AOI211xp5_ASAP7_75t_L g4012 ( 
.A1(n_3985),
.A2(n_2965),
.B(n_2971),
.C(n_3253),
.Y(n_4012)
);

INVxp67_ASAP7_75t_SL g4013 ( 
.A(n_3995),
.Y(n_4013)
);

NOR3xp33_ASAP7_75t_L g4014 ( 
.A(n_3985),
.B(n_2965),
.C(n_3011),
.Y(n_4014)
);

INVx2_ASAP7_75t_SL g4015 ( 
.A(n_4003),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_4013),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_4009),
.B(n_794),
.Y(n_4017)
);

OR2x2_ASAP7_75t_L g4018 ( 
.A(n_4000),
.B(n_794),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_4011),
.B(n_795),
.Y(n_4019)
);

HB1xp67_ASAP7_75t_L g4020 ( 
.A(n_4014),
.Y(n_4020)
);

OAI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_4007),
.A2(n_3701),
.B1(n_3448),
.B2(n_2994),
.Y(n_4021)
);

NAND2xp33_ASAP7_75t_SL g4022 ( 
.A(n_4018),
.B(n_4015),
.Y(n_4022)
);

NOR2xp33_ASAP7_75t_R g4023 ( 
.A(n_4016),
.B(n_797),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_4020),
.B(n_4001),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_4017),
.B(n_4012),
.Y(n_4025)
);

XNOR2xp5_ASAP7_75t_L g4026 ( 
.A(n_4021),
.B(n_4002),
.Y(n_4026)
);

NOR3xp33_ASAP7_75t_SL g4027 ( 
.A(n_4022),
.B(n_4005),
.C(n_4019),
.Y(n_4027)
);

AO22x2_ASAP7_75t_L g4028 ( 
.A1(n_4025),
.A2(n_4008),
.B1(n_4006),
.B2(n_4010),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_4028),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_4027),
.B(n_4026),
.Y(n_4030)
);

OAI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_4030),
.A2(n_4024),
.B1(n_4023),
.B2(n_4004),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_4029),
.B(n_797),
.Y(n_4032)
);

AOI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_4032),
.A2(n_3701),
.B1(n_3433),
.B2(n_3224),
.Y(n_4033)
);

AOI31xp33_ASAP7_75t_L g4034 ( 
.A1(n_4031),
.A2(n_801),
.A3(n_798),
.B(n_799),
.Y(n_4034)
);

XNOR2x1_ASAP7_75t_L g4035 ( 
.A(n_4034),
.B(n_798),
.Y(n_4035)
);

AOI222xp33_ASAP7_75t_L g4036 ( 
.A1(n_4035),
.A2(n_4033),
.B1(n_2923),
.B2(n_2960),
.C1(n_2903),
.C2(n_3433),
.Y(n_4036)
);

INVx4_ASAP7_75t_L g4037 ( 
.A(n_4036),
.Y(n_4037)
);

OAI221xp5_ASAP7_75t_R g4038 ( 
.A1(n_4037),
.A2(n_3022),
.B1(n_2979),
.B2(n_802),
.C(n_803),
.Y(n_4038)
);

AOI22xp33_ASAP7_75t_SL g4039 ( 
.A1(n_4038),
.A2(n_2953),
.B1(n_3529),
.B2(n_3024),
.Y(n_4039)
);


endmodule