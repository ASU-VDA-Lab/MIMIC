module fake_ibex_1037_n_1282 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1282);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1282;

wire n_1084;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1129;
wire n_1244;
wire n_449;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_485;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_996;
wire n_915;
wire n_1174;
wire n_542;
wire n_900;
wire n_377;
wire n_647;
wire n_317;
wire n_326;
wire n_270;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_277;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_632;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_987;
wire n_750;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1277;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_117),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_24),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_189),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_172),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_119),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_143),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_126),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_156),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_97),
.Y(n_282)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_37),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_54),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_168),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_99),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_109),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_152),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_70),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_13),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_42),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_155),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_198),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_163),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_132),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_205),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_134),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_140),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_59),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_47),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_157),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_47),
.B(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_118),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_7),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_179),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_34),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_3),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_90),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_107),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_31),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_241),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_167),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_26),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_146),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_123),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_147),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_65),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_225),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_16),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_220),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_66),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_89),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_149),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_125),
.B(n_184),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_190),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_49),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_38),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_234),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_249),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_33),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_108),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_29),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_5),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_211),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_166),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_199),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_24),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_136),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_77),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_35),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_11),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_237),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_122),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_238),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_160),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_28),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_76),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_265),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_203),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_151),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_232),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_221),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_173),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_120),
.Y(n_365)
);

BUFx8_ASAP7_75t_SL g366 ( 
.A(n_68),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_169),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_63),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_96),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_171),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_261),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_38),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_148),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_202),
.B(n_161),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_128),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_230),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_129),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_112),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_121),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_62),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_30),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_219),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_214),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_222),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_91),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_212),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_150),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_217),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_138),
.Y(n_390)
);

BUFx8_ASAP7_75t_SL g391 ( 
.A(n_264),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_183),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_130),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_46),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_95),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_187),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_182),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_208),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_247),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_174),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_197),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_73),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_13),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_42),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_0),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_51),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_181),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_116),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_27),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_200),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_88),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_178),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_41),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_131),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_256),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_188),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_40),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_75),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_245),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_61),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_175),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_159),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_139),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_259),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_58),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_81),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_45),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_31),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_85),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_106),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_3),
.B(n_33),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_162),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_207),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_83),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_18),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_176),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_193),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_254),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_153),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_250),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_251),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_12),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_32),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_206),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_1),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_227),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_74),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_248),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_195),
.Y(n_449)
);

OA22x2_ASAP7_75t_SL g450 ( 
.A1(n_366),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_296),
.Y(n_451)
);

AOI22x1_ASAP7_75t_SL g452 ( 
.A1(n_292),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_328),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_266),
.A2(n_87),
.B(n_86),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_444),
.A2(n_93),
.B(n_92),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_266),
.A2(n_98),
.B(n_94),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

OAI22x1_ASAP7_75t_R g461 ( 
.A1(n_292),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_296),
.Y(n_463)
);

OAI22x1_ASAP7_75t_R g464 ( 
.A1(n_297),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_306),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_394),
.B(n_9),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_352),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_300),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_352),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_300),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_269),
.B(n_10),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_297),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_300),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_306),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_352),
.Y(n_475)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_387),
.A2(n_101),
.B(n_100),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_352),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_387),
.A2(n_103),
.B(n_102),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_281),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_268),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_290),
.B(n_17),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_306),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_359),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_388),
.A2(n_105),
.B(n_104),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_281),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_368),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_350),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_418),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_274),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_393),
.B(n_20),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_300),
.Y(n_494)
);

AOI22x1_ASAP7_75t_SL g495 ( 
.A1(n_368),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_391),
.B(n_401),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_276),
.B(n_22),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_317),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_278),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_279),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_280),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_319),
.B(n_23),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_317),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_317),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_391),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_350),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_366),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_307),
.B(n_25),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_283),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_317),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_270),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_420),
.B(n_29),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_294),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_301),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_318),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_390),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_426),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_418),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_271),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_426),
.Y(n_527)
);

BUFx12f_ASAP7_75t_L g528 ( 
.A(n_284),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_390),
.B(n_30),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_430),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_400),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_388),
.A2(n_135),
.B(n_262),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_302),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_483),
.B(n_420),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_483),
.B(n_427),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_510),
.B(n_396),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_465),
.B(n_430),
.Y(n_537)
);

BUFx6f_ASAP7_75t_SL g538 ( 
.A(n_482),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_510),
.B(n_396),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_466),
.A2(n_285),
.B1(n_298),
.B2(n_295),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_466),
.A2(n_308),
.B1(n_315),
.B2(n_313),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_528),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g546 ( 
.A(n_482),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_487),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_467),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_453),
.B(n_427),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_466),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_510),
.B(n_423),
.Y(n_551)
);

CKINVDCx6p67_ASAP7_75t_R g552 ( 
.A(n_528),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_490),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_508),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_483),
.B(n_423),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_503),
.Y(n_559)
);

NOR3xp33_ASAP7_75t_L g560 ( 
.A(n_472),
.B(n_344),
.C(n_309),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_453),
.B(n_284),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_506),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_455),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_529),
.B(n_436),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_451),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_481),
.B(n_436),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_456),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_501),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_489),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_456),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_511),
.A2(n_496),
.B1(n_445),
.B2(n_434),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_460),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_462),
.B(n_287),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_469),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_507),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_507),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_489),
.B(n_419),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_477),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_465),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_530),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_475),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_485),
.B(n_304),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_492),
.B(n_430),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_517),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_492),
.B(n_419),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_499),
.A2(n_343),
.B1(n_348),
.B2(n_330),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_451),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_500),
.B(n_321),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_500),
.B(n_324),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_471),
.B(n_493),
.C(n_514),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_488),
.B(n_431),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_502),
.B(n_312),
.Y(n_600)
);

BUFx6f_ASAP7_75t_SL g601 ( 
.A(n_502),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_513),
.B(n_332),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_515),
.B(n_337),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_515),
.B(n_341),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_525),
.Y(n_605)
);

CKINVDCx11_ASAP7_75t_R g606 ( 
.A(n_522),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_516),
.B(n_533),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_533),
.B(n_381),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_497),
.B(n_406),
.C(n_404),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_477),
.A2(n_357),
.B1(n_358),
.B2(n_351),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_509),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_509),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_519),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_519),
.B(n_325),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_477),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_522),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_463),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_468),
.B(n_329),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_484),
.B(n_413),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_468),
.B(n_333),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_463),
.Y(n_622)
);

BUFx16f_ASAP7_75t_R g623 ( 
.A(n_461),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_468),
.B(n_340),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_463),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_491),
.B(n_447),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_463),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_470),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_468),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_470),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_491),
.B(n_347),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_468),
.B(n_353),
.Y(n_632)
);

CKINVDCx6p67_ASAP7_75t_R g633 ( 
.A(n_527),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_464),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_473),
.B(n_355),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_473),
.B(n_360),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_473),
.B(n_361),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_523),
.Y(n_638)
);

OAI22xp33_ASAP7_75t_L g639 ( 
.A1(n_480),
.A2(n_445),
.B1(n_434),
.B2(n_283),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

CKINVDCx6p67_ASAP7_75t_R g641 ( 
.A(n_527),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_523),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_512),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_479),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_494),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_454),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_494),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_494),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_494),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_486),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_450),
.B(n_372),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_512),
.B(n_267),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_494),
.B(n_282),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_457),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_512),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_454),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_454),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_512),
.B(n_362),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_498),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_458),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_592),
.B(n_272),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_553),
.B(n_275),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_607),
.B(n_288),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_550),
.A2(n_382),
.B1(n_403),
.B2(n_402),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_553),
.B(n_289),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_534),
.B(n_364),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_543),
.A2(n_286),
.B1(n_299),
.B2(n_282),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_555),
.A2(n_409),
.B1(n_425),
.B2(n_417),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_582),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_547),
.B(n_338),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_557),
.A2(n_559),
.B1(n_563),
.B2(n_561),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_595),
.B(n_596),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_603),
.B(n_291),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_604),
.B(n_608),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_535),
.B(n_293),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_597),
.B(n_369),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_539),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_543),
.B(n_303),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_591),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_605),
.B(n_305),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_581),
.B(n_310),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_616),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_565),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_562),
.B(n_314),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_544),
.B(n_320),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_602),
.B(n_322),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_588),
.B(n_323),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_588),
.B(n_326),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_570),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_558),
.B(n_327),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_558),
.B(n_331),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_556),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_573),
.Y(n_695)
);

AO22x2_ASAP7_75t_L g696 ( 
.A1(n_634),
.A2(n_495),
.B1(n_452),
.B2(n_429),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_563),
.A2(n_428),
.B1(n_442),
.B2(n_435),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_544),
.B(n_334),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_539),
.B(n_335),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_549),
.B(n_339),
.Y(n_700)
);

BUFx8_ASAP7_75t_L g701 ( 
.A(n_601),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_583),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_609),
.B(n_371),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_536),
.B(n_345),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_542),
.B(n_346),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_599),
.A2(n_574),
.B1(n_639),
.B2(n_299),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_614),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_577),
.B(n_286),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_552),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_572),
.A2(n_336),
.B1(n_367),
.B2(n_365),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_538),
.A2(n_365),
.B1(n_367),
.B2(n_336),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_538),
.A2(n_411),
.B1(n_437),
.B2(n_392),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_542),
.B(n_349),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_617),
.B(n_443),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_631),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_583),
.B(n_354),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_546),
.B(n_378),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_631),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_551),
.B(n_356),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_566),
.B(n_363),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_545),
.B(n_392),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_600),
.B(n_370),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_601),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_600),
.B(n_373),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_546),
.B(n_613),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_569),
.B(n_375),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_615),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_626),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_587),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_644),
.A2(n_650),
.B1(n_652),
.B2(n_655),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_593),
.B(n_376),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_569),
.B(n_379),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_654),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_568),
.B(n_380),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_610),
.A2(n_342),
.B1(n_311),
.B2(n_415),
.C(n_383),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_537),
.B(n_395),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_575),
.B(n_408),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_611),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_571),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_576),
.B(n_410),
.Y(n_742)
);

XNOR2xp5_ASAP7_75t_L g743 ( 
.A(n_574),
.B(n_452),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_657),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_578),
.B(n_412),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_584),
.B(n_385),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_639),
.B(n_316),
.C(n_414),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_610),
.A2(n_437),
.B1(n_411),
.B2(n_448),
.C(n_441),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_586),
.B(n_386),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_564),
.B(n_458),
.Y(n_751)
);

OR2x2_ASAP7_75t_SL g752 ( 
.A(n_623),
.B(n_606),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_651),
.A2(n_432),
.B1(n_439),
.B2(n_449),
.Y(n_753)
);

BUFx4_ASAP7_75t_L g754 ( 
.A(n_606),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_612),
.Y(n_755)
);

AND2x6_ASAP7_75t_SL g756 ( 
.A(n_599),
.B(n_495),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_560),
.A2(n_422),
.B1(n_433),
.B2(n_416),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_589),
.B(n_389),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_587),
.B(n_397),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_590),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_633),
.B(n_32),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_579),
.B(n_398),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_661),
.A2(n_532),
.B(n_476),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_590),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_641),
.B(n_34),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_580),
.B(n_407),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_580),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_619),
.B(n_273),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_599),
.A2(n_277),
.B(n_384),
.C(n_374),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_585),
.B(n_35),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_585),
.A2(n_421),
.B1(n_424),
.B2(n_521),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_540),
.B(n_438),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_619),
.B(n_440),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_541),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_541),
.B(n_446),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_648),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_621),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_624),
.B(n_36),
.C(n_39),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_624),
.B(n_421),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_632),
.B(n_518),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_632),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_548),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_518),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_635),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_636),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_636),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_637),
.B(n_521),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_659),
.B(n_521),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_653),
.B(n_521),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_659),
.B(n_643),
.Y(n_791)
);

AND2x2_ASAP7_75t_SL g792 ( 
.A(n_638),
.B(n_640),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_656),
.B(n_526),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_629),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_642),
.A2(n_526),
.B1(n_524),
.B2(n_520),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_660),
.B(n_526),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_567),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_701),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_678),
.A2(n_504),
.B(n_505),
.C(n_520),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_702),
.B(n_41),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_672),
.B(n_776),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_L g802 ( 
.A1(n_672),
.A2(n_747),
.B(n_671),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_694),
.B(n_43),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_679),
.B(n_43),
.Y(n_804)
);

NOR4xp25_ASAP7_75t_SL g805 ( 
.A(n_748),
.B(n_44),
.C(n_45),
.D(n_46),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_782),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_694),
.B(n_48),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_747),
.A2(n_649),
.B(n_647),
.C(n_645),
.Y(n_808)
);

AO21x1_ASAP7_75t_L g809 ( 
.A1(n_751),
.A2(n_622),
.B(n_618),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_681),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_710),
.A2(n_504),
.B1(n_505),
.B2(n_520),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_724),
.B(n_50),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_729),
.B(n_678),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_715),
.A2(n_505),
.B(n_520),
.C(n_524),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_730),
.B(n_51),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_776),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_700),
.B(n_52),
.Y(n_817)
);

OAI321xp33_ASAP7_75t_L g818 ( 
.A1(n_706),
.A2(n_524),
.A3(n_628),
.B1(n_627),
.B2(n_625),
.C(n_630),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_718),
.A2(n_524),
.B(n_598),
.C(n_594),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_730),
.B(n_52),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_673),
.B(n_53),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_701),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_673),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_783),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_708),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_667),
.B(n_55),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_667),
.B(n_56),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_767),
.A2(n_764),
.B(n_760),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_685),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_744),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_686),
.B(n_57),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_669),
.B(n_57),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_669),
.B(n_58),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_699),
.B(n_688),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_664),
.B(n_59),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_759),
.A2(n_170),
.B(n_258),
.Y(n_836)
);

O2A1O1Ixp5_ASAP7_75t_L g837 ( 
.A1(n_703),
.A2(n_164),
.B(n_257),
.C(n_253),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_706),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_721),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_711),
.B(n_63),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_774),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_709),
.B(n_64),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_746),
.A2(n_749),
.B(n_662),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_744),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_740),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_744),
.A2(n_766),
.B(n_762),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_737),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_697),
.B(n_67),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_665),
.B(n_69),
.Y(n_849)
);

INVx3_ASAP7_75t_SL g850 ( 
.A(n_752),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_723),
.B(n_70),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_772),
.A2(n_677),
.B(n_675),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_714),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_774),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_854)
);

OAI321xp33_ASAP7_75t_L g855 ( 
.A1(n_770),
.A2(n_75),
.A3(n_76),
.B1(n_78),
.B2(n_79),
.C(n_80),
.Y(n_855)
);

CKINVDCx10_ASAP7_75t_R g856 ( 
.A(n_754),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_755),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_665),
.A2(n_712),
.B1(n_738),
.B2(n_734),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_682),
.A2(n_693),
.B(n_692),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_739),
.A2(n_180),
.B(n_246),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_740),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_761),
.B(n_78),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_696),
.B(n_82),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_765),
.Y(n_864)
);

AO21x1_ASAP7_75t_L g865 ( 
.A1(n_778),
.A2(n_84),
.B(n_110),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_728),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_689),
.B(n_111),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_690),
.B(n_244),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_680),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_683),
.B(n_124),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_792),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_691),
.A2(n_695),
.B1(n_735),
.B2(n_742),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_753),
.A2(n_698),
.B(n_687),
.C(n_732),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_704),
.A2(n_127),
.B(n_133),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_705),
.A2(n_137),
.B(n_142),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_713),
.A2(n_144),
.B(n_145),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_719),
.A2(n_154),
.B(n_158),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_684),
.Y(n_878)
);

OAI21xp33_ASAP7_75t_L g879 ( 
.A1(n_745),
.A2(n_717),
.B(n_757),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_745),
.B(n_242),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_720),
.A2(n_185),
.B1(n_186),
.B2(n_191),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_790),
.A2(n_192),
.B(n_194),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_722),
.A2(n_196),
.B1(n_204),
.B2(n_209),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_725),
.A2(n_216),
.B(n_218),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_794),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_716),
.B(n_223),
.Y(n_886)
);

BUFx4f_ASAP7_75t_L g887 ( 
.A(n_791),
.Y(n_887)
);

OR2x6_ASAP7_75t_SL g888 ( 
.A(n_743),
.B(n_224),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_663),
.B(n_226),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_769),
.B(n_228),
.C(n_231),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_741),
.A2(n_235),
.B(n_750),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_794),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_666),
.B(n_758),
.C(n_726),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_726),
.B(n_775),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_736),
.A2(n_787),
.B(n_777),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_781),
.A2(n_786),
.B(n_785),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_768),
.A2(n_707),
.B1(n_773),
.B2(n_696),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_670),
.A2(n_733),
.B(n_727),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_768),
.B(n_773),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_779),
.A2(n_789),
.B(n_784),
.C(n_780),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_756),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_791),
.B(n_793),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_788),
.Y(n_903)
);

AOI21x1_ASAP7_75t_L g904 ( 
.A1(n_696),
.A2(n_797),
.B(n_796),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_771),
.B(n_796),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_795),
.B(n_797),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_797),
.A2(n_763),
.B(n_731),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_747),
.A2(n_706),
.B(n_737),
.C(n_714),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_678),
.A2(n_718),
.B(n_715),
.C(n_674),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_763),
.A2(n_731),
.B(n_658),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_763),
.A2(n_731),
.B(n_658),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_763),
.A2(n_731),
.B(n_658),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_674),
.B(n_676),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_672),
.B(n_702),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_861),
.B(n_839),
.Y(n_915)
);

OAI21x1_ASAP7_75t_SL g916 ( 
.A1(n_904),
.A2(n_860),
.B(n_843),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_852),
.A2(n_879),
.B(n_859),
.C(n_834),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_839),
.B(n_825),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_864),
.B(n_857),
.Y(n_919)
);

AO31x2_ASAP7_75t_L g920 ( 
.A1(n_809),
.A2(n_865),
.A3(n_799),
.B(n_814),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_846),
.A2(n_899),
.B(n_828),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_806),
.B(n_810),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_914),
.B(n_897),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_885),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_858),
.B(n_862),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_840),
.B(n_863),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_895),
.A2(n_896),
.B(n_898),
.Y(n_927)
);

AO31x2_ASAP7_75t_L g928 ( 
.A1(n_819),
.A2(n_872),
.A3(n_881),
.B(n_883),
.Y(n_928)
);

AOI211x1_ASAP7_75t_L g929 ( 
.A1(n_826),
.A2(n_827),
.B(n_823),
.C(n_821),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_893),
.B(n_892),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_804),
.Y(n_931)
);

AO31x2_ASAP7_75t_L g932 ( 
.A1(n_815),
.A2(n_820),
.A3(n_891),
.B(n_836),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_803),
.B(n_807),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_L g934 ( 
.A(n_818),
.B(n_886),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_817),
.B(n_831),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_863),
.B(n_888),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_900),
.A2(n_808),
.B(n_905),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_871),
.B(n_812),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_878),
.Y(n_939)
);

AOI31xp67_ASAP7_75t_L g940 ( 
.A1(n_880),
.A2(n_869),
.A3(n_830),
.B(n_844),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_894),
.B(n_804),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_866),
.B(n_887),
.Y(n_942)
);

AOI221xp5_ASAP7_75t_SL g943 ( 
.A1(n_847),
.A2(n_853),
.B1(n_838),
.B2(n_873),
.C(n_833),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_870),
.A2(n_868),
.B(n_867),
.Y(n_944)
);

AO22x2_ASAP7_75t_L g945 ( 
.A1(n_800),
.A2(n_886),
.B1(n_854),
.B2(n_841),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_SL g946 ( 
.A1(n_832),
.A2(n_849),
.B(n_848),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_835),
.B(n_829),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_851),
.B(n_901),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_837),
.A2(n_876),
.B(n_874),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_798),
.B(n_822),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_824),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_903),
.B(n_851),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_866),
.B(n_902),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_850),
.Y(n_954)
);

BUFx5_ASAP7_75t_L g955 ( 
.A(n_906),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_851),
.A2(n_805),
.B1(n_801),
.B2(n_811),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_842),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_875),
.A2(n_877),
.B(n_882),
.Y(n_958)
);

OA22x2_ASAP7_75t_L g959 ( 
.A1(n_856),
.A2(n_884),
.B1(n_818),
.B2(n_855),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_889),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_809),
.A2(n_911),
.A3(n_912),
.B(n_910),
.Y(n_962)
);

OAI21x1_ASAP7_75t_SL g963 ( 
.A1(n_904),
.A2(n_860),
.B(n_913),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_913),
.B(n_672),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_913),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_816),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_909),
.A2(n_913),
.B(n_843),
.C(n_852),
.Y(n_967)
);

NAND3x1_ASAP7_75t_L g968 ( 
.A(n_856),
.B(n_623),
.C(n_711),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_913),
.B(n_813),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_913),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_913),
.B(n_813),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_910),
.A2(n_912),
.B(n_911),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_798),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_SL g974 ( 
.A(n_913),
.B(n_668),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_913),
.B(n_672),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_913),
.B(n_672),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_913),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_798),
.B(n_679),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_909),
.A2(n_913),
.B(n_843),
.C(n_852),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_913),
.B(n_813),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_913),
.B(n_813),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_913),
.B(n_672),
.Y(n_986)
);

OAI21x1_ASAP7_75t_SL g987 ( 
.A1(n_904),
.A2(n_860),
.B(n_913),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_913),
.B(n_845),
.Y(n_988)
);

NOR2x1_ASAP7_75t_SL g989 ( 
.A(n_913),
.B(n_851),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_910),
.A2(n_912),
.B(n_911),
.Y(n_990)
);

AO31x2_ASAP7_75t_L g991 ( 
.A1(n_809),
.A2(n_911),
.A3(n_912),
.B(n_910),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_SL g992 ( 
.A1(n_913),
.A2(n_860),
.B(n_909),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_822),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_913),
.B(n_813),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_913),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_816),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_913),
.B(n_813),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_798),
.B(n_679),
.Y(n_998)
);

AO21x1_ASAP7_75t_L g999 ( 
.A1(n_860),
.A2(n_907),
.B(n_904),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_913),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_913),
.B(n_813),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_798),
.B(n_679),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_L g1003 ( 
.A(n_813),
.B(n_913),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_890),
.B(n_909),
.C(n_808),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_913),
.B(n_813),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_798),
.B(n_679),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_910),
.A2(n_912),
.B(n_911),
.Y(n_1007)
);

OAI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_913),
.A2(n_802),
.B(n_879),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_798),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_816),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_910),
.A2(n_912),
.B(n_911),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_913),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_816),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_913),
.B(n_813),
.Y(n_1015)
);

AOI221xp5_ASAP7_75t_SL g1016 ( 
.A1(n_909),
.A2(n_908),
.B1(n_879),
.B2(n_808),
.C(n_847),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_913),
.B(n_668),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_834),
.A2(n_672),
.B(n_908),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_913),
.B(n_813),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_913),
.B(n_813),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_913),
.A2(n_802),
.B1(n_747),
.B2(n_706),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_816),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_816),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_913),
.B(n_813),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_798),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_913),
.B(n_672),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_913),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_913),
.B(n_672),
.Y(n_1029)
);

AO32x2_ASAP7_75t_L g1030 ( 
.A1(n_823),
.A2(n_854),
.A3(n_841),
.B1(n_858),
.B2(n_646),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_913),
.B(n_672),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_913),
.A2(n_911),
.B(n_910),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_913),
.A2(n_802),
.B(n_879),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_913),
.A2(n_802),
.B1(n_747),
.B2(n_706),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_925),
.A2(n_936),
.B1(n_1017),
.B2(n_974),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_1034),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_977),
.B(n_1027),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_993),
.Y(n_1039)
);

AO21x2_ASAP7_75t_L g1040 ( 
.A1(n_916),
.A2(n_987),
.B(n_963),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_976),
.B(n_986),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_970),
.B(n_979),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_SL g1043 ( 
.A1(n_934),
.A2(n_992),
.B(n_959),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_995),
.B(n_1000),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_988),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_969),
.B(n_971),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1021),
.A2(n_1035),
.B1(n_945),
.B2(n_931),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_974),
.A2(n_1017),
.B1(n_1018),
.B2(n_1003),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_961),
.A2(n_978),
.B(n_975),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1021),
.A2(n_1035),
.B1(n_945),
.B2(n_931),
.Y(n_1050)
);

OA21x2_ASAP7_75t_L g1051 ( 
.A1(n_990),
.A2(n_1011),
.B(n_1007),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_924),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_993),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_917),
.A2(n_980),
.A3(n_981),
.B(n_1028),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_924),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_951),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_1009),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_984),
.B(n_985),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_994),
.A2(n_1005),
.B1(n_1019),
.B2(n_1024),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_966),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_964),
.B(n_1029),
.Y(n_1062)
);

OR3x4_ASAP7_75t_SL g1063 ( 
.A(n_968),
.B(n_989),
.C(n_954),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_982),
.Y(n_1064)
);

OAI211xp5_ASAP7_75t_L g1065 ( 
.A1(n_997),
.A2(n_1020),
.B(n_1001),
.C(n_1015),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1012),
.A2(n_1032),
.B(n_983),
.Y(n_1066)
);

BUFx4_ASAP7_75t_SL g1067 ( 
.A(n_950),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_915),
.B(n_918),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1008),
.A2(n_1033),
.B1(n_923),
.B2(n_926),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_957),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_927),
.A2(n_944),
.B(n_921),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_972),
.A2(n_958),
.B(n_949),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_937),
.A2(n_1004),
.B(n_946),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_SL g1074 ( 
.A(n_942),
.B(n_919),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_941),
.B(n_933),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_L g1076 ( 
.A(n_952),
.B(n_948),
.Y(n_1076)
);

BUFx5_ASAP7_75t_L g1077 ( 
.A(n_939),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_951),
.B(n_996),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_922),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_930),
.B(n_996),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_998),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_1002),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_930),
.B(n_953),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_1006),
.B(n_1025),
.Y(n_1084)
);

AOI222xp33_ASAP7_75t_L g1085 ( 
.A1(n_935),
.A2(n_973),
.B1(n_956),
.B2(n_947),
.C1(n_938),
.C2(n_960),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1016),
.A2(n_943),
.B(n_940),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_929),
.B(n_955),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_991),
.B(n_920),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1022),
.A2(n_1023),
.B(n_1030),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1023),
.A2(n_920),
.B(n_928),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1010),
.B(n_1014),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_932),
.A2(n_928),
.B(n_955),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_955),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_965),
.B(n_970),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_965),
.B(n_970),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_R g1096 ( 
.A(n_965),
.B(n_856),
.Y(n_1096)
);

BUFx12f_ASAP7_75t_L g1097 ( 
.A(n_1034),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_925),
.A2(n_936),
.B1(n_863),
.B2(n_974),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1013),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_967),
.A2(n_983),
.B(n_917),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1013),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_965),
.B(n_970),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_999),
.A2(n_917),
.A3(n_809),
.B(n_961),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_965),
.B(n_970),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_977),
.B(n_1027),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_965),
.B(n_970),
.Y(n_1106)
);

CKINVDCx6p67_ASAP7_75t_R g1107 ( 
.A(n_1037),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1067),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1078),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1099),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1060),
.B(n_1046),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1077),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_1067),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1055),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1065),
.A2(n_1062),
.B(n_1059),
.C(n_1036),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1059),
.B(n_1062),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1078),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1077),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1079),
.B(n_1065),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1087),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1086),
.A2(n_1071),
.B(n_1100),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1055),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1049),
.A2(n_1066),
.B(n_1072),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_1045),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1073),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1068),
.B(n_1104),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1073),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1041),
.B(n_1053),
.Y(n_1128)
);

AO21x2_ASAP7_75t_L g1129 ( 
.A1(n_1049),
.A2(n_1066),
.B(n_1090),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1101),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1093),
.B(n_1091),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1042),
.A2(n_1095),
.B(n_1094),
.C(n_1106),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1044),
.B(n_1094),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1051),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1101),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1091),
.B(n_1089),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1047),
.B(n_1050),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_1097),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_SL g1139 ( 
.A(n_1039),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1044),
.B(n_1095),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1061),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1048),
.A2(n_1036),
.B(n_1098),
.Y(n_1142)
);

NAND4xp25_ASAP7_75t_SL g1143 ( 
.A(n_1098),
.B(n_1085),
.C(n_1076),
.D(n_1102),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_L g1144 ( 
.A(n_1141),
.B(n_1057),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1111),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1129),
.B(n_1120),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1118),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1129),
.B(n_1088),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1134),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1129),
.B(n_1092),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1111),
.B(n_1103),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1112),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1137),
.B(n_1119),
.Y(n_1154)
);

INVx4_ASAP7_75t_R g1155 ( 
.A(n_1108),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1136),
.B(n_1040),
.Y(n_1156)
);

AND2x4_ASAP7_75t_SL g1157 ( 
.A(n_1131),
.B(n_1080),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1131),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1140),
.B(n_1069),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1121),
.B(n_1040),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1150),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_1158),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1144),
.B(n_1109),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1146),
.B(n_1137),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1152),
.B(n_1123),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1152),
.B(n_1123),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1149),
.B(n_1123),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1146),
.B(n_1128),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_1158),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1156),
.B(n_1114),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_1157),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1153),
.B(n_1115),
.C(n_1085),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1151),
.B(n_1122),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1145),
.B(n_1159),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1148),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1157),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1158),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1161),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1174),
.B(n_1147),
.Y(n_1179)
);

OR3x2_ASAP7_75t_L g1180 ( 
.A(n_1168),
.B(n_1155),
.C(n_1107),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1174),
.B(n_1154),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1165),
.B(n_1166),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1172),
.A2(n_1132),
.B(n_1133),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_L g1184 ( 
.A(n_1163),
.B(n_1158),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1170),
.B(n_1156),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1161),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1165),
.B(n_1166),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1165),
.B(n_1160),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1175),
.Y(n_1189)
);

BUFx2_ASAP7_75t_SL g1190 ( 
.A(n_1171),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1166),
.B(n_1160),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1173),
.B(n_1147),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1167),
.B(n_1160),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1190),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1182),
.B(n_1167),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1182),
.B(n_1164),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1178),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_1180),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1178),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1193),
.B(n_1179),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1186),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1190),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1187),
.B(n_1167),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1189),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1184),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1193),
.B(n_1179),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1204),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1202),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1195),
.B(n_1187),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1198),
.Y(n_1210)
);

AOI21xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1205),
.A2(n_1180),
.B(n_1155),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1197),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1198),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1195),
.B(n_1193),
.Y(n_1214)
);

OAI32xp33_ASAP7_75t_L g1215 ( 
.A1(n_1198),
.A2(n_1176),
.A3(n_1171),
.B1(n_1180),
.B2(n_1113),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1198),
.A2(n_1184),
.B(n_1163),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1196),
.Y(n_1217)
);

OAI31xp33_ASAP7_75t_L g1218 ( 
.A1(n_1205),
.A2(n_1172),
.A3(n_1176),
.B(n_1143),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1196),
.B(n_1188),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1197),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_1194),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1199),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1203),
.A2(n_1142),
.B1(n_1183),
.B2(n_1126),
.Y(n_1223)
);

AOI211xp5_ASAP7_75t_L g1224 ( 
.A1(n_1200),
.A2(n_1183),
.B(n_1142),
.C(n_1096),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1223),
.A2(n_1191),
.B1(n_1188),
.B2(n_1185),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1207),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1210),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1210),
.A2(n_1206),
.B1(n_1203),
.B2(n_1162),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1213),
.Y(n_1229)
);

OAI21xp33_ASAP7_75t_L g1230 ( 
.A1(n_1223),
.A2(n_1213),
.B(n_1221),
.Y(n_1230)
);

OAI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1218),
.A2(n_1181),
.B1(n_1164),
.B2(n_1168),
.C(n_1189),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_L g1232 ( 
.A(n_1213),
.B(n_1083),
.C(n_1116),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1211),
.A2(n_1162),
.B1(n_1181),
.B2(n_1107),
.Y(n_1233)
);

AOI32xp33_ASAP7_75t_L g1234 ( 
.A1(n_1224),
.A2(n_1188),
.A3(n_1191),
.B1(n_1177),
.B2(n_1169),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1233),
.A2(n_1215),
.B(n_1216),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1226),
.Y(n_1236)
);

OAI211xp5_ASAP7_75t_L g1237 ( 
.A1(n_1230),
.A2(n_1215),
.B(n_1096),
.C(n_1211),
.Y(n_1237)
);

AOI211xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1231),
.A2(n_1208),
.B(n_1139),
.C(n_1217),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1225),
.A2(n_1219),
.B1(n_1209),
.B2(n_1214),
.Y(n_1239)
);

OAI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1234),
.A2(n_1214),
.B(n_1212),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1229),
.B(n_1227),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1228),
.A2(n_1209),
.B(n_1212),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1232),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1230),
.A2(n_1043),
.B(n_1222),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1231),
.A2(n_1220),
.B1(n_1222),
.B2(n_1191),
.Y(n_1245)
);

OA211x2_ASAP7_75t_L g1246 ( 
.A1(n_1230),
.A2(n_1074),
.B(n_1063),
.C(n_1083),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1238),
.B(n_1110),
.C(n_1220),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_L g1248 ( 
.A(n_1237),
.B(n_1244),
.C(n_1243),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1236),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1245),
.B(n_1199),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1235),
.B(n_1138),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1241),
.B(n_1192),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_L g1253 ( 
.A(n_1240),
.B(n_1058),
.C(n_1081),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1242),
.Y(n_1254)
);

NAND4xp25_ASAP7_75t_L g1255 ( 
.A(n_1251),
.B(n_1246),
.C(n_1239),
.D(n_1064),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1248),
.B(n_1056),
.C(n_1052),
.Y(n_1256)
);

NOR3xp33_ASAP7_75t_L g1257 ( 
.A(n_1248),
.B(n_1082),
.C(n_1057),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_SL g1258 ( 
.A(n_1254),
.B(n_1063),
.C(n_1075),
.Y(n_1258)
);

NOR2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1247),
.B(n_1054),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_SL g1260 ( 
.A(n_1249),
.B(n_1084),
.Y(n_1260)
);

NOR2x1_ASAP7_75t_L g1261 ( 
.A(n_1252),
.B(n_1070),
.Y(n_1261)
);

NOR2x1_ASAP7_75t_L g1262 ( 
.A(n_1250),
.B(n_1109),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1256),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1255),
.B(n_1253),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_SL g1265 ( 
.A(n_1258),
.B(n_1124),
.Y(n_1265)
);

NOR3xp33_ASAP7_75t_L g1266 ( 
.A(n_1257),
.B(n_1056),
.C(n_1052),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_1259),
.B(n_1201),
.Y(n_1267)
);

NOR2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1261),
.B(n_1109),
.Y(n_1268)
);

NAND3xp33_ASAP7_75t_SL g1269 ( 
.A(n_1260),
.B(n_1105),
.C(n_1038),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1263),
.B(n_1201),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1269),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1266),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1268),
.Y(n_1273)
);

OAI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1273),
.A2(n_1265),
.B1(n_1264),
.B2(n_1267),
.C(n_1271),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1273),
.A2(n_1262),
.B1(n_1080),
.B2(n_1126),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1274),
.A2(n_1272),
.B(n_1270),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1276),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1277),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1278),
.B(n_1276),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1279),
.B(n_1117),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1280),
.B(n_1117),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1281),
.A2(n_1275),
.B1(n_1135),
.B2(n_1130),
.Y(n_1282)
);


endmodule