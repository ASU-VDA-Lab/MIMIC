module fake_jpeg_18611_n_295 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_295);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_41),
.B1(n_42),
.B2(n_27),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_26),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_25),
.B1(n_13),
.B2(n_12),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_31),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_31),
.C(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_58),
.B(n_62),
.Y(n_74)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_61),
.B1(n_43),
.B2(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_34),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_31),
.B(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_31),
.C(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_38),
.B1(n_44),
.B2(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_56),
.B1(n_44),
.B2(n_60),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_85),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_64),
.C(n_62),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_31),
.C(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_74),
.B1(n_86),
.B2(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_47),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_100),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_85),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_56),
.B1(n_44),
.B2(n_59),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_105),
.B1(n_48),
.B2(n_72),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_31),
.B(n_32),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_68),
.B1(n_72),
.B2(n_78),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_61),
.B1(n_52),
.B2(n_55),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_40),
.B1(n_35),
.B2(n_36),
.Y(n_122)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_45),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_40),
.B1(n_29),
.B2(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_78),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_66),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_83),
.B(n_73),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_123),
.B1(n_124),
.B2(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_40),
.B1(n_72),
.B2(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_122),
.B1(n_101),
.B2(n_67),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_41),
.B1(n_42),
.B2(n_35),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_45),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_45),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_47),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_91),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_102),
.B1(n_93),
.B2(n_96),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_140),
.B1(n_146),
.B2(n_33),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_47),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_139),
.B1(n_151),
.B2(n_118),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_90),
.C(n_100),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_144),
.C(n_110),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_103),
.B1(n_105),
.B2(n_88),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_127),
.B1(n_115),
.B2(n_112),
.Y(n_140)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_100),
.C(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_34),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_150),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_28),
.B1(n_27),
.B2(n_30),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_153),
.B1(n_30),
.B2(n_28),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_50),
.B1(n_48),
.B2(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_76),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_175),
.B1(n_178),
.B2(n_180),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_108),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_164),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_115),
.C(n_128),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_170),
.C(n_177),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_126),
.B(n_113),
.C(n_130),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_16),
.B(n_12),
.C(n_22),
.Y(n_205)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_183),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_131),
.A2(n_121),
.B1(n_33),
.B2(n_30),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_47),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_139),
.B1(n_144),
.B2(n_137),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_121),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_182),
.C(n_63),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_121),
.C(n_63),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_137),
.B(n_147),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_202),
.B(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_28),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_204),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_53),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_174),
.B1(n_168),
.B2(n_175),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_220),
.B1(n_185),
.B2(n_192),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_179),
.B1(n_158),
.B2(n_164),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_219),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_177),
.B1(n_160),
.B2(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_226),
.B1(n_187),
.B2(n_185),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_163),
.B1(n_13),
.B2(n_14),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_14),
.B1(n_19),
.B2(n_22),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_12),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_194),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_188),
.A2(n_19),
.B1(n_22),
.B2(n_16),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_22),
.B1(n_16),
.B2(n_3),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_24),
.C(n_15),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_223),
.C(n_189),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_16),
.B1(n_15),
.B2(n_3),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_24),
.C(n_15),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_229),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_236),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_190),
.C(n_193),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_186),
.C(n_24),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_237),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_187),
.B1(n_207),
.B2(n_206),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_239),
.B1(n_223),
.B2(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_198),
.B1(n_199),
.B2(n_205),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_210),
.C(n_214),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_205),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_220),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_250),
.B(n_242),
.Y(n_257)
);

OAI322xp33_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_186),
.A3(n_24),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_1),
.B(n_2),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_24),
.C(n_5),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_262),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_240),
.B1(n_231),
.B2(n_238),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_232),
.C(n_8),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_265),
.C(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_6),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_6),
.C(n_8),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_6),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_8),
.C(n_9),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_259),
.C(n_10),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_8),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_256),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_257),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_265),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_272),
.C(n_277),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_268),
.B(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_282),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_280),
.C(n_283),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_288),
.B(n_10),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_9),
.C(n_10),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_292),
.B(n_9),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_11),
.B(n_290),
.C(n_271),
.D(n_287),
.Y(n_295)
);


endmodule