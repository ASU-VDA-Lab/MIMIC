module fake_jpeg_31785_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_53),
.Y(n_80)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_52),
.Y(n_71)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_26),
.B(n_28),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_1),
.C(n_2),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_36),
.B1(n_22),
.B2(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_79),
.B1(n_34),
.B2(n_16),
.Y(n_99)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_13),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_76),
.B1(n_32),
.B2(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_31),
.B1(n_49),
.B2(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_22),
.B1(n_32),
.B2(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_16),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_92),
.Y(n_120)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_24),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_16),
.B(n_32),
.C(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_44),
.B1(n_33),
.B2(n_35),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_66),
.B1(n_67),
.B2(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_10),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_74),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_R g117 ( 
.A(n_100),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_11),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_34),
.Y(n_102)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_76),
.C(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_70),
.B1(n_74),
.B2(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_9),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_12),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_57),
.B(n_10),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_87),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_130),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_135),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_126),
.B1(n_133),
.B2(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_70),
.B(n_67),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_85),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_98),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_6),
.B1(n_66),
.B2(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_6),
.B1(n_94),
.B2(n_112),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_103),
.B1(n_113),
.B2(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_6),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_88),
.Y(n_159)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_101),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_137),
.C(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_156),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_152),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_113),
.B1(n_123),
.B2(n_91),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_119),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_90),
.B(n_103),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_161),
.B(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_141),
.Y(n_178)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_155),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_88),
.B(n_127),
.C(n_124),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_122),
.B1(n_136),
.B2(n_127),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_172),
.B(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_122),
.B1(n_133),
.B2(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_171),
.B1(n_148),
.B2(n_160),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_169),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_121),
.B1(n_129),
.B2(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_161),
.B(n_144),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_146),
.C(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_178),
.C(n_145),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_181),
.C(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_142),
.C(n_150),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_156),
.B1(n_152),
.B2(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_187),
.B1(n_162),
.B2(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_142),
.B1(n_148),
.B2(n_149),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_162),
.B1(n_170),
.B2(n_168),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_171),
.B(n_164),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_190),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_196),
.B(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_169),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_181),
.C(n_180),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.C(n_198),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_172),
.C(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_200),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_184),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_195),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_188),
.A3(n_191),
.B(n_165),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_192),
.C(n_185),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_199),
.B(n_200),
.Y(n_212)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_203),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_218),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_216),
.C(n_215),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_204),
.C(n_194),
.Y(n_220)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_221),
.B(n_211),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_194),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

OAI221xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_202),
.B1(n_223),
.B2(n_215),
.C(n_196),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_173),
.Y(n_226)
);


endmodule