module fake_jpeg_280_n_655 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_655);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_655;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_67),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_79),
.Y(n_171)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_8),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_86),
.A2(n_58),
.B(n_20),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_8),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_33),
.Y(n_141)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

BUFx2_ASAP7_75t_R g153 ( 
.A(n_114),
.Y(n_153)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_117),
.B(n_118),
.Y(n_197)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_54),
.Y(n_125)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_59),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_127),
.B(n_143),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_159),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_47),
.B1(n_57),
.B2(n_55),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_136),
.A2(n_142),
.B1(n_165),
.B2(n_19),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_141),
.B(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_64),
.A2(n_57),
.B1(n_53),
.B2(n_33),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_59),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_30),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_146),
.B(n_152),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_30),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_68),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_72),
.A2(n_33),
.B1(n_57),
.B2(n_50),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_77),
.A2(n_53),
.B1(n_19),
.B2(n_50),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_166),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_73),
.B(n_58),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_82),
.B(n_37),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_183),
.B(n_185),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_67),
.B(n_54),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_79),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_83),
.B(n_37),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_117),
.B(n_40),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_84),
.B(n_45),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_87),
.A2(n_98),
.B1(n_99),
.B2(n_113),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_50),
.B1(n_19),
.B2(n_166),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_100),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_36),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_67),
.B(n_36),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_123),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_111),
.B1(n_107),
.B2(n_112),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_208),
.A2(n_216),
.B1(n_223),
.B2(n_247),
.Y(n_330)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_212),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_213),
.Y(n_285)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_228),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_171),
.A2(n_34),
.B1(n_31),
.B2(n_38),
.Y(n_216)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_221),
.B(n_250),
.Y(n_297)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_171),
.A2(n_38),
.B1(n_34),
.B2(n_45),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_225),
.Y(n_319)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_227),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_126),
.B(n_133),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_229),
.Y(n_307)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_132),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_245),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_234),
.B(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_236),
.A2(n_276),
.B1(n_189),
.B2(n_195),
.Y(n_293)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

INVx4_ASAP7_75t_SL g238 ( 
.A(n_140),
.Y(n_238)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

OA22x2_ASAP7_75t_L g326 ( 
.A1(n_239),
.A2(n_277),
.B1(n_0),
.B2(n_1),
.Y(n_326)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_240),
.Y(n_332)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_241),
.Y(n_346)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_182),
.A2(n_53),
.B1(n_20),
.B2(n_40),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_273),
.B1(n_164),
.B2(n_195),
.Y(n_288)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_135),
.B(n_65),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_139),
.B(n_94),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_246),
.B(n_0),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_197),
.A2(n_90),
.B1(n_115),
.B2(n_105),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_200),
.Y(n_250)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_167),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_251),
.A2(n_255),
.B1(n_260),
.B2(n_264),
.Y(n_336)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_158),
.Y(n_252)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_252),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_253),
.Y(n_337)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_254),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_197),
.A2(n_118),
.B1(n_104),
.B2(n_101),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_258),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_263),
.Y(n_324)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_144),
.B(n_44),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_267),
.C(n_270),
.Y(n_292)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_147),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_134),
.A2(n_35),
.B1(n_8),
.B2(n_9),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_265),
.B(n_269),
.Y(n_329)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_266),
.B(n_272),
.Y(n_348)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_145),
.B(n_0),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_268),
.B(n_275),
.Y(n_305)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_147),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_149),
.B(n_193),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_162),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_271),
.B(n_274),
.Y(n_341)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_174),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_166),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_129),
.Y(n_275)
);

BUFx6f_ASAP7_75t_SL g276 ( 
.A(n_175),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_134),
.A2(n_7),
.B1(n_17),
.B2(n_15),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_206),
.B1(n_157),
.B2(n_177),
.Y(n_296)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_151),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_279),
.B(n_280),
.Y(n_343)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_155),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_165),
.B(n_6),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_137),
.C(n_161),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_131),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_282),
.B(n_283),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_164),
.A2(n_6),
.B(n_17),
.C(n_13),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_209),
.A2(n_206),
.B(n_179),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_284),
.B(n_326),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_288),
.A2(n_301),
.B1(n_304),
.B2(n_311),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_293),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_162),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_299),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_151),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_168),
.B1(n_192),
.B2(n_190),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_239),
.A2(n_168),
.B1(n_192),
.B2(n_190),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_189),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_315),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_137),
.B1(n_161),
.B2(n_198),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_254),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_218),
.B(n_158),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_211),
.B(n_174),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_317),
.B(n_320),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_229),
.B(n_177),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_277),
.A2(n_198),
.B1(n_175),
.B2(n_172),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_328),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_220),
.A2(n_224),
.B1(n_228),
.B2(n_230),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_245),
.A2(n_172),
.B1(n_1),
.B2(n_2),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_245),
.A2(n_262),
.B1(n_208),
.B2(n_229),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_334),
.B(n_344),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_11),
.C(n_17),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_340),
.C(n_347),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_217),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_338),
.A2(n_339),
.B1(n_276),
.B2(n_238),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_232),
.A2(n_3),
.B1(n_4),
.B2(n_18),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_232),
.B(n_11),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_4),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_270),
.B(n_11),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_316),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_350),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_309),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_317),
.B(n_225),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_351),
.B(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_343),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_284),
.A2(n_215),
.B(n_227),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_356),
.A2(n_375),
.B(n_392),
.Y(n_437)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_307),
.A2(n_270),
.B1(n_279),
.B2(n_269),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_366),
.A2(n_378),
.B1(n_398),
.B2(n_339),
.Y(n_428)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_368),
.B(n_369),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_290),
.B(n_258),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_379),
.Y(n_410)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_328),
.A2(n_263),
.B1(n_240),
.B2(n_241),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_387),
.B1(n_303),
.B2(n_342),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_327),
.A2(n_259),
.B(n_242),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_377),
.A2(n_333),
.B1(n_302),
.B2(n_345),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_307),
.A2(n_219),
.B1(n_214),
.B2(n_222),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_315),
.B(n_256),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_381),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_308),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_295),
.B(n_248),
.Y(n_382)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_389),
.B(n_400),
.Y(n_417)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_386),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_384),
.B(n_289),
.Y(n_440)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_304),
.A2(n_237),
.B1(n_210),
.B2(n_282),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_298),
.B(n_252),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_394),
.C(n_340),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_321),
.A2(n_271),
.B1(n_272),
.B2(n_266),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_294),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_396),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_308),
.A2(n_226),
.B(n_244),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_393),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_292),
.B(n_233),
.C(n_248),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_341),
.Y(n_395)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_305),
.B(n_13),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_308),
.A2(n_251),
.B(n_260),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_397),
.A2(n_320),
.B(n_330),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_299),
.A2(n_4),
.B1(n_18),
.B2(n_306),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_334),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_347),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_311),
.A2(n_4),
.B1(n_18),
.B2(n_288),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_371),
.A2(n_344),
.B1(n_297),
.B2(n_301),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_402),
.A2(n_423),
.B(n_427),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_292),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_405),
.C(n_408),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_404),
.B(n_431),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_388),
.C(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

OA22x2_ASAP7_75t_L g411 ( 
.A1(n_357),
.A2(n_326),
.B1(n_336),
.B2(n_319),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_411),
.B(n_369),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_367),
.A2(n_326),
.B1(n_312),
.B2(n_319),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_415),
.A2(n_420),
.B1(n_398),
.B2(n_366),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_367),
.A2(n_326),
.B1(n_300),
.B2(n_325),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_356),
.A2(n_335),
.B(n_337),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_371),
.A2(n_337),
.B(n_300),
.Y(n_427)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_429),
.B(n_414),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_357),
.A2(n_338),
.B1(n_325),
.B2(n_286),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_430),
.A2(n_434),
.B1(n_443),
.B2(n_363),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_371),
.A2(n_303),
.B(n_323),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_375),
.A2(n_318),
.B(n_314),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_432),
.A2(n_397),
.B(n_379),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_342),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_436),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_372),
.A2(n_318),
.B1(n_286),
.B2(n_302),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_333),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_438),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_393),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_368),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_442),
.C(n_392),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_285),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_372),
.A2(n_286),
.B1(n_287),
.B2(n_289),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_287),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_353),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_376),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_446),
.B(n_458),
.C(n_464),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_401),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_447),
.B(n_448),
.Y(n_519)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_385),
.C(n_351),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_442),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_451),
.B(n_437),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_454),
.A2(n_467),
.B1(n_468),
.B2(n_473),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_456),
.A2(n_469),
.B(n_475),
.Y(n_492)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_401),
.Y(n_457)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_362),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_444),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_462),
.Y(n_503)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_463),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_405),
.B(n_385),
.C(n_395),
.Y(n_464)
);

AOI21xp33_ASAP7_75t_L g465 ( 
.A1(n_413),
.A2(n_359),
.B(n_352),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_465),
.A2(n_422),
.B(n_419),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_407),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_466),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_406),
.B(n_349),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_427),
.A2(n_374),
.B(n_354),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_410),
.Y(n_472)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_420),
.A2(n_415),
.B1(n_430),
.B2(n_431),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_414),
.A2(n_399),
.B1(n_363),
.B2(n_378),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_436),
.B(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_476),
.Y(n_518)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_477),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_407),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_478),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_386),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_479),
.Y(n_516)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_426),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_480),
.A2(n_481),
.B1(n_421),
.B2(n_412),
.Y(n_510)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_445),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_364),
.Y(n_482)
);

NAND4xp25_ASAP7_75t_SL g493 ( 
.A(n_482),
.B(n_483),
.C(n_443),
.D(n_434),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_419),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_484),
.A2(n_409),
.B(n_411),
.C(n_423),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_455),
.A2(n_404),
.B1(n_424),
.B2(n_417),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_487),
.A2(n_501),
.B1(n_488),
.B2(n_490),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_511),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_493),
.Y(n_534)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_458),
.B(n_429),
.Y(n_497)
);

XNOR2x2_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_514),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_453),
.A2(n_437),
.B(n_402),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_498),
.A2(n_478),
.B(n_479),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_505),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_452),
.B1(n_484),
.B2(n_473),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_449),
.B(n_435),
.C(n_406),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_507),
.C(n_508),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_456),
.C(n_453),
.Y(n_528)
);

XNOR2x1_ASAP7_75t_L g505 ( 
.A(n_450),
.B(n_411),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_452),
.A2(n_454),
.B1(n_447),
.B2(n_457),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_506),
.A2(n_513),
.B1(n_468),
.B2(n_477),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_449),
.B(n_419),
.C(n_439),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_450),
.B(n_416),
.C(n_422),
.Y(n_508)
);

XNOR2x1_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_411),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_471),
.Y(n_532)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_416),
.C(n_432),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_481),
.A2(n_428),
.B1(n_424),
.B2(n_411),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_471),
.B(n_421),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_412),
.C(n_425),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_517),
.B(n_482),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_483),
.Y(n_522)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_522),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_523),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_502),
.B(n_472),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_524),
.B(n_526),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_462),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_466),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_530),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_528),
.A2(n_536),
.B(n_537),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_519),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_532),
.B(n_498),
.Y(n_568)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_519),
.Y(n_533)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_533),
.Y(n_574)
);

OAI22x1_ASAP7_75t_L g535 ( 
.A1(n_501),
.A2(n_475),
.B1(n_470),
.B2(n_461),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_535),
.A2(n_545),
.B1(n_513),
.B2(n_489),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_492),
.A2(n_470),
.B(n_469),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_547),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_486),
.B(n_459),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_550),
.Y(n_551)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_510),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_541),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_503),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_543),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_500),
.B(n_460),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_504),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_492),
.Y(n_563)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_495),
.Y(n_546)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_546),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_518),
.B(n_459),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_516),
.A2(n_470),
.B1(n_467),
.B2(n_448),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_548),
.A2(n_506),
.B1(n_518),
.B2(n_488),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_549),
.A2(n_496),
.B1(n_515),
.B2(n_495),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_486),
.B(n_480),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_553),
.A2(n_555),
.B1(n_558),
.B2(n_562),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_517),
.C(n_511),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_560),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_522),
.A2(n_536),
.B(n_537),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_557),
.B(n_523),
.C(n_531),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_545),
.A2(n_490),
.B1(n_487),
.B2(n_494),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_539),
.B(n_499),
.C(n_508),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_549),
.A2(n_534),
.B1(n_525),
.B2(n_548),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_563),
.B(n_565),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_550),
.B(n_505),
.C(n_514),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_521),
.B(n_509),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_567),
.B(n_568),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_521),
.B(n_491),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_570),
.B(n_571),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_540),
.B(n_497),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_575),
.A2(n_576),
.B1(n_533),
.B2(n_546),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_534),
.A2(n_515),
.B1(n_474),
.B2(n_463),
.Y(n_576)
);

BUFx24_ASAP7_75t_SL g578 ( 
.A(n_566),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_578),
.B(n_591),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_572),
.B(n_538),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_580),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_529),
.C(n_532),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_551),
.B(n_560),
.C(n_529),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_583),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_582),
.A2(n_588),
.B(n_598),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_541),
.C(n_531),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_584),
.Y(n_600)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_556),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_585),
.B(n_586),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_570),
.C(n_565),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_562),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_564),
.A2(n_525),
.B(n_574),
.Y(n_588)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_569),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_575),
.A2(n_535),
.B1(n_547),
.B2(n_520),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_592),
.A2(n_597),
.B1(n_598),
.B2(n_596),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_573),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_593),
.B(n_588),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_559),
.B(n_425),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_594),
.B(n_355),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_561),
.A2(n_520),
.B1(n_493),
.B2(n_387),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_564),
.A2(n_418),
.B(n_358),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_599),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_559),
.C(n_561),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_601),
.B(n_606),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_583),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_610),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_561),
.C(n_553),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_580),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_596),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_595),
.B(n_558),
.C(n_567),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_609),
.B(n_613),
.C(n_603),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_593),
.A2(n_569),
.B1(n_555),
.B2(n_576),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_611),
.A2(n_616),
.B1(n_587),
.B2(n_597),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_377),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_595),
.B(n_568),
.C(n_418),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_589),
.A2(n_383),
.B(n_360),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_615),
.A2(n_291),
.B(n_345),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_617),
.B(n_622),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_618),
.B(n_620),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_614),
.A2(n_586),
.B(n_589),
.Y(n_620)
);

INVxp33_ASAP7_75t_L g637 ( 
.A(n_621),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_373),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_602),
.B(n_291),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_624),
.B(n_628),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_625),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_605),
.B(n_4),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_627),
.Y(n_639)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_604),
.A2(n_601),
.B(n_606),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_629),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_599),
.B(n_609),
.C(n_613),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_630),
.B(n_610),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_629),
.B(n_608),
.Y(n_631)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_631),
.Y(n_643)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_634),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_619),
.B(n_600),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_638),
.B(n_630),
.Y(n_642)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_640),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_641),
.B(n_642),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_636),
.B(n_619),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_644),
.B(n_645),
.C(n_640),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_639),
.B(n_626),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_647),
.B(n_648),
.C(n_646),
.Y(n_650)
);

OAI311xp33_ASAP7_75t_L g648 ( 
.A1(n_641),
.A2(n_623),
.A3(n_633),
.B1(n_632),
.C1(n_617),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_650),
.B(n_651),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_647),
.B(n_643),
.C(n_623),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_649),
.C(n_635),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_637),
.C(n_621),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_654),
.B(n_622),
.Y(n_655)
);


endmodule