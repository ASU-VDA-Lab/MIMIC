module fake_netlist_6_3922_n_1978 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1978);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1978;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_1970;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_231),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_198),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_103),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_252),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_329),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_328),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_189),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_235),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_162),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_392),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_214),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_68),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_303),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_224),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_495),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_481),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_234),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_429),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_71),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_331),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_485),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_353),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_102),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_157),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_384),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_428),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_39),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_382),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_29),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_248),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_317),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_76),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_337),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_446),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_245),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_37),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_199),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_113),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_500),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_227),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_1),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_34),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_298),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_435),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_83),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_44),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_217),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_265),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_251),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_395),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_162),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_355),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_98),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_318),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_158),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_387),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_0),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_206),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_349),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_326),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_402),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_399),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_400),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_76),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_299),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_362),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_301),
.Y(n_578)
);

BUFx2_ASAP7_75t_SL g579 ( 
.A(n_20),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_70),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_479),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_383),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_122),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_480),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_398),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_499),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_51),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_177),
.Y(n_588)
);

BUFx5_ASAP7_75t_L g589 ( 
.A(n_221),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_397),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_4),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_357),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_474),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_149),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_394),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_233),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_82),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_109),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_35),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_99),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_339),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_292),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_493),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_309),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_6),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_267),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_273),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_413),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_270),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_406),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_322),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_268),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_255),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_361),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_360),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_79),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_38),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_489),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_53),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_332),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_390),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_265),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_409),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_178),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_458),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_294),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_116),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_344),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_63),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_125),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_483),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_173),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_10),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_248),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_263),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_186),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_285),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_219),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_222),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_23),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_192),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_187),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_244),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_295),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_62),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_304),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_347),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_386),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_235),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_165),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_74),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_27),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_230),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_150),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_0),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_155),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_281),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_330),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_312),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_153),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_112),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_482),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_351),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_238),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_31),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_420),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_257),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_214),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_216),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_359),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_130),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_391),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_228),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_507),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_501),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_217),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_449),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_323),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_87),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_198),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_171),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_68),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_146),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_13),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_277),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_358),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_363),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_340),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_117),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_112),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_46),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_502),
.Y(n_692)
);

BUFx10_ASAP7_75t_L g693 ( 
.A(n_92),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_336),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_41),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_354),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_192),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_64),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_468),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_424),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_174),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_403),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_103),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_24),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_155),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_102),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_587),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_589),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_589),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_589),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

CKINVDCx16_ASAP7_75t_R g713 ( 
.A(n_511),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_513),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_535),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_536),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_512),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_589),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_544),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_554),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_512),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_551),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_589),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_520),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_698),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_536),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_520),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_629),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_681),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_629),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_633),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_633),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_682),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_703),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_592),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_548),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_703),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_592),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_681),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_561),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_563),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_681),
.Y(n_742)
);

INVxp33_ASAP7_75t_SL g743 ( 
.A(n_695),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_681),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_510),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_516),
.Y(n_746)
);

CKINVDCx14_ASAP7_75t_R g747 ( 
.A(n_599),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_704),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_548),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_571),
.Y(n_750)
);

INVxp33_ASAP7_75t_SL g751 ( 
.A(n_525),
.Y(n_751)
);

INVxp33_ASAP7_75t_SL g752 ( 
.A(n_525),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_650),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_650),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_565),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_517),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_572),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_546),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_693),
.Y(n_759)
);

INVxp33_ASAP7_75t_L g760 ( 
.A(n_546),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_676),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_676),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_519),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_522),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_527),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_533),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_581),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_701),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_602),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_684),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_540),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_580),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_542),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_684),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_509),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_514),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_518),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_693),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_552),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_558),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_559),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_530),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_602),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_598),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_574),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_600),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_576),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_581),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_606),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_693),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_619),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_649),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_664),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_534),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_669),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_783),
.Y(n_796)
);

CKINVDCx6p67_ASAP7_75t_R g797 ( 
.A(n_713),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_729),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_735),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_729),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_767),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_739),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_767),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_767),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_767),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_708),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_743),
.A2(n_543),
.B1(n_573),
.B2(n_529),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_747),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_709),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_783),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_710),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_717),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_SL g813 ( 
.A1(n_717),
.A2(n_543),
.B1(n_573),
.B2(n_529),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_711),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_712),
.A2(n_608),
.B(n_582),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_718),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_723),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_778),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_744),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_758),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_758),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_788),
.Y(n_823)
);

NOR2x1_ASAP7_75t_L g824 ( 
.A(n_788),
.B(n_538),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_725),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_788),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_735),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_772),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_735),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_716),
.B(n_652),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_721),
.A2(n_646),
.B1(n_706),
.B2(n_701),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_714),
.B(n_526),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_775),
.B(n_776),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_735),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_738),
.Y(n_836)
);

CKINVDCx8_ASAP7_75t_R g837 ( 
.A(n_722),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_748),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_745),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_746),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_777),
.B(n_782),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_768),
.A2(n_646),
.B1(n_515),
.B2(n_532),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_756),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_763),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_715),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_764),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_SL g847 ( 
.A1(n_721),
.A2(n_706),
.B1(n_537),
.B2(n_630),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_738),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_765),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_766),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_768),
.A2(n_539),
.B1(n_545),
.B2(n_508),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_771),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_719),
.B(n_526),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_773),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_800),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_831),
.B(n_582),
.Y(n_856)
);

AND3x1_ASAP7_75t_L g857 ( 
.A(n_842),
.B(n_652),
.C(n_671),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_830),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_834),
.A2(n_740),
.B1(n_741),
.B2(n_720),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_834),
.B(n_755),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_835),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_800),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_801),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_836),
.B(n_726),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_835),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_806),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_806),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_809),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_801),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_815),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_817),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_836),
.B(n_779),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_818),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_821),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_SL g875 ( 
.A1(n_832),
.A2(n_749),
.B1(n_753),
.B2(n_736),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_811),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_834),
.B(n_608),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_821),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_827),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_799),
.B(n_780),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_799),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_807),
.A2(n_749),
.B1(n_753),
.B2(n_736),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_821),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_821),
.Y(n_884)
);

BUFx6f_ASAP7_75t_SL g885 ( 
.A(n_848),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_839),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_821),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_847),
.A2(n_761),
.B1(n_762),
.B2(n_754),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_839),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_825),
.B(n_747),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_840),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_SL g892 ( 
.A(n_831),
.B(n_707),
.Y(n_892)
);

XOR2xp5_ASAP7_75t_L g893 ( 
.A(n_838),
.B(n_754),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_848),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_798),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_840),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_841),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_841),
.B(n_844),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_841),
.B(n_853),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_833),
.B(n_757),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_824),
.B(n_618),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_850),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_801),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_SL g904 ( 
.A(n_796),
.B(n_707),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_854),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_843),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_843),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_796),
.B(n_769),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_801),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_803),
.B(n_618),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_812),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_813),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_808),
.B(n_769),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_851),
.B(n_623),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_845),
.B(n_623),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_808),
.B(n_750),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_843),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_843),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_843),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_849),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_846),
.B(n_781),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_803),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_845),
.A2(n_787),
.B1(n_785),
.B2(n_752),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_801),
.Y(n_924)
);

INVx8_ASAP7_75t_L g925 ( 
.A(n_885),
.Y(n_925)
);

INVxp67_ASAP7_75t_SL g926 ( 
.A(n_917),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_897),
.B(n_816),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_897),
.B(n_816),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_911),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_900),
.B(n_751),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_864),
.B(n_810),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_864),
.B(n_760),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_894),
.Y(n_933)
);

INVxp33_ASAP7_75t_L g934 ( 
.A(n_893),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_898),
.B(n_816),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_899),
.B(n_837),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_SL g937 ( 
.A(n_890),
.B(n_760),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_864),
.B(n_810),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_898),
.B(n_810),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_908),
.B(n_837),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_899),
.B(n_819),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_859),
.B(n_819),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_877),
.B(n_804),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_860),
.B(n_819),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_886),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_894),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_916),
.B(n_759),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_915),
.B(n_797),
.Y(n_948)
);

NOR2xp67_ASAP7_75t_L g949 ( 
.A(n_923),
.B(n_790),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_889),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_877),
.B(n_856),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_855),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_862),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_892),
.A2(n_625),
.B(n_595),
.C(n_794),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_915),
.B(n_797),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_914),
.B(n_761),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_891),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_892),
.B(n_521),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_880),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_856),
.B(n_804),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_856),
.B(n_826),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_872),
.B(n_521),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_880),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_880),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_856),
.B(n_826),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_896),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_856),
.B(n_826),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_901),
.B(n_578),
.Y(n_968)
);

AND2x6_ASAP7_75t_SL g969 ( 
.A(n_913),
.B(n_683),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_902),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_904),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_905),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_862),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_921),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_914),
.B(n_762),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_L g976 ( 
.A(n_882),
.B(n_656),
.C(n_616),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_921),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_895),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_857),
.B(n_580),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_869),
.Y(n_980)
);

XOR2xp5_ASAP7_75t_L g981 ( 
.A(n_888),
.B(n_875),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_917),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_921),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_881),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_922),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_858),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_904),
.B(n_770),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_876),
.B(n_866),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_922),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_872),
.B(n_523),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_867),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_872),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_879),
.B(n_523),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_912),
.B(n_724),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_885),
.A2(n_666),
.B1(n_586),
.B2(n_590),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_868),
.B(n_774),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_861),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_870),
.B(n_524),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_871),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_873),
.B(n_524),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_865),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_874),
.B(n_823),
.Y(n_1002)
);

BUFx5_ASAP7_75t_L g1003 ( 
.A(n_910),
.Y(n_1003)
);

BUFx8_ASAP7_75t_L g1004 ( 
.A(n_901),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_869),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_901),
.B(n_602),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_874),
.B(n_823),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_906),
.B(n_774),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_907),
.B(n_528),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_918),
.B(n_531),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_919),
.B(n_727),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_878),
.B(n_852),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_869),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_878),
.B(n_852),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_920),
.B(n_531),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_883),
.B(n_728),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_883),
.B(n_699),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_884),
.B(n_887),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_884),
.B(n_852),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_887),
.B(n_852),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_863),
.B(n_699),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_901),
.B(n_805),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_901),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_869),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_903),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_903),
.B(n_700),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_903),
.B(n_700),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_924),
.B(n_805),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_903),
.B(n_702),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_910),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_863),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_924),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_909),
.B(n_730),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_909),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_910),
.B(n_702),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_L g1036 ( 
.A(n_910),
.B(n_585),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_910),
.B(n_732),
.C(n_731),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_SL g1038 ( 
.A(n_894),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_900),
.B(n_547),
.Y(n_1039)
);

AO22x2_ASAP7_75t_L g1040 ( 
.A1(n_981),
.A2(n_976),
.B1(n_942),
.B2(n_931),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_959),
.B(n_805),
.Y(n_1041)
);

OAI221xp5_ASAP7_75t_L g1042 ( 
.A1(n_930),
.A2(n_705),
.B1(n_846),
.B2(n_550),
.C(n_560),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_SL g1043 ( 
.A(n_979),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_978),
.Y(n_1044)
);

AO22x2_ASAP7_75t_L g1045 ( 
.A1(n_938),
.A2(n_579),
.B1(n_635),
.B2(n_622),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_929),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1016),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_951),
.A2(n_637),
.B1(n_625),
.B2(n_595),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

AO22x2_ASAP7_75t_L g1050 ( 
.A1(n_958),
.A2(n_635),
.B1(n_641),
.B2(n_622),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_945),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_950),
.Y(n_1052)
);

AO22x2_ASAP7_75t_L g1053 ( 
.A1(n_939),
.A2(n_641),
.B1(n_680),
.B2(n_637),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_1038),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_971),
.A2(n_680),
.B1(n_549),
.B2(n_553),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_957),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_947),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_966),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_994),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_970),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_959),
.B(n_805),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_972),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_SL g1063 ( 
.A(n_933),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_988),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_988),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1033),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1011),
.Y(n_1067)
);

NAND2x1_ASAP7_75t_L g1068 ( 
.A(n_980),
.B(n_805),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_974),
.B(n_593),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_986),
.Y(n_1070)
);

OAI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_992),
.A2(n_555),
.B1(n_567),
.B2(n_541),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_997),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_953),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_733),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_973),
.Y(n_1075)
);

AO22x2_ASAP7_75t_L g1076 ( 
.A1(n_1023),
.A2(n_577),
.B1(n_584),
.B2(n_570),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_991),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_933),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_985),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1039),
.B(n_603),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_964),
.B(n_822),
.Y(n_1081)
);

AO22x2_ASAP7_75t_L g1082 ( 
.A1(n_956),
.A2(n_614),
.B1(n_644),
.B2(n_604),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_964),
.B(n_822),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_926),
.B(n_657),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_975),
.A2(n_562),
.B1(n_564),
.B2(n_557),
.C(n_556),
.Y(n_1085)
);

AO22x2_ASAP7_75t_L g1086 ( 
.A1(n_962),
.A2(n_659),
.B1(n_662),
.B2(n_658),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_989),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_982),
.B(n_670),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_999),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_963),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_974),
.Y(n_1091)
);

AO22x2_ASAP7_75t_L g1092 ( 
.A1(n_990),
.A2(n_1006),
.B1(n_928),
.B2(n_927),
.Y(n_1092)
);

AO22x2_ASAP7_75t_L g1093 ( 
.A1(n_1006),
.A2(n_688),
.B1(n_692),
.B2(n_672),
.Y(n_1093)
);

OAI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_936),
.A2(n_569),
.B1(n_575),
.B2(n_568),
.C(n_566),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1001),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_984),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1034),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_940),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_964),
.B(n_828),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1002),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1002),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1007),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1034),
.Y(n_1103)
);

AO22x2_ASAP7_75t_L g1104 ( 
.A1(n_987),
.A2(n_696),
.B1(n_737),
.B2(n_734),
.Y(n_1104)
);

XNOR2xp5_ASAP7_75t_SL g1105 ( 
.A(n_934),
.B(n_1),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_977),
.B(n_601),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1007),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_977),
.B(n_940),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_977),
.B(n_607),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_933),
.B(n_828),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_946),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_943),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1018),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1032),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_941),
.A2(n_611),
.B1(n_615),
.B2(n_610),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1018),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_935),
.B(n_829),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_935),
.B(n_829),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_954),
.B(n_802),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_925),
.Y(n_1120)
);

AO22x2_ASAP7_75t_L g1121 ( 
.A1(n_1009),
.A2(n_786),
.B1(n_789),
.B2(n_784),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1031),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1012),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_996),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1015),
.B(n_802),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_925),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1012),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1014),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1014),
.Y(n_1129)
);

AO22x2_ASAP7_75t_L g1130 ( 
.A1(n_1010),
.A2(n_792),
.B1(n_793),
.B2(n_791),
.Y(n_1130)
);

OR2x6_ASAP7_75t_SL g1131 ( 
.A(n_1004),
.B(n_583),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_937),
.A2(n_621),
.B1(n_626),
.B2(n_620),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_946),
.B(n_980),
.Y(n_1133)
);

AO22x2_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_795),
.B1(n_10),
.B2(n_18),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1019),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_1038),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1019),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1005),
.B(n_814),
.Y(n_1138)
);

NAND2xp33_ASAP7_75t_L g1139 ( 
.A(n_1003),
.B(n_628),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1020),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1030),
.B(n_274),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1008),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1013),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_949),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_948),
.B(n_814),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_944),
.A2(n_647),
.B1(n_648),
.B2(n_631),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1024),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1025),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1028),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_961),
.Y(n_1151)
);

AO22x2_ASAP7_75t_L g1152 ( 
.A1(n_1026),
.A2(n_11),
.B1(n_19),
.B2(n_2),
.Y(n_1152)
);

AO22x2_ASAP7_75t_L g1153 ( 
.A1(n_1027),
.A2(n_11),
.B1(n_19),
.B2(n_2),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_961),
.A2(n_674),
.B1(n_675),
.B2(n_663),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_965),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_955),
.A2(n_678),
.B1(n_685),
.B2(n_677),
.Y(n_1156)
);

AO22x2_ASAP7_75t_L g1157 ( 
.A1(n_1029),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_998),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_965),
.A2(n_687),
.B1(n_694),
.B2(n_686),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_960),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_960),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_995),
.B(n_275),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_1021),
.B(n_1022),
.Y(n_1163)
);

AO22x2_ASAP7_75t_L g1164 ( 
.A1(n_1000),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_R g1165 ( 
.A(n_968),
.B(n_1004),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_967),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_SL g1167 ( 
.A1(n_969),
.A2(n_591),
.B1(n_594),
.B2(n_588),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_993),
.B(n_596),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1037),
.Y(n_1169)
);

AO22x2_ASAP7_75t_L g1170 ( 
.A1(n_1035),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_SL g1171 ( 
.A(n_1036),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1003),
.A2(n_605),
.B1(n_609),
.B2(n_597),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1003),
.Y(n_1173)
);

AND2x2_ASAP7_75t_SL g1174 ( 
.A(n_929),
.B(n_814),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_974),
.B(n_612),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1039),
.A2(n_820),
.B1(n_617),
.B2(n_624),
.Y(n_1176)
);

OAI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_930),
.A2(n_632),
.B1(n_634),
.B2(n_627),
.C(n_613),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_978),
.Y(n_1178)
);

CKINVDCx16_ASAP7_75t_R g1179 ( 
.A(n_940),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1039),
.A2(n_820),
.B1(n_638),
.B2(n_639),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_932),
.B(n_636),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_983),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_983),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_959),
.B(n_820),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_974),
.B(n_640),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_983),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_929),
.Y(n_1187)
);

AO22x2_ASAP7_75t_L g1188 ( 
.A1(n_981),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_930),
.A2(n_645),
.B1(n_651),
.B2(n_643),
.C(n_642),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_959),
.B(n_276),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_929),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_930),
.B(n_653),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1039),
.A2(n_655),
.B(n_660),
.C(n_654),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_983),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_978),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_983),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_983),
.Y(n_1197)
);

AO22x2_ASAP7_75t_L g1198 ( 
.A1(n_981),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_983),
.Y(n_1199)
);

AO22x2_ASAP7_75t_L g1200 ( 
.A1(n_981),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_929),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1174),
.B(n_661),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1064),
.A2(n_667),
.B1(n_668),
.B2(n_665),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1065),
.B(n_673),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1192),
.A2(n_689),
.B1(n_690),
.B2(n_679),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1059),
.B(n_691),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_1139),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1116),
.B(n_697),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1113),
.A2(n_279),
.B(n_278),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1046),
.B(n_280),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1098),
.B(n_282),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1063),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1051),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1163),
.A2(n_284),
.B(n_283),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1090),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_L g1216 ( 
.A(n_1080),
.B(n_286),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1166),
.A2(n_288),
.B(n_287),
.Y(n_1217)
);

INVx5_ASAP7_75t_L g1218 ( 
.A(n_1074),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1182),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1124),
.B(n_15),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1100),
.B(n_16),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1183),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1078),
.B(n_289),
.Y(n_1223)
);

NOR3xp33_ASAP7_75t_L g1224 ( 
.A(n_1177),
.B(n_17),
.C(n_18),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1151),
.A2(n_291),
.B1(n_293),
.B2(n_290),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1101),
.B(n_17),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1085),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1179),
.B(n_1057),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1187),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1054),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1173),
.A2(n_297),
.B(n_296),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1191),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1155),
.A2(n_302),
.B(n_300),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1201),
.Y(n_1234)
);

AO32x1_ASAP7_75t_L g1235 ( 
.A1(n_1048),
.A2(n_23),
.A3(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1102),
.B(n_1107),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1173),
.A2(n_306),
.B(n_305),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1123),
.B(n_25),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1127),
.B(n_25),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1047),
.B(n_26),
.Y(n_1240)
);

AO32x2_ASAP7_75t_L g1241 ( 
.A1(n_1092),
.A2(n_1050),
.A3(n_1172),
.B1(n_1055),
.B2(n_1154),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1128),
.B(n_26),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1108),
.A2(n_308),
.B1(n_310),
.B2(n_307),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1142),
.B(n_1066),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1052),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1173),
.A2(n_313),
.B(n_311),
.Y(n_1246)
);

BUFx12f_ASAP7_75t_L g1247 ( 
.A(n_1136),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1181),
.B(n_27),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1067),
.B(n_28),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1168),
.B(n_28),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1056),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1160),
.A2(n_315),
.B1(n_316),
.B2(n_314),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1111),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1129),
.B(n_29),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1145),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1042),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1161),
.A2(n_320),
.B1(n_321),
.B2(n_319),
.Y(n_1257)
);

AO21x1_ASAP7_75t_L g1258 ( 
.A1(n_1119),
.A2(n_32),
.B(n_33),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1189),
.B(n_33),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1120),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1040),
.A2(n_325),
.B1(n_327),
.B2(n_324),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1112),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1186),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1158),
.B(n_40),
.Y(n_1264)
);

AOI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1094),
.A2(n_40),
.B(n_41),
.Y(n_1265)
);

AO22x1_ASAP7_75t_L g1266 ( 
.A1(n_1136),
.A2(n_1091),
.B1(n_1141),
.B2(n_1060),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1096),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1135),
.B(n_42),
.Y(n_1268)
);

AOI33xp33_ASAP7_75t_L g1269 ( 
.A1(n_1058),
.A2(n_45),
.A3(n_47),
.B1(n_43),
.B2(n_44),
.B3(n_46),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1137),
.B(n_43),
.Y(n_1270)
);

NOR3xp33_ASAP7_75t_L g1271 ( 
.A(n_1175),
.B(n_45),
.C(n_47),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1062),
.B(n_333),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1140),
.B(n_48),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_335),
.B(n_334),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1126),
.B(n_338),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1150),
.A2(n_342),
.B(n_341),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1194),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1086),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_L g1279 ( 
.A1(n_1125),
.A2(n_345),
.B(n_346),
.C(n_343),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1040),
.A2(n_350),
.B1(n_352),
.B2(n_348),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1193),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1156),
.B(n_52),
.C(n_53),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1043),
.B(n_52),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1196),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1069),
.A2(n_1109),
.B(n_1106),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1197),
.B(n_54),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1185),
.A2(n_364),
.B(n_356),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1044),
.A2(n_366),
.B(n_365),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1199),
.B(n_1070),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1074),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_L g1291 ( 
.A(n_1141),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1171),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1072),
.B(n_367),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1071),
.A2(n_55),
.B(n_56),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1077),
.B(n_55),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1133),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_L g1297 ( 
.A1(n_1084),
.A2(n_369),
.B(n_370),
.C(n_368),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1105),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1298)
);

BUFx4_ASAP7_75t_SL g1299 ( 
.A(n_1146),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1089),
.B(n_58),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1088),
.B(n_59),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1095),
.B(n_59),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1180),
.B(n_371),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1146),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_1304)
);

OR2x6_ASAP7_75t_SL g1305 ( 
.A(n_1169),
.B(n_60),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1121),
.B(n_60),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1104),
.B(n_61),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1068),
.A2(n_376),
.B(n_375),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1147),
.B(n_61),
.Y(n_1309)
);

NAND3x1_ASAP7_75t_L g1310 ( 
.A(n_1188),
.B(n_62),
.C(n_63),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_SL g1311 ( 
.A1(n_1114),
.A2(n_378),
.B(n_379),
.C(n_377),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1121),
.B(n_64),
.Y(n_1312)
);

BUFx8_ASAP7_75t_SL g1313 ( 
.A(n_1178),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1130),
.B(n_65),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1115),
.B(n_65),
.Y(n_1315)
);

OA22x2_ASAP7_75t_L g1316 ( 
.A1(n_1188),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1073),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1075),
.A2(n_381),
.B(n_380),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1167),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1045),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1068),
.A2(n_388),
.B(n_385),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1162),
.B(n_389),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1184),
.A2(n_396),
.B(n_393),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1097),
.A2(n_404),
.B1(n_405),
.B2(n_401),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1041),
.A2(n_1061),
.B(n_1103),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1049),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1195),
.A2(n_410),
.B(n_408),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1122),
.A2(n_412),
.B1(n_414),
.B2(n_411),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1079),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1190),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1081),
.A2(n_416),
.B(n_415),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1083),
.A2(n_418),
.B(n_417),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1110),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1176),
.B(n_66),
.C(n_67),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1130),
.B(n_69),
.Y(n_1335)
);

AOI21xp33_ASAP7_75t_L g1336 ( 
.A1(n_1082),
.A2(n_70),
.B(n_71),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1099),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1159),
.B(n_419),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1087),
.A2(n_422),
.B(n_421),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_R g1340 ( 
.A(n_1148),
.B(n_423),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1143),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1053),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1149),
.A2(n_426),
.B(n_425),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1132),
.B(n_72),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1138),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1050),
.B(n_72),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1076),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1131),
.B(n_73),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1053),
.Y(n_1349)
);

AO22x1_ASAP7_75t_L g1350 ( 
.A1(n_1198),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1093),
.A2(n_430),
.B(n_427),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1076),
.A2(n_432),
.B(n_431),
.Y(n_1352)
);

BUFx8_ASAP7_75t_L g1353 ( 
.A(n_1198),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1165),
.B(n_1086),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1055),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1082),
.A2(n_434),
.B(n_433),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1104),
.B(n_75),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1200),
.B(n_77),
.Y(n_1358)
);

AOI21xp33_ASAP7_75t_L g1359 ( 
.A1(n_1134),
.A2(n_77),
.B(n_78),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1200),
.B(n_78),
.Y(n_1360)
);

OAI21xp33_ASAP7_75t_L g1361 ( 
.A1(n_1134),
.A2(n_79),
.B(n_80),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1170),
.A2(n_437),
.B(n_436),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1164),
.B(n_80),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1152),
.A2(n_440),
.B1(n_441),
.B2(n_439),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1153),
.A2(n_443),
.B(n_442),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1164),
.B(n_81),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1153),
.Y(n_1367)
);

CKINVDCx10_ASAP7_75t_R g1368 ( 
.A(n_1157),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_SL g1369 ( 
.A(n_1157),
.B(n_444),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1064),
.A2(n_448),
.B1(n_450),
.B2(n_447),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1215),
.B(n_81),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1260),
.Y(n_1372)
);

AND3x1_ASAP7_75t_SL g1373 ( 
.A(n_1353),
.B(n_1368),
.C(n_1310),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1236),
.B(n_82),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1298),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1213),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1245),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1251),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1229),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1277),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1247),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1367),
.B(n_1221),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1226),
.B(n_84),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1215),
.B(n_85),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1212),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1250),
.B(n_86),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1292),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1289),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1291),
.B(n_86),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1264),
.B(n_87),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1291),
.B(n_88),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1248),
.B(n_88),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1219),
.B(n_89),
.Y(n_1393)
);

AND3x1_ASAP7_75t_SL g1394 ( 
.A(n_1353),
.B(n_89),
.C(n_90),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1222),
.B(n_91),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1309),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1315),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1358),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1204),
.B(n_96),
.Y(n_1399)
);

AND3x1_ASAP7_75t_SL g1400 ( 
.A(n_1368),
.B(n_97),
.C(n_98),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1208),
.B(n_99),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1284),
.B(n_100),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1238),
.B(n_100),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1317),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1249),
.B(n_101),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1326),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1333),
.B(n_452),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1239),
.B(n_101),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1215),
.B(n_506),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1329),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1242),
.B(n_1254),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1360),
.B(n_104),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1268),
.B(n_104),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1355),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1296),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1266),
.B(n_453),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1292),
.Y(n_1417)
);

AOI22x1_ASAP7_75t_L g1418 ( 
.A1(n_1285),
.A2(n_455),
.B1(n_456),
.B2(n_454),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1313),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1341),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1270),
.B(n_105),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1234),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1296),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1296),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1273),
.B(n_106),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1267),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1218),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1286),
.Y(n_1428)
);

AND3x1_ASAP7_75t_SL g1429 ( 
.A(n_1350),
.B(n_107),
.C(n_108),
.Y(n_1429)
);

AND3x1_ASAP7_75t_SL g1430 ( 
.A(n_1305),
.B(n_108),
.C(n_109),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1349),
.B(n_110),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1316),
.A2(n_113),
.B1(n_110),
.B2(n_111),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1302),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1228),
.B(n_111),
.Y(n_1434)
);

AND3x1_ASAP7_75t_SL g1435 ( 
.A(n_1369),
.B(n_114),
.C(n_115),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1295),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1307),
.B(n_114),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1203),
.B(n_115),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1244),
.B(n_116),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1347),
.B(n_117),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1203),
.B(n_118),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1232),
.B(n_118),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1253),
.B(n_119),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1342),
.B(n_120),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1337),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1223),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1223),
.Y(n_1447)
);

AND3x1_ASAP7_75t_SL g1448 ( 
.A(n_1359),
.B(n_120),
.C(n_121),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1300),
.Y(n_1449)
);

AND3x1_ASAP7_75t_SL g1450 ( 
.A(n_1361),
.B(n_121),
.C(n_122),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1301),
.B(n_123),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1320),
.B(n_1207),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1230),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1346),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1344),
.B(n_123),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1319),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1259),
.B(n_124),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1220),
.B(n_124),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1345),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1218),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1211),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1240),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1210),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1269),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1330),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1306),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_SL g1467 ( 
.A(n_1205),
.B(n_128),
.C(n_129),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1330),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1218),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1206),
.B(n_130),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1255),
.B(n_131),
.Y(n_1471)
);

OR2x6_ASAP7_75t_SL g1472 ( 
.A(n_1334),
.B(n_132),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1312),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1314),
.Y(n_1474)
);

NAND2xp33_ASAP7_75t_L g1475 ( 
.A(n_1224),
.B(n_457),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1357),
.B(n_132),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1335),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1290),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1214),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_L g1480 ( 
.A(n_1340),
.B(n_459),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1202),
.B(n_133),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1338),
.B(n_133),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1258),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1363),
.Y(n_1484)
);

AND3x1_ASAP7_75t_SL g1485 ( 
.A(n_1348),
.B(n_134),
.C(n_135),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1275),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1303),
.B(n_134),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1299),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1365),
.B(n_135),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1283),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1354),
.B(n_136),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1366),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1241),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1362),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1263),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1272),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1271),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1262),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1325),
.B(n_137),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1278),
.B(n_138),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1293),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1322),
.B(n_139),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1261),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1282),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1280),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1336),
.B(n_139),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1352),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1265),
.B(n_140),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1227),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1331),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1364),
.B(n_141),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1332),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1294),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1281),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1256),
.B(n_142),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1243),
.Y(n_1516)
);

A2O1A1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1233),
.A2(n_143),
.B(n_144),
.C(n_145),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1276),
.B(n_143),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1279),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1311),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1304),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1356),
.B(n_144),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1288),
.B(n_147),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1297),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1328),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1231),
.B(n_505),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1225),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1318),
.B(n_147),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1351),
.B(n_148),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1388),
.B(n_1287),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1416),
.B(n_1237),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1385),
.B(n_1370),
.Y(n_1532)
);

NAND2xp33_ASAP7_75t_L g1533 ( 
.A(n_1503),
.B(n_1327),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1376),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1411),
.B(n_1428),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1505),
.A2(n_1216),
.B1(n_1252),
.B2(n_1257),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1372),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1446),
.B(n_1246),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1465),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1510),
.A2(n_1209),
.B(n_1217),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1379),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1377),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1512),
.A2(n_1274),
.B(n_1343),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1512),
.A2(n_1339),
.B(n_1323),
.Y(n_1544)
);

NAND2x1_ASAP7_75t_L g1545 ( 
.A(n_1520),
.B(n_1308),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1524),
.A2(n_1519),
.B(n_1452),
.Y(n_1546)
);

AOI221x1_ASAP7_75t_L g1547 ( 
.A1(n_1511),
.A2(n_1324),
.B1(n_1321),
.B2(n_1235),
.C(n_151),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1378),
.Y(n_1548)
);

AOI21xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1455),
.A2(n_148),
.B(n_149),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1436),
.B(n_150),
.Y(n_1550)
);

BUFx2_ASAP7_75t_SL g1551 ( 
.A(n_1453),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1416),
.B(n_1235),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1415),
.Y(n_1553)
);

BUFx2_ASAP7_75t_SL g1554 ( 
.A(n_1422),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1449),
.B(n_151),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1478),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1456),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1415),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1494),
.A2(n_1235),
.B(n_154),
.C(n_156),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1504),
.A2(n_152),
.B(n_156),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1484),
.B(n_157),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1452),
.A2(n_504),
.B(n_461),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1492),
.B(n_158),
.Y(n_1563)
);

INVx8_ASAP7_75t_L g1564 ( 
.A(n_1427),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1380),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1404),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1462),
.B(n_1454),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_SL g1568 ( 
.A1(n_1483),
.A2(n_159),
.B(n_160),
.C(n_161),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1516),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1415),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1460),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1475),
.B(n_163),
.C(n_164),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1465),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1466),
.B(n_163),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1490),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1457),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.C(n_168),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1423),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1473),
.B(n_1474),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1437),
.B(n_166),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1491),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1457),
.A2(n_169),
.B(n_170),
.C(n_171),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1375),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1477),
.B(n_172),
.Y(n_1583)
);

AO22x1_ASAP7_75t_L g1584 ( 
.A1(n_1432),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1507),
.A2(n_462),
.B(n_460),
.Y(n_1585)
);

AO22x2_ASAP7_75t_L g1586 ( 
.A1(n_1432),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1426),
.Y(n_1587)
);

O2A1O1Ixp5_ASAP7_75t_L g1588 ( 
.A1(n_1515),
.A2(n_178),
.B(n_179),
.C(n_180),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1481),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1416),
.B(n_463),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1423),
.Y(n_1591)
);

OAI21xp33_ASAP7_75t_L g1592 ( 
.A1(n_1489),
.A2(n_181),
.B(n_182),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1467),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1451),
.B(n_183),
.Y(n_1594)
);

BUFx5_ASAP7_75t_L g1595 ( 
.A(n_1526),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1518),
.A2(n_184),
.B(n_185),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1516),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_1597)
);

INVx4_ASAP7_75t_L g1598 ( 
.A(n_1465),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1433),
.B(n_188),
.Y(n_1599)
);

AOI222xp33_ASAP7_75t_L g1600 ( 
.A1(n_1398),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.C1(n_191),
.C2(n_193),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1406),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1410),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1447),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_1603)
);

AOI21xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1397),
.A2(n_194),
.B(n_195),
.Y(n_1604)
);

O2A1O1Ixp5_ASAP7_75t_SL g1605 ( 
.A1(n_1513),
.A2(n_194),
.B(n_195),
.C(n_196),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1464),
.B(n_196),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1387),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1424),
.B(n_1468),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1469),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_L g1610 ( 
.A(n_1417),
.Y(n_1610)
);

INVx4_ASAP7_75t_L g1611 ( 
.A(n_1424),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1486),
.B(n_464),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1420),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1374),
.B(n_197),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1419),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1399),
.B(n_465),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1480),
.A2(n_503),
.B(n_498),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1374),
.B(n_197),
.Y(n_1618)
);

AOI21xp33_ASAP7_75t_L g1619 ( 
.A1(n_1514),
.A2(n_199),
.B(n_200),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1382),
.B(n_200),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1382),
.B(n_201),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1393),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1518),
.A2(n_201),
.B(n_202),
.C(n_203),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1389),
.B(n_1391),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1393),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_SL g1626 ( 
.A1(n_1517),
.A2(n_204),
.B(n_205),
.C(n_207),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1521),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1401),
.B(n_208),
.Y(n_1628)
);

AND2x4_ASAP7_75t_SL g1629 ( 
.A(n_1409),
.B(n_466),
.Y(n_1629)
);

AOI221x1_ASAP7_75t_L g1630 ( 
.A1(n_1489),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.C(n_212),
.Y(n_1630)
);

NAND2x1p5_ASAP7_75t_L g1631 ( 
.A(n_1488),
.B(n_467),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1451),
.B(n_209),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1389),
.B(n_210),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1391),
.B(n_469),
.Y(n_1634)
);

BUFx8_ASAP7_75t_SL g1635 ( 
.A(n_1381),
.Y(n_1635)
);

INVx3_ASAP7_75t_SL g1636 ( 
.A(n_1488),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1412),
.B(n_212),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1500),
.B(n_213),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1445),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1409),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_L g1641 ( 
.A(n_1482),
.B(n_215),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1395),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1373),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1459),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1442),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1390),
.B(n_218),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1443),
.Y(n_1647)
);

NOR2x1p5_ASAP7_75t_L g1648 ( 
.A(n_1482),
.B(n_470),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1434),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1523),
.A2(n_218),
.B(n_219),
.C(n_220),
.Y(n_1650)
);

INVx5_ASAP7_75t_L g1651 ( 
.A(n_1526),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1527),
.A2(n_497),
.B(n_496),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1528),
.A2(n_220),
.B(n_221),
.C(n_222),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1407),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1499),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1529),
.A2(n_223),
.B(n_224),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1438),
.B(n_223),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1407),
.B(n_471),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1431),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1525),
.A2(n_1479),
.B(n_1496),
.Y(n_1660)
);

AOI222xp33_ASAP7_75t_L g1661 ( 
.A1(n_1441),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.C1(n_228),
.C2(n_229),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1470),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1553),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1533),
.A2(n_1536),
.B(n_1616),
.C(n_1656),
.Y(n_1664)
);

CKINVDCx16_ASAP7_75t_R g1665 ( 
.A(n_1551),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1651),
.B(n_1431),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1596),
.A2(n_1509),
.B(n_1396),
.C(n_1497),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1535),
.B(n_1506),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1613),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1582),
.A2(n_1651),
.B1(n_1593),
.B2(n_1472),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1649),
.B(n_1476),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1659),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1541),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1575),
.B(n_1371),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1580),
.A2(n_1461),
.B1(n_1463),
.B2(n_1444),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1572),
.A2(n_1487),
.B(n_1408),
.C(n_1383),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_SL g1677 ( 
.A(n_1635),
.B(n_1397),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1587),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1537),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1640),
.B(n_1522),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1655),
.B(n_1444),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1540),
.A2(n_1487),
.B(n_1498),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1662),
.B(n_1386),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1592),
.A2(n_1383),
.B(n_1403),
.C(n_1408),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1637),
.B(n_1405),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1622),
.B(n_1508),
.Y(n_1686)
);

A2O1A1Ixp33_ASAP7_75t_SL g1687 ( 
.A1(n_1560),
.A2(n_1439),
.B(n_1495),
.C(n_1414),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1641),
.A2(n_1414),
.B(n_1471),
.C(n_1458),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1640),
.B(n_1440),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1534),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1640),
.B(n_1440),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1579),
.B(n_1392),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1384),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1578),
.B(n_1403),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1543),
.A2(n_1501),
.B(n_1418),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1542),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1548),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1567),
.B(n_1594),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1625),
.B(n_1413),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1556),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1642),
.B(n_1421),
.Y(n_1701)
);

CKINVDCx6p67_ASAP7_75t_R g1702 ( 
.A(n_1636),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1554),
.Y(n_1703)
);

NOR2x2_ASAP7_75t_L g1704 ( 
.A(n_1590),
.B(n_1400),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1581),
.A2(n_1425),
.B(n_1502),
.C(n_1402),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1565),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1607),
.B(n_1435),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1598),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1590),
.A2(n_1658),
.B(n_1630),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1658),
.A2(n_1630),
.B(n_1617),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1601),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1634),
.A2(n_1450),
.B(n_1429),
.C(n_1485),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1602),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1544),
.A2(n_1493),
.B(n_1448),
.Y(n_1714)
);

CKINVDCx14_ASAP7_75t_R g1715 ( 
.A(n_1610),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1615),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1557),
.B(n_472),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1624),
.B(n_1430),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1614),
.B(n_225),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1600),
.A2(n_1394),
.B(n_229),
.C(n_230),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1643),
.Y(n_1721)
);

CKINVDCx20_ASAP7_75t_R g1722 ( 
.A(n_1645),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1618),
.B(n_226),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1566),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1650),
.A2(n_231),
.B(n_232),
.C(n_233),
.Y(n_1725)
);

OR2x4_ASAP7_75t_L g1726 ( 
.A(n_1553),
.B(n_232),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1608),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1564),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1620),
.B(n_234),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1621),
.B(n_236),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1577),
.B(n_494),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1632),
.B(n_236),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_SL g1733 ( 
.A1(n_1619),
.A2(n_237),
.B(n_238),
.C(n_239),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1553),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1646),
.B(n_492),
.Y(n_1735)
);

O2A1O1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1653),
.A2(n_237),
.B(n_239),
.C(n_240),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1638),
.B(n_491),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1546),
.A2(n_490),
.B(n_488),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1564),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1530),
.A2(n_487),
.B(n_486),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1604),
.A2(n_1628),
.B(n_1623),
.C(n_1576),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1561),
.B(n_241),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1647),
.B(n_1639),
.Y(n_1743)
);

INVx6_ASAP7_75t_L g1744 ( 
.A(n_1558),
.Y(n_1744)
);

OR2x2_ASAP7_75t_SL g1745 ( 
.A(n_1583),
.B(n_241),
.Y(n_1745)
);

OR2x6_ASAP7_75t_SL g1746 ( 
.A(n_1563),
.B(n_242),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1574),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1549),
.A2(n_242),
.B(n_243),
.C(n_244),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1591),
.B(n_484),
.Y(n_1749)
);

BUFx5_ASAP7_75t_L g1750 ( 
.A(n_1538),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1690),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1664),
.A2(n_1586),
.B1(n_1589),
.B2(n_1648),
.Y(n_1752)
);

BUFx4f_ASAP7_75t_SL g1753 ( 
.A(n_1702),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1696),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1720),
.A2(n_1661),
.B(n_1597),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1697),
.B(n_1552),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1677),
.A2(n_1532),
.B1(n_1547),
.B2(n_1552),
.Y(n_1757)
);

BUFx4f_ASAP7_75t_SL g1758 ( 
.A(n_1722),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1706),
.B(n_1711),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1668),
.B(n_1681),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1675),
.A2(n_1531),
.B1(n_1586),
.B2(n_1595),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1670),
.A2(n_1569),
.B1(n_1538),
.B2(n_1531),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1707),
.A2(n_1595),
.B1(n_1627),
.B2(n_1633),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1746),
.A2(n_1631),
.B1(n_1612),
.B2(n_1606),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1712),
.A2(n_1629),
.B(n_1603),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1713),
.B(n_1559),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1725),
.A2(n_1652),
.B(n_1562),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1665),
.B(n_1571),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1669),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1667),
.A2(n_1612),
.B1(n_1555),
.B2(n_1550),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1741),
.A2(n_1595),
.B1(n_1584),
.B2(n_1609),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1678),
.Y(n_1772)
);

BUFx4f_ASAP7_75t_SL g1773 ( 
.A(n_1716),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1724),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1709),
.A2(n_1599),
.B1(n_1644),
.B2(n_1611),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1739),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1734),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1721),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1694),
.B(n_1660),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1734),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1700),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_SL g1782 ( 
.A1(n_1718),
.A2(n_1585),
.B1(n_1626),
.B2(n_1568),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1698),
.B(n_1545),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1672),
.B(n_1605),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1715),
.Y(n_1785)
);

CKINVDCx11_ASAP7_75t_R g1786 ( 
.A(n_1703),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1666),
.A2(n_1680),
.B1(n_1674),
.B2(n_1693),
.Y(n_1787)
);

BUFx12f_ASAP7_75t_L g1788 ( 
.A(n_1728),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1673),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1710),
.A2(n_1573),
.B1(n_1539),
.B2(n_1570),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1684),
.A2(n_1570),
.B1(n_1558),
.B2(n_1588),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1680),
.A2(n_1570),
.B1(n_1558),
.B2(n_247),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1693),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1689),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1747),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1752),
.A2(n_1736),
.B1(n_1748),
.B2(n_1688),
.C(n_1687),
.Y(n_1796)
);

INVx3_ASAP7_75t_SL g1797 ( 
.A(n_1785),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1751),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1751),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1754),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1756),
.B(n_1743),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1755),
.A2(n_1689),
.B1(n_1691),
.B2(n_1717),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1789),
.B(n_1671),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1772),
.B(n_1686),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1781),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1754),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1756),
.B(n_1727),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_R g1808 ( 
.A(n_1785),
.B(n_1685),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_L g1809 ( 
.A(n_1770),
.B(n_1676),
.C(n_1705),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_L g1810 ( 
.A(n_1761),
.B(n_1730),
.C(n_1729),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1774),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1788),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1777),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1757),
.A2(n_1732),
.B1(n_1742),
.B2(n_1733),
.C(n_1701),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1767),
.A2(n_1682),
.B(n_1738),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1774),
.Y(n_1816)
);

NAND2xp33_ASAP7_75t_L g1817 ( 
.A(n_1771),
.B(n_1750),
.Y(n_1817)
);

INVxp33_ASAP7_75t_L g1818 ( 
.A(n_1768),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1775),
.B(n_1699),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1788),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1760),
.B(n_1719),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1765),
.A2(n_1740),
.B(n_1714),
.C(n_1695),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1759),
.B(n_1727),
.Y(n_1823)
);

INVx4_ASAP7_75t_L g1824 ( 
.A(n_1777),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1779),
.B(n_1750),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1780),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1764),
.B(n_1691),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1805),
.B(n_1769),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1799),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1825),
.B(n_1783),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1812),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1826),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1799),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1800),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1800),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1809),
.A2(n_1762),
.B1(n_1793),
.B2(n_1795),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1811),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1798),
.Y(n_1839)
);

CKINVDCx14_ASAP7_75t_R g1840 ( 
.A(n_1803),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1806),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1807),
.B(n_1823),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1801),
.B(n_1787),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1801),
.B(n_1784),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1801),
.B(n_1784),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1807),
.B(n_1766),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1807),
.B(n_1823),
.Y(n_1847)
);

OR2x6_ASAP7_75t_SL g1848 ( 
.A(n_1831),
.B(n_1778),
.Y(n_1848)
);

INVxp67_ASAP7_75t_SL g1849 ( 
.A(n_1830),
.Y(n_1849)
);

OAI21x1_ASAP7_75t_L g1850 ( 
.A1(n_1834),
.A2(n_1815),
.B(n_1816),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1833),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1846),
.B(n_1823),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1844),
.B(n_1819),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1838),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1838),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1838),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1852),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1853),
.B(n_1844),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1851),
.B(n_1845),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1850),
.B(n_1845),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1849),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1854),
.Y(n_1862)
);

OAI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1859),
.A2(n_1837),
.B1(n_1818),
.B2(n_1848),
.Y(n_1863)
);

INVx2_ASAP7_75t_SL g1864 ( 
.A(n_1861),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1858),
.B(n_1831),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1857),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1861),
.Y(n_1867)
);

AND2x4_ASAP7_75t_SL g1868 ( 
.A(n_1862),
.B(n_1832),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1860),
.Y(n_1869)
);

INVx4_ASAP7_75t_L g1870 ( 
.A(n_1861),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1859),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1868),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1867),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1864),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1871),
.B(n_1821),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1871),
.B(n_1846),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1870),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1870),
.Y(n_1878)
);

AOI32xp33_ASAP7_75t_L g1879 ( 
.A1(n_1863),
.A2(n_1817),
.A3(n_1818),
.B1(n_1796),
.B2(n_1819),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1866),
.B(n_1833),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1865),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1863),
.B(n_1849),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1877),
.B(n_1797),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1878),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1878),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1875),
.B(n_1869),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1873),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1872),
.B(n_1832),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1880),
.B(n_1881),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1876),
.Y(n_1890)
);

AOI21xp33_ASAP7_75t_L g1891 ( 
.A1(n_1889),
.A2(n_1882),
.B(n_1874),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1884),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_SL g1893 ( 
.A1(n_1885),
.A2(n_1882),
.B(n_1879),
.C(n_1794),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1890),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1891),
.B(n_1883),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1892),
.B(n_1888),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1894),
.B(n_1888),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1893),
.B(n_1886),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1897),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1895),
.B(n_1887),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1896),
.B(n_1887),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1898),
.A2(n_1837),
.B(n_1810),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1898),
.A2(n_1822),
.B(n_1814),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1899),
.Y(n_1904)
);

NAND2x1_ASAP7_75t_L g1905 ( 
.A(n_1901),
.B(n_1900),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1902),
.B(n_1797),
.Y(n_1906)
);

INVxp67_ASAP7_75t_L g1907 ( 
.A(n_1903),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1899),
.B(n_1778),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1899),
.B(n_1832),
.Y(n_1909)
);

INVxp67_ASAP7_75t_SL g1910 ( 
.A(n_1899),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1899),
.B(n_1832),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1899),
.Y(n_1912)
);

NOR2xp67_ASAP7_75t_SL g1913 ( 
.A(n_1899),
.B(n_1776),
.Y(n_1913)
);

AOI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1907),
.A2(n_1832),
.B1(n_1812),
.B2(n_1820),
.C(n_1679),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1910),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1832),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1906),
.A2(n_1776),
.B1(n_1758),
.B2(n_1840),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1913),
.A2(n_1820),
.B1(n_1753),
.B2(n_1786),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1904),
.B(n_1773),
.Y(n_1919)
);

OAI211xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1912),
.A2(n_1786),
.B(n_1723),
.C(n_1822),
.Y(n_1920)
);

AOI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1905),
.A2(n_1817),
.B1(n_1828),
.B2(n_1737),
.C(n_1692),
.Y(n_1921)
);

AOI221x1_ASAP7_75t_SL g1922 ( 
.A1(n_1909),
.A2(n_1726),
.B1(n_1855),
.B2(n_1854),
.C(n_1856),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1911),
.A2(n_1808),
.B(n_1828),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1906),
.A2(n_1745),
.B1(n_1802),
.B2(n_1856),
.Y(n_1924)
);

NOR3xp33_ASAP7_75t_L g1925 ( 
.A(n_1919),
.B(n_1735),
.C(n_1683),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1915),
.B(n_1847),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1914),
.B(n_1792),
.C(n_1731),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1917),
.B(n_1916),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1918),
.Y(n_1929)
);

OAI21xp33_ASAP7_75t_SL g1930 ( 
.A1(n_1923),
.A2(n_1855),
.B(n_1843),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1922),
.B(n_1839),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1924),
.Y(n_1932)
);

AND3x1_ASAP7_75t_L g1933 ( 
.A(n_1921),
.B(n_1708),
.C(n_1843),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1920),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1928),
.Y(n_1935)
);

AO22x2_ASAP7_75t_L g1936 ( 
.A1(n_1934),
.A2(n_1790),
.B1(n_1749),
.B2(n_1731),
.Y(n_1936)
);

AO22x2_ASAP7_75t_L g1937 ( 
.A1(n_1926),
.A2(n_1749),
.B1(n_1663),
.B2(n_1813),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1931),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1929),
.A2(n_1933),
.B1(n_1932),
.B2(n_1927),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1930),
.B(n_253),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1925),
.B(n_1663),
.C(n_1791),
.Y(n_1941)
);

A2O1A1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1940),
.A2(n_1827),
.B(n_254),
.C(n_255),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1939),
.B(n_1734),
.Y(n_1943)
);

AOI31xp33_ASAP7_75t_L g1944 ( 
.A1(n_1935),
.A2(n_1704),
.A3(n_1782),
.B(n_1763),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1937),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1938),
.B(n_1804),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_L g1947 ( 
.A(n_1941),
.B(n_253),
.C(n_254),
.Y(n_1947)
);

XOR2x2_ASAP7_75t_L g1948 ( 
.A(n_1936),
.B(n_256),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1948),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1942),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1946),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1945),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1947),
.Y(n_1953)
);

NAND5xp2_ASAP7_75t_L g1954 ( 
.A(n_1952),
.B(n_1943),
.C(n_1944),
.D(n_258),
.E(n_259),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1949),
.B(n_256),
.Y(n_1955)
);

AOI211xp5_ASAP7_75t_L g1956 ( 
.A1(n_1950),
.A2(n_257),
.B(n_258),
.C(n_259),
.Y(n_1956)
);

AOI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1953),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.C(n_263),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1955),
.A2(n_1951),
.B(n_261),
.Y(n_1958)
);

XNOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1956),
.B(n_260),
.Y(n_1959)
);

NAND4xp25_ASAP7_75t_L g1960 ( 
.A(n_1954),
.B(n_262),
.C(n_264),
.D(n_266),
.Y(n_1960)
);

XOR2xp5_ASAP7_75t_L g1961 ( 
.A(n_1957),
.B(n_264),
.Y(n_1961)
);

OAI222xp33_ASAP7_75t_L g1962 ( 
.A1(n_1955),
.A2(n_1813),
.B1(n_1824),
.B2(n_1839),
.C1(n_1835),
.C2(n_1836),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1961),
.A2(n_1744),
.B1(n_267),
.B2(n_268),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1960),
.A2(n_1829),
.B1(n_1744),
.B2(n_1842),
.Y(n_1964)
);

NAND4xp25_ASAP7_75t_L g1965 ( 
.A(n_1958),
.B(n_266),
.C(n_269),
.D(n_270),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1959),
.A2(n_1829),
.B1(n_1842),
.B2(n_1813),
.Y(n_1966)
);

INVxp67_ASAP7_75t_SL g1967 ( 
.A(n_1963),
.Y(n_1967)
);

AOI222xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1965),
.A2(n_1962),
.B1(n_1964),
.B2(n_1966),
.C1(n_269),
.C2(n_271),
.Y(n_1968)
);

NAND3xp33_ASAP7_75t_L g1969 ( 
.A(n_1965),
.B(n_271),
.C(n_272),
.Y(n_1969)
);

XNOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1969),
.B(n_1967),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1968),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1969),
.A2(n_272),
.B(n_473),
.Y(n_1972)
);

OAI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1970),
.A2(n_1847),
.B(n_1842),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1972),
.B(n_475),
.Y(n_1974)
);

OR2x6_ASAP7_75t_L g1975 ( 
.A(n_1974),
.B(n_1971),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1975),
.A2(n_1973),
.B(n_1842),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1976),
.A2(n_1827),
.B1(n_1824),
.B2(n_1841),
.Y(n_1977)
);

AOI211xp5_ASAP7_75t_L g1978 ( 
.A1(n_1977),
.A2(n_476),
.B(n_477),
.C(n_478),
.Y(n_1978)
);


endmodule