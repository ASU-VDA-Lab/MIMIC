module real_jpeg_4958_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_1),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_1),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_36),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_143),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_1),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_2),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_2),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_2),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_2),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_2),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_2),
.B(n_235),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_3),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_3),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_4),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_5),
.B(n_69),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_6),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_6),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_6),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_6),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_6),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_7),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_7),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_8),
.B(n_149),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_8),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_8),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_9),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_9),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_9),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_9),
.B(n_363),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_10),
.B(n_147),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_10),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_10),
.B(n_351),
.Y(n_350)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_12),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_12),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_12),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_13),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_13),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_13),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_13),
.B(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_13),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_14),
.Y(n_126)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_16),
.Y(n_320)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_17),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_324),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_272),
.B(n_323),
.Y(n_20)
);

AOI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_227),
.B(n_271),
.Y(n_21)
);

AO21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_152),
.B(n_226),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_136),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_24),
.B(n_136),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_74),
.B2(n_135),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_25),
.B(n_75),
.C(n_115),
.Y(n_270)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_49),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_27),
.B(n_50),
.C(n_73),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.C(n_45),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_28),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_141)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_31),
.Y(n_160)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_33),
.Y(n_149)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_38),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_39),
.B(n_45),
.Y(n_151)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_43),
.Y(n_268)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_44),
.Y(n_289)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_44),
.Y(n_365)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_47),
.B(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B1(n_72),
.B2(n_73),
.Y(n_49)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_55),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_55),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_55),
.B(n_232),
.C(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_57),
.B(n_63),
.C(n_68),
.Y(n_269)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_67),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_67),
.Y(n_349)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_70),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_71),
.Y(n_286)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_115),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_93),
.C(n_105),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_83),
.C(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_82),
.Y(n_258)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_82),
.Y(n_346)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_94),
.B1(n_105),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.C(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_219)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_98),
.B(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2x1_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_132),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_116),
.B(n_133),
.C(n_134),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_117),
.B(n_127),
.C(n_130),
.Y(n_243)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_126),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_129),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_150),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_137),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_140),
.B(n_150),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.C(n_144),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_141),
.B(n_142),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_148),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_221),
.B(n_225),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_206),
.B(n_220),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_190),
.B(n_205),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_181),
.B(n_189),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_168),
.C(n_173),
.Y(n_204)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_179),
.Y(n_194)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B(n_188),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_204),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_204),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_194),
.C(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_201),
.C(n_203),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_216),
.C(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_270),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_245),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_231),
.C(n_245),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_242),
.B2(n_244),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_290)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_248),
.C(n_262),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_249),
.B(n_255),
.C(n_259),
.Y(n_306)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.C(n_269),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_274),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_275),
.B(n_292),
.C(n_321),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_292),
.B1(n_321),
.B2(n_322),
.Y(n_276)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_291),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_327)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_284),
.B(n_287),
.C(n_290),
.Y(n_358)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_305),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_293),
.B(n_306),
.C(n_307),
.Y(n_356)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_293),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_298),
.CI(n_301),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_298),
.C(n_301),
.Y(n_368)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_318),
.B2(n_319),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_317),
.C(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_314),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_314),
.A2(n_317),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_371),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_370),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_370),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_354),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_339),
.B2(n_353),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_339),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_350),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_369),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_368),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_366),
.B2(n_367),
.Y(n_360)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_362),
.Y(n_367)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);


endmodule