module real_aes_7512_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g170 ( .A1(n_0), .A2(n_171), .B(n_174), .C(n_178), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_1), .B(n_162), .Y(n_181) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_3), .B(n_172), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_4), .A2(n_135), .B(n_138), .C(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_5), .A2(n_130), .B(n_544), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_6), .A2(n_100), .B1(n_111), .B2(n_749), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_7), .A2(n_130), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_8), .B(n_162), .Y(n_550) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_9), .A2(n_164), .B(n_236), .Y(n_235) );
AND2x6_ASAP7_75t_L g135 ( .A(n_10), .B(n_136), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_11), .A2(n_135), .B(n_138), .C(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g510 ( .A(n_12), .Y(n_510) );
INVx1_ASAP7_75t_L g103 ( .A(n_13), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_13), .B(n_40), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_14), .B(n_177), .Y(n_521) );
INVx1_ASAP7_75t_L g156 ( .A(n_15), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_16), .B(n_172), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_17), .A2(n_173), .B(n_530), .C(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_18), .B(n_162), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_19), .B(n_150), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_20), .A2(n_138), .B(n_141), .C(n_149), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_21), .A2(n_176), .B(n_244), .C(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_22), .B(n_177), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_23), .A2(n_75), .B1(n_453), .B2(n_741), .C1(n_744), .C2(n_745), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_24), .B(n_177), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_25), .Y(n_491) );
INVx1_ASAP7_75t_L g471 ( .A(n_26), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_27), .A2(n_138), .B(n_149), .C(n_239), .Y(n_238) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_28), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_29), .Y(n_517) );
INVx1_ASAP7_75t_L g485 ( .A(n_30), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_31), .A2(n_130), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g133 ( .A(n_32), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_33), .A2(n_188), .B(n_189), .C(n_193), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_34), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_35), .A2(n_176), .B(n_547), .C(n_549), .Y(n_546) );
INVxp67_ASAP7_75t_L g486 ( .A(n_36), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_37), .B(n_241), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_38), .A2(n_138), .B(n_149), .C(n_470), .Y(n_469) );
CKINVDCx14_ASAP7_75t_R g545 ( .A(n_39), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_40), .B(n_103), .Y(n_102) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_41), .A2(n_178), .B(n_508), .C(n_509), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_42), .B(n_129), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_43), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_44), .B(n_172), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_45), .B(n_130), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_46), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_47), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_48), .B(n_449), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_49), .A2(n_188), .B(n_193), .C(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g175 ( .A(n_50), .Y(n_175) );
INVx1_ASAP7_75t_L g219 ( .A(n_51), .Y(n_219) );
INVx1_ASAP7_75t_L g558 ( .A(n_52), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_53), .B(n_130), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_54), .Y(n_158) );
CKINVDCx14_ASAP7_75t_R g506 ( .A(n_55), .Y(n_506) );
INVx1_ASAP7_75t_L g136 ( .A(n_56), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_57), .B(n_130), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_58), .B(n_162), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_59), .A2(n_148), .B(n_204), .C(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
INVx1_ASAP7_75t_SL g548 ( .A(n_61), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_62), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_63), .B(n_172), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_64), .B(n_162), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_65), .B(n_173), .Y(n_254) );
INVx1_ASAP7_75t_L g494 ( .A(n_66), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g168 ( .A(n_67), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_68), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_69), .A2(n_138), .B(n_193), .C(n_202), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_70), .Y(n_228) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_72), .A2(n_130), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_73), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_74), .A2(n_130), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_75), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_76), .A2(n_129), .B(n_481), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_77), .Y(n_468) );
INVx1_ASAP7_75t_L g528 ( .A(n_78), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_79), .B(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_80), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_81), .A2(n_130), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g531 ( .A(n_82), .Y(n_531) );
INVx2_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx1_ASAP7_75t_L g520 ( .A(n_84), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_85), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_86), .B(n_177), .Y(n_255) );
INVx2_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
OR2x2_ASAP7_75t_L g444 ( .A(n_87), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g456 ( .A(n_87), .B(n_446), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_88), .A2(n_138), .B(n_193), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_89), .B(n_130), .Y(n_186) );
INVx1_ASAP7_75t_L g190 ( .A(n_90), .Y(n_190) );
INVxp67_ASAP7_75t_L g231 ( .A(n_91), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_92), .A2(n_118), .B1(n_440), .B2(n_441), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_92), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_93), .B(n_164), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_94), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g203 ( .A(n_95), .Y(n_203) );
INVx1_ASAP7_75t_L g250 ( .A(n_96), .Y(n_250) );
INVx2_ASAP7_75t_L g561 ( .A(n_97), .Y(n_561) );
AND2x2_ASAP7_75t_L g221 ( .A(n_98), .B(n_152), .Y(n_221) );
INVx2_ASAP7_75t_L g750 ( .A(n_100), .Y(n_750) );
AND2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_104), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_106), .B(n_107), .C(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g446 ( .A(n_106), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g460 ( .A(n_107), .B(n_446), .Y(n_460) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_107), .B(n_445), .Y(n_747) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_451), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g748 ( .A(n_113), .Y(n_748) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_442), .B(n_448), .Y(n_116) );
INVx1_ASAP7_75t_L g441 ( .A(n_118), .Y(n_441) );
INVx2_ASAP7_75t_L g457 ( .A(n_118), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_118), .A2(n_454), .B1(n_742), .B2(n_743), .Y(n_741) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_395), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_330), .Y(n_119) );
NAND4xp25_ASAP7_75t_SL g120 ( .A(n_121), .B(n_275), .C(n_299), .D(n_322), .Y(n_120) );
AOI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_212), .B1(n_246), .B2(n_259), .C(n_262), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_182), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_124), .A2(n_160), .B1(n_213), .B2(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_124), .B(n_183), .Y(n_333) );
AND2x2_ASAP7_75t_L g352 ( .A(n_124), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_124), .B(n_336), .Y(n_422) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
AND2x2_ASAP7_75t_L g290 ( .A(n_125), .B(n_183), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_125), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g313 ( .A(n_125), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g318 ( .A(n_125), .B(n_161), .Y(n_318) );
INVx2_ASAP7_75t_L g350 ( .A(n_125), .Y(n_350) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_125), .Y(n_394) );
AND2x2_ASAP7_75t_L g411 ( .A(n_125), .B(n_288), .Y(n_411) );
INVx5_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g329 ( .A(n_126), .B(n_288), .Y(n_329) );
AND2x4_ASAP7_75t_L g343 ( .A(n_126), .B(n_160), .Y(n_343) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_126), .Y(n_347) );
AND2x2_ASAP7_75t_L g367 ( .A(n_126), .B(n_282), .Y(n_367) );
AND2x2_ASAP7_75t_L g417 ( .A(n_126), .B(n_184), .Y(n_417) );
AND2x2_ASAP7_75t_L g427 ( .A(n_126), .B(n_161), .Y(n_427) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_157), .Y(n_126) );
AOI21xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_137), .B(n_150), .Y(n_127) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_131), .B(n_135), .Y(n_251) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g245 ( .A(n_133), .Y(n_245) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_134), .Y(n_144) );
INVx3_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g241 ( .A(n_134), .Y(n_241) );
BUFx3_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
INVx4_ASAP7_75t_SL g180 ( .A(n_135), .Y(n_180) );
INVx5_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx3_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_147), .Y(n_141) );
INVx2_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_146), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_146), .A2(n_192), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_146), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
O2A1O1Ixp5_ASAP7_75t_L g519 ( .A1(n_146), .A2(n_496), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_147), .A2(n_172), .B(n_471), .C(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_148), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_151), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_152), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_152), .A2(n_216), .B(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_152), .A2(n_251), .B(n_468), .C(n_469), .Y(n_467) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_152), .A2(n_504), .B(n_511), .Y(n_503) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g165 ( .A(n_153), .B(n_154), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_159), .A2(n_516), .B(n_522), .Y(n_515) );
AND2x2_ASAP7_75t_L g283 ( .A(n_160), .B(n_183), .Y(n_283) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_160), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_160), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g373 ( .A(n_160), .Y(n_373) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g261 ( .A(n_161), .B(n_198), .Y(n_261) );
AND2x2_ASAP7_75t_L g288 ( .A(n_161), .B(n_199), .Y(n_288) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_166), .B(n_181), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_163), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_200), .B(n_210), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_163), .B(n_211), .Y(n_210) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_163), .A2(n_249), .B(n_256), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_163), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_163), .A2(n_490), .B(n_497), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_163), .B(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_164), .A2(n_237), .B(n_238), .Y(n_236) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g258 ( .A(n_165), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_180), .Y(n_167) );
INVx2_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_169), .A2(n_180), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_169), .A2(n_180), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_169), .A2(n_180), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_169), .A2(n_180), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_169), .A2(n_180), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g557 ( .A1(n_169), .A2(n_180), .B(n_558), .C(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_172), .B(n_231), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_172), .A2(n_205), .B1(n_485), .B2(n_486), .Y(n_484) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_173), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_176), .B(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g508 ( .A(n_177), .Y(n_508) );
INVx2_ASAP7_75t_L g496 ( .A(n_178), .Y(n_496) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_179), .Y(n_192) );
INVx1_ASAP7_75t_L g532 ( .A(n_179), .Y(n_532) );
INVx1_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_182), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_196), .Y(n_182) );
OR2x2_ASAP7_75t_L g314 ( .A(n_183), .B(n_197), .Y(n_314) );
AND2x2_ASAP7_75t_L g351 ( .A(n_183), .B(n_261), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_183), .B(n_282), .Y(n_362) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_183), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_183), .B(n_318), .Y(n_435) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx2_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
AND2x2_ASAP7_75t_L g269 ( .A(n_184), .B(n_197), .Y(n_269) );
AND2x2_ASAP7_75t_L g385 ( .A(n_184), .B(n_280), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_184), .B(n_318), .Y(n_407) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_194), .Y(n_184) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_197), .Y(n_353) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_198), .Y(n_305) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx2_ASAP7_75t_L g282 ( .A(n_199), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_209), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_206), .C(n_207), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_205), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_205), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g549 ( .A(n_208), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_222), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_213), .B(n_295), .Y(n_414) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_214), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g266 ( .A(n_214), .B(n_267), .Y(n_266) );
INVx5_ASAP7_75t_SL g274 ( .A(n_214), .Y(n_274) );
OR2x2_ASAP7_75t_L g297 ( .A(n_214), .B(n_267), .Y(n_297) );
OR2x2_ASAP7_75t_L g307 ( .A(n_214), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g370 ( .A(n_214), .B(n_224), .Y(n_370) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_214), .B(n_223), .Y(n_408) );
NOR4xp25_ASAP7_75t_L g429 ( .A(n_214), .B(n_350), .C(n_430), .D(n_431), .Y(n_429) );
AND2x2_ASAP7_75t_L g439 ( .A(n_214), .B(n_271), .Y(n_439) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .Y(n_214) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g264 ( .A(n_223), .B(n_260), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_223), .B(n_266), .Y(n_433) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_233), .Y(n_223) );
OR2x2_ASAP7_75t_L g273 ( .A(n_224), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_224), .B(n_248), .Y(n_292) );
INVxp67_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_224), .B(n_267), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_224), .B(n_234), .Y(n_361) );
AND2x2_ASAP7_75t_L g376 ( .A(n_224), .B(n_271), .Y(n_376) );
OR2x2_ASAP7_75t_L g405 ( .A(n_224), .B(n_234), .Y(n_405) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_225), .A2(n_526), .B(n_533), .Y(n_525) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_225), .A2(n_543), .B(n_550), .Y(n_542) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_225), .A2(n_556), .B(n_562), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_233), .B(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_233), .B(n_274), .Y(n_413) );
OR2x2_ASAP7_75t_L g434 ( .A(n_233), .B(n_311), .Y(n_434) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g247 ( .A(n_234), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g271 ( .A(n_234), .B(n_267), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_234), .B(n_248), .Y(n_286) );
AND2x2_ASAP7_75t_L g356 ( .A(n_234), .B(n_280), .Y(n_356) );
AND2x2_ASAP7_75t_L g390 ( .A(n_234), .B(n_274), .Y(n_390) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_235), .B(n_274), .Y(n_293) );
AND2x2_ASAP7_75t_L g321 ( .A(n_235), .B(n_248), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_242), .B(n_243), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_243), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_246), .B(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_247), .A2(n_336), .B1(n_372), .B2(n_389), .C(n_391), .Y(n_388) );
INVx5_ASAP7_75t_SL g267 ( .A(n_248), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_252), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_251), .A2(n_491), .B(n_492), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_251), .A2(n_517), .B(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g479 ( .A(n_258), .Y(n_479) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OAI33xp33_ASAP7_75t_L g287 ( .A1(n_260), .A2(n_288), .A3(n_289), .B1(n_291), .B2(n_294), .B3(n_298), .Y(n_287) );
OR2x2_ASAP7_75t_L g303 ( .A(n_260), .B(n_304), .Y(n_303) );
AOI322xp5_ASAP7_75t_L g412 ( .A1(n_260), .A2(n_329), .A3(n_336), .B1(n_413), .B2(n_414), .C1(n_415), .C2(n_418), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_260), .B(n_288), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_SL g436 ( .A1(n_260), .A2(n_288), .B(n_437), .C(n_439), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_261), .A2(n_276), .B1(n_281), .B2(n_284), .C(n_287), .Y(n_275) );
INVx1_ASAP7_75t_L g368 ( .A(n_261), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_261), .B(n_417), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B1(n_268), .B2(n_270), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g345 ( .A(n_266), .B(n_280), .Y(n_345) );
AND2x2_ASAP7_75t_L g403 ( .A(n_266), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g311 ( .A(n_267), .B(n_274), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_267), .B(n_280), .Y(n_339) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_269), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_269), .B(n_347), .Y(n_401) );
OAI321xp33_ASAP7_75t_L g420 ( .A1(n_269), .A2(n_342), .A3(n_421), .B1(n_422), .B2(n_423), .C(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g387 ( .A(n_270), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_271), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g326 ( .A(n_271), .B(n_274), .Y(n_326) );
AOI321xp33_ASAP7_75t_L g384 ( .A1(n_271), .A2(n_288), .A3(n_385), .B1(n_386), .B2(n_387), .C(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g301 ( .A(n_273), .B(n_286), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_274), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_274), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_274), .B(n_360), .Y(n_397) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g320 ( .A(n_278), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g285 ( .A(n_279), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g393 ( .A(n_280), .Y(n_393) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_283), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_290), .B(n_325), .Y(n_374) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OR2x2_ASAP7_75t_L g338 ( .A(n_293), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g383 ( .A(n_293), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_294), .A2(n_341), .B1(n_344), .B2(n_346), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g438 ( .A(n_297), .B(n_361), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_302), .B1(n_306), .B2(n_312), .C(n_315), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g336 ( .A(n_305), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_SL g382 ( .A(n_308), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_310), .B(n_360), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_310), .A2(n_378), .B(n_380), .Y(n_377) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g423 ( .A(n_311), .B(n_405), .Y(n_423) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_SL g325 ( .A(n_314), .Y(n_325) );
AOI21xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_319), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g369 ( .A(n_321), .B(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g431 ( .A(n_321), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_325), .B(n_343), .Y(n_379) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g400 ( .A(n_329), .Y(n_400) );
NAND5xp2_ASAP7_75t_L g330 ( .A(n_331), .B(n_348), .C(n_357), .D(n_377), .E(n_384), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_337), .C(n_340), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_344), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
OAI21xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_352), .B(n_354), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_349), .A2(n_403), .B1(n_406), .B2(n_408), .C(n_409), .Y(n_402) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AOI321xp33_ASAP7_75t_L g357 ( .A1(n_350), .A2(n_358), .A3(n_362), .B1(n_363), .B2(n_369), .C(n_371), .Y(n_357) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g428 ( .A(n_362), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_364), .B(n_368), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g380 ( .A(n_365), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NOR2xp67_ASAP7_75t_SL g392 ( .A(n_366), .B(n_373), .Y(n_392) );
AOI321xp33_ASAP7_75t_SL g424 ( .A1(n_369), .A2(n_425), .A3(n_426), .B1(n_427), .B2(n_428), .C(n_429), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_374), .C(n_375), .Y(n_371) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_382), .B(n_390), .Y(n_419) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .C(n_394), .Y(n_391) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_420), .C(n_432), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_398), .B(n_402), .C(n_412), .Y(n_396) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_400), .B(n_401), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_401), .A2(n_433), .B1(n_434), .B2(n_435), .C(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g421 ( .A(n_403), .Y(n_421) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g425 ( .A(n_423), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_444), .Y(n_450) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_448), .A2(n_452), .B(n_748), .Y(n_451) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B1(n_458), .B2(n_461), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g743 ( .A(n_459), .Y(n_743) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g742 ( .A(n_461), .Y(n_742) );
OR4x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_631), .C(n_678), .D(n_718), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_577), .C(n_606), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_499), .B(n_534), .C(n_570), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_464), .A2(n_590), .B(n_607), .C(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_466), .B(n_569), .Y(n_568) );
INVx3_ASAP7_75t_SL g573 ( .A(n_466), .Y(n_573) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_466), .Y(n_585) );
AND2x4_ASAP7_75t_L g589 ( .A(n_466), .B(n_541), .Y(n_589) );
AND2x2_ASAP7_75t_L g600 ( .A(n_466), .B(n_489), .Y(n_600) );
OR2x2_ASAP7_75t_L g624 ( .A(n_466), .B(n_537), .Y(n_624) );
AND2x2_ASAP7_75t_L g637 ( .A(n_466), .B(n_542), .Y(n_637) );
AND2x2_ASAP7_75t_L g677 ( .A(n_466), .B(n_663), .Y(n_677) );
AND2x2_ASAP7_75t_L g684 ( .A(n_466), .B(n_647), .Y(n_684) );
AND2x2_ASAP7_75t_L g714 ( .A(n_466), .B(n_476), .Y(n_714) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_475), .B(n_641), .Y(n_653) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_488), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_476), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g591 ( .A(n_476), .B(n_488), .Y(n_591) );
BUFx3_ASAP7_75t_L g599 ( .A(n_476), .Y(n_599) );
OR2x2_ASAP7_75t_L g620 ( .A(n_476), .B(n_502), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_476), .B(n_641), .Y(n_731) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_480), .B(n_487), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_478), .A2(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g538 ( .A(n_480), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_487), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_488), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g584 ( .A(n_488), .Y(n_584) );
AND2x2_ASAP7_75t_L g647 ( .A(n_488), .B(n_542), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_488), .A2(n_650), .B1(n_652), .B2(n_654), .C(n_655), .Y(n_649) );
AND2x2_ASAP7_75t_L g663 ( .A(n_488), .B(n_537), .Y(n_663) );
AND2x2_ASAP7_75t_L g689 ( .A(n_488), .B(n_573), .Y(n_689) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g569 ( .A(n_489), .B(n_542), .Y(n_569) );
BUFx2_ASAP7_75t_L g703 ( .A(n_489), .Y(n_703) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI32xp33_ASAP7_75t_L g669 ( .A1(n_500), .A2(n_630), .A3(n_644), .B1(n_670), .B2(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
AND2x2_ASAP7_75t_L g610 ( .A(n_501), .B(n_554), .Y(n_610) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g592 ( .A(n_502), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_502), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g664 ( .A(n_502), .B(n_554), .Y(n_664) );
AND2x2_ASAP7_75t_L g675 ( .A(n_502), .B(n_567), .Y(n_675) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g576 ( .A(n_503), .B(n_555), .Y(n_576) );
AND2x2_ASAP7_75t_L g580 ( .A(n_503), .B(n_555), .Y(n_580) );
AND2x2_ASAP7_75t_L g615 ( .A(n_503), .B(n_566), .Y(n_615) );
AND2x2_ASAP7_75t_L g622 ( .A(n_503), .B(n_524), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g627 ( .A1(n_503), .A2(n_573), .B(n_584), .C(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g681 ( .A(n_503), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_503), .B(n_514), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_512), .B(n_564), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_512), .B(n_580), .Y(n_670) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g575 ( .A(n_513), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
AND2x2_ASAP7_75t_L g567 ( .A(n_514), .B(n_525), .Y(n_567) );
OR2x2_ASAP7_75t_L g582 ( .A(n_514), .B(n_525), .Y(n_582) );
AND2x2_ASAP7_75t_L g605 ( .A(n_514), .B(n_566), .Y(n_605) );
INVx1_ASAP7_75t_L g609 ( .A(n_514), .Y(n_609) );
AND2x2_ASAP7_75t_L g628 ( .A(n_514), .B(n_565), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_514), .A2(n_593), .B1(n_639), .B2(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_514), .B(n_681), .Y(n_705) );
AND2x2_ASAP7_75t_L g720 ( .A(n_514), .B(n_580), .Y(n_720) );
INVx4_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx3_ASAP7_75t_L g552 ( .A(n_515), .Y(n_552) );
AND2x2_ASAP7_75t_L g594 ( .A(n_515), .B(n_525), .Y(n_594) );
AND2x2_ASAP7_75t_L g596 ( .A(n_515), .B(n_554), .Y(n_596) );
AND3x2_ASAP7_75t_L g658 ( .A(n_515), .B(n_622), .C(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g693 ( .A(n_524), .B(n_565), .Y(n_693) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g554 ( .A(n_525), .B(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_525), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_525), .B(n_564), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_525), .B(n_605), .C(n_681), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_551), .B1(n_563), .B2(n_568), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_537), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g645 ( .A(n_537), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g661 ( .A1(n_540), .A2(n_662), .A3(n_663), .B(n_664), .Y(n_661) );
AND2x2_ASAP7_75t_L g686 ( .A(n_540), .B(n_573), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_540), .B(n_599), .Y(n_732) );
AND2x2_ASAP7_75t_L g641 ( .A(n_541), .B(n_573), .Y(n_641) );
AND2x2_ASAP7_75t_L g702 ( .A(n_541), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g572 ( .A(n_542), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g630 ( .A(n_542), .Y(n_630) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
CKINVDCx16_ASAP7_75t_R g651 ( .A(n_552), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_553), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AOI221x1_ASAP7_75t_SL g618 ( .A1(n_554), .A2(n_619), .B1(n_621), .B2(n_623), .C(n_625), .Y(n_618) );
INVx2_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_555), .Y(n_660) );
INVx1_ASAP7_75t_L g648 ( .A(n_563), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_564), .B(n_581), .Y(n_673) );
INVx1_ASAP7_75t_SL g736 ( .A(n_564), .Y(n_736) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g654 ( .A(n_567), .B(n_580), .Y(n_654) );
INVx1_ASAP7_75t_L g722 ( .A(n_568), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_568), .B(n_651), .Y(n_735) );
INVx2_ASAP7_75t_SL g574 ( .A(n_569), .Y(n_574) );
AND2x2_ASAP7_75t_L g617 ( .A(n_569), .B(n_573), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_569), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_569), .B(n_644), .Y(n_671) );
AOI21xp33_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_574), .B(n_575), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_572), .B(n_644), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_572), .B(n_599), .Y(n_740) );
OR2x2_ASAP7_75t_L g612 ( .A(n_573), .B(n_591), .Y(n_612) );
AND2x2_ASAP7_75t_L g711 ( .A(n_573), .B(n_702), .Y(n_711) );
OAI22xp5_ASAP7_75t_SL g586 ( .A1(n_574), .A2(n_587), .B1(n_592), .B2(n_595), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_574), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g634 ( .A(n_576), .B(n_582), .Y(n_634) );
INVx1_ASAP7_75t_L g698 ( .A(n_576), .Y(n_698) );
AOI311xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_583), .A3(n_585), .B(n_586), .C(n_597), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_581), .A2(n_713), .B1(n_725), .B2(n_728), .C(n_730), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_581), .B(n_736), .Y(n_738) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_584), .A2(n_626), .B(n_627), .C(n_629), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_SL g694 ( .A1(n_588), .A2(n_590), .B(n_695), .C(n_696), .Y(n_694) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_589), .B(n_663), .Y(n_729) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_592), .A2(n_612), .B1(n_613), .B2(n_616), .C(n_618), .Y(n_611) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g614 ( .A(n_594), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g697 ( .A(n_594), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_598), .A2(n_656), .B(n_657), .C(n_661), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_599), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_599), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVxp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g621 ( .A(n_605), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_609), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g723 ( .A(n_612), .Y(n_723) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_615), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g650 ( .A(n_615), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g727 ( .A(n_615), .Y(n_727) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g668 ( .A(n_617), .B(n_644), .Y(n_668) );
INVx1_ASAP7_75t_SL g662 ( .A(n_624), .Y(n_662) );
INVx1_ASAP7_75t_L g639 ( .A(n_630), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g631 ( .A(n_632), .B(n_649), .C(n_665), .Y(n_631) );
AOI322xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .A3(n_636), .B1(n_638), .B2(n_642), .C1(n_646), .C2(n_648), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_633), .A2(n_686), .B(n_687), .C(n_694), .Y(n_685) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_636), .A2(n_657), .B1(n_688), .B2(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g646 ( .A(n_644), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g683 ( .A(n_644), .B(n_684), .Y(n_683) );
AOI32xp33_ASAP7_75t_L g734 ( .A1(n_644), .A2(n_735), .A3(n_736), .B1(n_737), .B2(n_739), .Y(n_734) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g656 ( .A(n_647), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_647), .A2(n_700), .B1(n_704), .B2(n_706), .C(n_709), .Y(n_699) );
AND2x2_ASAP7_75t_L g713 ( .A(n_647), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g716 ( .A(n_651), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g726 ( .A(n_651), .B(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g717 ( .A(n_660), .B(n_681), .Y(n_717) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_669), .C(n_672), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI211xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_682), .B(n_685), .C(n_699), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_693), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g708 ( .A(n_705), .Y(n_708) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B(n_715), .Y(n_709) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI211xp5_ASAP7_75t_SL g718 ( .A1(n_719), .A2(n_721), .B(n_724), .C(n_734), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI21xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
BUFx4f_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
endmodule