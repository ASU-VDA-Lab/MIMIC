module fake_jpeg_28930_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_9),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_9),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_56),
.Y(n_70)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_36),
.Y(n_76)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_17),
.B1(n_29),
.B2(n_38),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_47),
.B1(n_17),
.B2(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_37),
.B1(n_27),
.B2(n_29),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_52),
.B1(n_55),
.B2(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_36),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_38),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_86),
.Y(n_117)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_103),
.B(n_53),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_52),
.B1(n_41),
.B2(n_55),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_100),
.B1(n_105),
.B2(n_51),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_26),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_118)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_66),
.B1(n_69),
.B2(n_47),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_31),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_22),
.B(n_23),
.C(n_34),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_22),
.C(n_23),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_28),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_48),
.B(n_45),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_49),
.B1(n_39),
.B2(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_31),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_59),
.B(n_34),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_99),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_89),
.B1(n_98),
.B2(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_131),
.B1(n_134),
.B2(n_87),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_105),
.B1(n_113),
.B2(n_96),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_67),
.B1(n_73),
.B2(n_68),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_68),
.B1(n_48),
.B2(n_47),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_97),
.B1(n_112),
.B2(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_51),
.B1(n_17),
.B2(n_32),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_97),
.B(n_88),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_87),
.B(n_103),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_154),
.B(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_152),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_150),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_153),
.B1(n_158),
.B2(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_94),
.C(n_82),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_109),
.B1(n_106),
.B2(n_84),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_140),
.B1(n_119),
.B2(n_122),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_88),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_85),
.B1(n_101),
.B2(n_93),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_32),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_137),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_30),
.B1(n_24),
.B2(n_80),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_24),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_78),
.C(n_30),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_0),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_169),
.B1(n_178),
.B2(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_129),
.B1(n_127),
.B2(n_134),
.Y(n_169)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_117),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_175),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_132),
.B1(n_136),
.B2(n_123),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_115),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_186),
.B1(n_155),
.B2(n_147),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_127),
.B(n_116),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_181),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_119),
.B1(n_122),
.B2(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

XOR2x2_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_135),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_130),
.B1(n_132),
.B2(n_137),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_138),
.B(n_33),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_189),
.B(n_138),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_130),
.B1(n_132),
.B2(n_33),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_145),
.A2(n_138),
.B(n_1),
.Y(n_189)
);

AND2x4_ASAP7_75t_SL g190 ( 
.A(n_188),
.B(n_154),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_201),
.B(n_208),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_186),
.B1(n_187),
.B2(n_168),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_147),
.B1(n_153),
.B2(n_148),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_198),
.B1(n_204),
.B2(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_161),
.B1(n_158),
.B2(n_164),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_156),
.C(n_164),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_165),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_164),
.B1(n_162),
.B2(n_152),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_150),
.B(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_184),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_138),
.B(n_1),
.Y(n_208)
);

AND2x4_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_0),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_203),
.C(n_202),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_187),
.B(n_199),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_183),
.B(n_169),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_201),
.B(n_195),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_224),
.B1(n_215),
.B2(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_190),
.B1(n_220),
.B2(n_182),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_207),
.B1(n_199),
.B2(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_10),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_242),
.C(n_225),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_203),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_240),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_181),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_177),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_209),
.B1(n_223),
.B2(n_216),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_185),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_251),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_212),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_221),
.B1(n_212),
.B2(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_235),
.C(n_240),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_209),
.B1(n_182),
.B2(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_171),
.B1(n_172),
.B2(n_3),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_171),
.B1(n_2),
.B2(n_4),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_238),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_256),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_255),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_242),
.B(n_229),
.C(n_0),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_11),
.B(n_2),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_246),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_264),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_243),
.B1(n_254),
.B2(n_249),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_274),
.C(n_12),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_244),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_267),
.A2(n_263),
.B(n_265),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_262),
.B(n_4),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_279),
.C(n_271),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_274),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_280),
.C(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

AOI321xp33_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_284),
.A3(n_7),
.B1(n_10),
.B2(n_13),
.C(n_15),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_289),
.A2(n_288),
.B(n_10),
.C(n_16),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_16),
.B(n_0),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_16),
.Y(n_292)
);


endmodule