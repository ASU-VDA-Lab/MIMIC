module fake_jpeg_15953_n_74 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_14),
.B1(n_22),
.B2(n_21),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_36),
.B(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_29),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_25),
.B(n_30),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_52),
.B(n_53),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_15),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_45),
.B(n_3),
.C(n_6),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_4),
.B(n_8),
.C(n_9),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_12),
.B(n_13),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_62),
.B(n_60),
.Y(n_68)
);

BUFx24_ASAP7_75t_SL g69 ( 
.A(n_68),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_67),
.CI(n_49),
.CON(n_70),
.SN(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_70),
.B(n_59),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_61),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);


endmodule