module fake_ariane_253_n_1772 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1772);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1772;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_1),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_55),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_42),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_54),
.B(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_43),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_70),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_24),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_93),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_134),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_46),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_56),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_58),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_57),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_53),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_65),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_84),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_68),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_78),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_108),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_39),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_114),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_47),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_2),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_157),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_35),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_62),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_59),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_40),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_85),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_123),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_48),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_104),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_26),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_29),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_122),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_15),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_135),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_96),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_118),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_0),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_59),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_158),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_61),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_89),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_51),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_9),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_76),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_47),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_17),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_81),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_44),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_88),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_97),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_52),
.Y(n_242)
);

BUFx2_ASAP7_75t_SL g243 ( 
.A(n_155),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_45),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_148),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_110),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_136),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_29),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_46),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_13),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_34),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_113),
.Y(n_259)
);

BUFx2_ASAP7_75t_SL g260 ( 
.A(n_16),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_156),
.Y(n_262)
);

BUFx8_ASAP7_75t_SL g263 ( 
.A(n_145),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_21),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_24),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_117),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_64),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_129),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_133),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_127),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_77),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_54),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_73),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_99),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_124),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g282 ( 
.A(n_44),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_32),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_91),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_19),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_82),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_52),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_106),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_139),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_41),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_144),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_57),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_151),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_126),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_121),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_132),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_25),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_72),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_33),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_2),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_87),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_95),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_147),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_55),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_42),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_143),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_152),
.Y(n_314)
);

BUFx2_ASAP7_75t_SL g315 ( 
.A(n_5),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_263),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_287),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_184),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_208),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_221),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_299),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_252),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_181),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_196),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_204),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_264),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_204),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_159),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_205),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_303),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_211),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_159),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_217),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_179),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_222),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_277),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_223),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_224),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_231),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_179),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_233),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_239),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_199),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_163),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_199),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_164),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_244),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_294),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_306),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_245),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_204),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_167),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_173),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_177),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_178),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_194),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_246),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_203),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_206),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_247),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_161),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_210),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_226),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_226),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_226),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_161),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_260),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_214),
.B(n_0),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_165),
.B(n_169),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_163),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_230),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_253),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_171),
.B(n_3),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_254),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_235),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_255),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_256),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_261),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_238),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_183),
.B(n_3),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_248),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_R g388 ( 
.A(n_160),
.B(n_102),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_257),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_197),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_265),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_195),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_331),
.B(n_266),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_197),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_202),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_291),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_202),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_240),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_386),
.B(n_182),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_345),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_348),
.B(n_240),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_297),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_351),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_351),
.A2(n_234),
.B(n_228),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_352),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_307),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_358),
.A2(n_273),
.B(n_250),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_213),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_274),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_364),
.B(n_207),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_364),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_328),
.B(n_182),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_368),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_376),
.B(n_328),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_320),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_220),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_322),
.Y(n_441)
);

CKINVDCx6p67_ASAP7_75t_R g442 ( 
.A(n_321),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_323),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_321),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_332),
.B(n_275),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_332),
.B(n_213),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_357),
.B(n_213),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_327),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_417),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_462),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_438),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_404),
.B(n_357),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_325),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_403),
.A2(n_317),
.B1(n_350),
.B2(n_369),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_403),
.A2(n_370),
.B1(n_371),
.B2(n_315),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_430),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_417),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_404),
.B(n_451),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_404),
.B(n_334),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_403),
.A2(n_462),
.B1(n_402),
.B2(n_424),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_455),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_336),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_404),
.B(n_338),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_340),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_342),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_343),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_462),
.A2(n_282),
.B1(n_242),
.B2(n_382),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_344),
.Y(n_490)
);

NOR2x1p5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_316),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_462),
.A2(n_384),
.B1(n_383),
.B2(n_380),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_438),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_425),
.Y(n_494)
);

BUFx6f_ASAP7_75t_SL g495 ( 
.A(n_463),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_207),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_346),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_462),
.B(n_347),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_207),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_426),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_424),
.B(n_353),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_462),
.B(n_356),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g507 ( 
.A(n_396),
.B(n_366),
.C(n_363),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_454),
.B(n_378),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_462),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_438),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_463),
.B(n_272),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_463),
.B(n_318),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_402),
.A2(n_175),
.B1(n_191),
.B2(n_220),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_393),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_393),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_463),
.B(n_276),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_438),
.B(n_460),
.C(n_459),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_232),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_431),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_433),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_424),
.B(n_434),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_393),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_463),
.B(n_319),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_456),
.B(n_279),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_459),
.A2(n_460),
.B1(n_355),
.B2(n_326),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_454),
.B(n_160),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_459),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_454),
.B(n_170),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_406),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_456),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_437),
.B(n_168),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_402),
.A2(n_243),
.B1(n_166),
.B2(n_278),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_421),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_396),
.B(n_281),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_406),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_406),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_454),
.B(n_170),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_421),
.B(n_436),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_432),
.A2(n_269),
.B1(n_270),
.B2(n_284),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_396),
.B(n_304),
.Y(n_552)
);

AND3x2_ASAP7_75t_L g553 ( 
.A(n_460),
.B(n_308),
.C(n_354),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_431),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_431),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_454),
.B(n_168),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_406),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_456),
.B(n_207),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_411),
.B(n_174),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_411),
.B(n_174),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_444),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_431),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_448),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_421),
.Y(n_566)
);

AND2x2_ASAP7_75t_SL g567 ( 
.A(n_460),
.B(n_207),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_406),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_411),
.B(n_185),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_406),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_448),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_411),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_406),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_448),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_448),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_432),
.A2(n_180),
.B1(n_176),
.B2(n_172),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_456),
.B(n_241),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_431),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_432),
.A2(n_189),
.B1(n_180),
.B2(n_176),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_411),
.B(n_185),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_456),
.B(n_241),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_411),
.B(n_186),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g584 ( 
.A(n_458),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_452),
.A2(n_341),
.B1(n_312),
.B2(n_311),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_458),
.B(n_186),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_411),
.B(n_187),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_442),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_445),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_456),
.B(n_187),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_402),
.B(n_188),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_406),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_445),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_394),
.B(n_172),
.Y(n_598)
);

INVxp33_ASAP7_75t_SL g599 ( 
.A(n_458),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_402),
.B(n_188),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_402),
.B(n_452),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_421),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_406),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_SL g604 ( 
.A1(n_437),
.A2(n_312),
.B1(n_311),
.B2(n_305),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_402),
.A2(n_189),
.B1(n_305),
.B2(n_301),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_421),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_402),
.A2(n_192),
.B1(n_285),
.B2(n_288),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_398),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_534),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_456),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_584),
.B(n_437),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_442),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_493),
.B(n_457),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_524),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_442),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_468),
.B(n_477),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_452),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_524),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_480),
.B(n_440),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_527),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_512),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_482),
.B(n_453),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_480),
.B(n_440),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_497),
.B(n_453),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_464),
.B(n_453),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_464),
.B(n_440),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_503),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_567),
.A2(n_442),
.B1(n_400),
.B2(n_440),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_554),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_478),
.A2(n_440),
.B1(n_419),
.B2(n_450),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_503),
.B(n_457),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_440),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_440),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_483),
.B(n_442),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_565),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_557),
.B(n_440),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_480),
.B(n_421),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_484),
.B(n_485),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_574),
.Y(n_642)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_469),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_470),
.B(n_400),
.C(n_427),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_575),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_486),
.B(n_400),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_490),
.B(n_400),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_480),
.B(n_436),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_557),
.B(n_395),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_557),
.B(n_395),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_476),
.B(n_395),
.Y(n_651)
);

AO221x1_ASAP7_75t_L g652 ( 
.A1(n_586),
.A2(n_461),
.B1(n_457),
.B2(n_241),
.C(n_262),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_473),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_567),
.A2(n_395),
.B1(n_427),
.B2(n_394),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_523),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_480),
.B(n_436),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_475),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_523),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_586),
.A2(n_461),
.B1(n_457),
.B2(n_427),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_489),
.B(n_436),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_534),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_467),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_489),
.B(n_436),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_489),
.B(n_466),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_494),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_508),
.B(n_392),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_521),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_513),
.B(n_392),
.C(n_285),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_541),
.B(n_395),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_471),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_498),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_541),
.B(n_395),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_491),
.B(n_457),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_586),
.B(n_461),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_489),
.B(n_436),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_489),
.B(n_436),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_500),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_502),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_481),
.B(n_461),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_505),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_466),
.B(n_608),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_536),
.B(n_461),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_594),
.A2(n_532),
.B1(n_517),
.B2(n_543),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_534),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_515),
.B(n_419),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_395),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_506),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_522),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_598),
.B(n_413),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_598),
.B(n_471),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_552),
.B(n_398),
.Y(n_691)
);

BUFx6f_ASAP7_75t_SL g692 ( 
.A(n_471),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_507),
.B(n_419),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_555),
.B(n_398),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_601),
.B(n_419),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_466),
.B(n_436),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_564),
.B(n_398),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_535),
.B(n_398),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_479),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_538),
.B(n_398),
.Y(n_700)
);

BUFx5_ASAP7_75t_L g701 ( 
.A(n_496),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_479),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_466),
.B(n_436),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_572),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_479),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_572),
.B(n_436),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_548),
.B(n_398),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_526),
.B(n_422),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_542),
.B(n_413),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_542),
.B(n_413),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_526),
.B(n_398),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_572),
.B(n_436),
.Y(n_712)
);

NAND2x1p5_ASAP7_75t_L g713 ( 
.A(n_608),
.B(n_401),
.Y(n_713)
);

AND2x6_ASAP7_75t_SL g714 ( 
.A(n_531),
.B(n_413),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_472),
.B(n_418),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_526),
.B(n_530),
.Y(n_716)
);

BUFx5_ASAP7_75t_L g717 ( 
.A(n_496),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_530),
.B(n_401),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_578),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_533),
.B(n_418),
.Y(n_721)
);

AND2x6_ASAP7_75t_L g722 ( 
.A(n_465),
.B(n_394),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_465),
.B(n_401),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_556),
.B(n_422),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_487),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_556),
.B(n_587),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_585),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_487),
.B(n_401),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_511),
.B(n_401),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_511),
.B(n_401),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_516),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_592),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_593),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_516),
.B(n_401),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_518),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_492),
.B(n_446),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_587),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_469),
.Y(n_740)
);

OAI22x1_ASAP7_75t_SL g741 ( 
.A1(n_467),
.A2(n_288),
.B1(n_192),
.B2(n_290),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_518),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_590),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_519),
.B(n_422),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_519),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_579),
.B(n_301),
.C(n_296),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_529),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_488),
.A2(n_450),
.B1(n_449),
.B2(n_447),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_509),
.B(n_446),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_520),
.A2(n_420),
.B(n_449),
.Y(n_750)
);

AOI221xp5_ASAP7_75t_L g751 ( 
.A1(n_586),
.A2(n_290),
.B1(n_296),
.B2(n_418),
.C(n_397),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_510),
.B(n_446),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_560),
.B(n_422),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_532),
.A2(n_418),
.B1(n_449),
.B2(n_447),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_562),
.B(n_423),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_510),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_604),
.B(n_405),
.C(n_449),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_520),
.A2(n_450),
.B1(n_449),
.B2(n_447),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_553),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_595),
.B(n_423),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_569),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_581),
.B(n_423),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_576),
.A2(n_450),
.B1(n_447),
.B2(n_423),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_510),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_600),
.A2(n_450),
.B1(n_447),
.B2(n_423),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_509),
.B(n_446),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_583),
.A2(n_428),
.B1(n_443),
.B2(n_439),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_589),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_539),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_510),
.B(n_446),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_605),
.B(n_428),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_514),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_616),
.A2(n_607),
.B1(n_495),
.B2(n_551),
.Y(n_773)
);

OA21x2_ASAP7_75t_L g774 ( 
.A1(n_750),
.A2(n_416),
.B(n_420),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_708),
.A2(n_504),
.B(n_499),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_653),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_616),
.B(n_499),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_716),
.A2(n_504),
.B(n_549),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_666),
.B(n_590),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_612),
.A2(n_495),
.B1(n_559),
.B2(n_577),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_661),
.B(n_514),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_657),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_681),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_666),
.B(n_428),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_646),
.B(n_428),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_611),
.B(n_428),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_716),
.A2(n_549),
.B(n_546),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_655),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_613),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_681),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_611),
.B(n_495),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_738),
.A2(n_416),
.B(n_420),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_710),
.B(n_429),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_610),
.A2(n_646),
.B(n_647),
.C(n_655),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_658),
.B(n_429),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_658),
.B(n_429),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_647),
.B(n_429),
.Y(n_797)
);

NOR2x1_ASAP7_75t_R g798 ( 
.A(n_702),
.B(n_190),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_679),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_696),
.A2(n_546),
.B(n_539),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_725),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_612),
.A2(n_582),
.B1(n_577),
.B2(n_559),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_665),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_632),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_732),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_703),
.A2(n_648),
.B(n_639),
.Y(n_806)
);

OAI321xp33_ASAP7_75t_L g807 ( 
.A1(n_751),
.A2(n_408),
.A3(n_410),
.B1(n_409),
.B2(n_407),
.C(n_415),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_661),
.B(n_514),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_737),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_681),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_640),
.B(n_429),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_671),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_703),
.A2(n_550),
.B(n_547),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_639),
.A2(n_550),
.B(n_547),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_708),
.A2(n_561),
.B(n_603),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_648),
.A2(n_568),
.B(n_603),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_640),
.B(n_435),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_617),
.A2(n_439),
.B(n_443),
.C(n_435),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_622),
.A2(n_540),
.B1(n_568),
.B2(n_596),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_644),
.A2(n_420),
.B(n_416),
.C(n_435),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_615),
.B(n_540),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_681),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_677),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_656),
.A2(n_558),
.B(n_596),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_624),
.A2(n_629),
.B1(n_683),
.B2(n_633),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_621),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_656),
.A2(n_558),
.B(n_573),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_760),
.A2(n_573),
.B(n_561),
.Y(n_828)
);

OAI321xp33_ASAP7_75t_L g829 ( 
.A1(n_674),
.A2(n_410),
.A3(n_407),
.B1(n_408),
.B2(n_409),
.C(n_399),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_742),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_615),
.B(n_559),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_628),
.B(n_540),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_690),
.B(n_435),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_636),
.B(n_435),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_684),
.B(n_704),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_660),
.A2(n_570),
.B(n_602),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_660),
.A2(n_570),
.B(n_602),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_692),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_SL g839 ( 
.A(n_692),
.B(n_514),
.Y(n_839)
);

AOI21x1_ASAP7_75t_L g840 ( 
.A1(n_619),
.A2(n_420),
.B(n_416),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_681),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_689),
.B(n_721),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_636),
.B(n_439),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_609),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_614),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_663),
.A2(n_602),
.B(n_537),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_618),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_625),
.B(n_439),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_695),
.A2(n_416),
.B(n_443),
.C(n_439),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_760),
.A2(n_525),
.B(n_501),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_693),
.A2(n_525),
.B(n_410),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_745),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_709),
.B(n_443),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_761),
.B(n_443),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_662),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_663),
.A2(n_602),
.B(n_537),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_682),
.B(n_405),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_675),
.A2(n_537),
.B(n_566),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_740),
.B(n_643),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_768),
.B(n_405),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_695),
.A2(n_496),
.B(n_501),
.Y(n_861)
);

INVx5_ASAP7_75t_L g862 ( 
.A(n_722),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_684),
.B(n_537),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_675),
.A2(n_606),
.B(n_566),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_756),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_676),
.A2(n_606),
.B(n_566),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_715),
.B(n_654),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_626),
.A2(n_606),
.B1(n_566),
.B2(n_544),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_682),
.B(n_405),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_609),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_676),
.A2(n_606),
.B(n_566),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_722),
.B(n_405),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_747),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_635),
.A2(n_405),
.B(n_407),
.C(n_408),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_619),
.A2(n_501),
.B(n_496),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_722),
.B(n_405),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_714),
.B(n_397),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_686),
.A2(n_606),
.B1(n_544),
.B2(n_446),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_704),
.B(n_544),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_746),
.A2(n_409),
.B(n_410),
.C(n_407),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_749),
.A2(n_544),
.B(n_501),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_667),
.B(n_474),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_749),
.A2(n_544),
.B(n_501),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_766),
.A2(n_501),
.B(n_496),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_685),
.B(n_559),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_668),
.B(n_397),
.Y(n_886)
);

AO21x1_ASAP7_75t_L g887 ( 
.A1(n_693),
.A2(n_399),
.B(n_415),
.Y(n_887)
);

NOR2x1_ASAP7_75t_R g888 ( 
.A(n_670),
.B(n_190),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_766),
.A2(n_755),
.B(n_753),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_769),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_642),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_673),
.B(n_474),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_620),
.B(n_446),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_623),
.A2(n_496),
.B(n_582),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_711),
.A2(n_582),
.B(n_577),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_649),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_739),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_756),
.B(n_446),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_645),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_678),
.B(n_582),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_762),
.A2(n_446),
.B(n_193),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_664),
.A2(n_412),
.B(n_582),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_744),
.A2(n_446),
.B(n_193),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_680),
.B(n_582),
.Y(n_904)
);

BUFx4f_ASAP7_75t_L g905 ( 
.A(n_673),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_687),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_638),
.A2(n_412),
.B(n_414),
.C(n_313),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_743),
.B(n_412),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_664),
.A2(n_412),
.B(n_232),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_688),
.B(n_412),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_673),
.B(n_474),
.Y(n_911)
);

NOR2x1_ASAP7_75t_L g912 ( 
.A(n_627),
.B(n_414),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_756),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_691),
.B(n_414),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_740),
.B(n_414),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_718),
.A2(n_236),
.B(n_237),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_630),
.B(n_414),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_659),
.A2(n_236),
.B1(n_237),
.B2(n_286),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_699),
.B(n_414),
.Y(n_919)
);

AO21x1_ASAP7_75t_L g920 ( 
.A1(n_738),
.A2(n_232),
.B(n_414),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_651),
.A2(n_286),
.B(n_289),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_705),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_713),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_698),
.A2(n_289),
.B(n_292),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_726),
.A2(n_724),
.B1(n_672),
.B2(n_669),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_SL g926 ( 
.A(n_759),
.B(n_292),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_634),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_650),
.A2(n_293),
.B1(n_295),
.B2(n_298),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_700),
.A2(n_293),
.B(n_295),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_637),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_641),
.B(n_414),
.Y(n_931)
);

AO21x1_ASAP7_75t_L g932 ( 
.A1(n_763),
.A2(n_232),
.B(n_414),
.Y(n_932)
);

NOR2x1_ASAP7_75t_L g933 ( 
.A(n_694),
.B(n_241),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_707),
.A2(n_298),
.B(n_300),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_697),
.B(n_300),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_756),
.B(n_474),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_739),
.B(n_302),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_706),
.A2(n_302),
.B(n_314),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_723),
.A2(n_4),
.B(n_8),
.C(n_10),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_764),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_713),
.B(n_719),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_712),
.A2(n_310),
.B(n_313),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_712),
.A2(n_229),
.B(n_200),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_770),
.A2(n_198),
.B(n_212),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_720),
.Y(n_945)
);

AOI21x1_ASAP7_75t_L g946 ( 
.A1(n_770),
.A2(n_730),
.B(n_736),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_724),
.B(n_201),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_727),
.A2(n_209),
.B(n_215),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_764),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_674),
.B(n_8),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_731),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_779),
.A2(n_631),
.B1(n_734),
.B2(n_733),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_791),
.A2(n_631),
.B1(n_735),
.B2(n_772),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_786),
.B(n_674),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_838),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_SL g956 ( 
.A1(n_826),
.A2(n_741),
.B1(n_771),
.B2(n_754),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_887),
.A2(n_729),
.B(n_728),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_834),
.A2(n_752),
.B(n_764),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_791),
.A2(n_821),
.B1(n_773),
.B2(n_817),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_842),
.B(n_757),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_794),
.A2(n_763),
.B(n_748),
.C(n_765),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_843),
.A2(n_772),
.B(n_764),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_825),
.A2(n_748),
.B(n_767),
.C(n_652),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_804),
.B(n_772),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_838),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_776),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_788),
.B(n_789),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_811),
.A2(n_772),
.B(n_758),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_905),
.B(n_701),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_833),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_784),
.A2(n_717),
.B(n_701),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_782),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_804),
.B(n_717),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_862),
.B(n_701),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_833),
.A2(n_12),
.B(n_14),
.C(n_17),
.Y(n_975)
);

BUFx8_ASAP7_75t_SL g976 ( 
.A(n_855),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_777),
.A2(n_717),
.B(n_701),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_SL g978 ( 
.A1(n_821),
.A2(n_717),
.B(n_701),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_896),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_889),
.A2(n_717),
.B(n_701),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_803),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_945),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_785),
.A2(n_14),
.B(n_18),
.C(n_19),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_789),
.B(n_717),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_812),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_797),
.A2(n_241),
.B(n_309),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_892),
.B(n_18),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_799),
.B(n_20),
.Y(n_988)
);

OAI22x1_ASAP7_75t_L g989 ( 
.A1(n_918),
.A2(n_225),
.B1(n_227),
.B2(n_249),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_823),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_928),
.A2(n_251),
.B(n_259),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_891),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_826),
.B(n_267),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_810),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_799),
.B(n_20),
.Y(n_995)
);

CKINVDCx8_ASAP7_75t_R g996 ( 
.A(n_892),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_951),
.Y(n_997)
);

AOI33xp33_ASAP7_75t_L g998 ( 
.A1(n_899),
.A2(n_21),
.A3(n_22),
.B1(n_23),
.B2(n_26),
.B3(n_27),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_810),
.B(n_262),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_783),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_783),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_853),
.B(n_28),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_L g1003 ( 
.A(n_783),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_822),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_915),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_795),
.B(n_30),
.Y(n_1006)
);

BUFx2_ASAP7_75t_R g1007 ( 
.A(n_950),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_874),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_927),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_783),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_796),
.B(n_31),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_862),
.B(n_280),
.Y(n_1012)
);

INVx5_ASAP7_75t_L g1013 ( 
.A(n_822),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_841),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_793),
.B(n_896),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_859),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_857),
.B(n_34),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_930),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_857),
.B(n_35),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_839),
.B(n_283),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_909),
.A2(n_232),
.B(n_309),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_841),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_925),
.A2(n_309),
.B(n_271),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_905),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_790),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_SL g1026 ( 
.A1(n_877),
.A2(n_262),
.B1(n_271),
.B2(n_309),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_941),
.A2(n_862),
.B1(n_935),
.B2(n_867),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_908),
.B(n_36),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_862),
.A2(n_262),
.B1(n_271),
.B2(n_38),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_926),
.B(n_232),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_877),
.B(n_36),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_923),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_878),
.A2(n_271),
.B(n_232),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_828),
.A2(n_232),
.B(n_430),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_SL g1035 ( 
.A1(n_922),
.A2(n_37),
.B1(n_41),
.B2(n_48),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_815),
.A2(n_430),
.B(n_50),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_831),
.B(n_49),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_775),
.A2(n_430),
.B(n_51),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_923),
.B(n_50),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_869),
.A2(n_56),
.B1(n_60),
.B2(n_430),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_886),
.A2(n_430),
.B(n_60),
.C(n_66),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_778),
.A2(n_430),
.B(n_71),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_906),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_809),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_911),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_947),
.A2(n_430),
.B1(n_74),
.B2(n_75),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_911),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_888),
.B(n_63),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_830),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_937),
.A2(n_430),
.B1(n_90),
.B2(n_98),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_937),
.B(n_430),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_807),
.A2(n_430),
.B1(n_103),
.B2(n_111),
.C(n_112),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_886),
.B(n_430),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_852),
.B(n_430),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_882),
.B(n_86),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_914),
.A2(n_430),
.B(n_119),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_897),
.B(n_430),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_845),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_829),
.B(n_115),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_902),
.A2(n_130),
.B(n_140),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_873),
.B(n_141),
.Y(n_1061)
);

OAI22x1_ASAP7_75t_L g1062 ( 
.A1(n_847),
.A2(n_780),
.B1(n_802),
.B2(n_801),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_874),
.A2(n_880),
.B(n_939),
.C(n_854),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_830),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_868),
.A2(n_850),
.B(n_849),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_849),
.A2(n_861),
.B(n_787),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_832),
.B(n_897),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_805),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_832),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_890),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_910),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_882),
.B(n_848),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_917),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_860),
.A2(n_844),
.B1(n_870),
.B2(n_872),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_798),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_835),
.B(n_948),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_790),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_844),
.B(n_870),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_865),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_919),
.B(n_938),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_865),
.B(n_913),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_865),
.B(n_913),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_839),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_814),
.A2(n_816),
.B(n_827),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_819),
.A2(n_806),
.B(n_800),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_876),
.B(n_835),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_865),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_781),
.A2(n_863),
.B(n_808),
.C(n_879),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_913),
.B(n_949),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_913),
.B(n_949),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_949),
.B(n_940),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_949),
.B(n_940),
.Y(n_1092)
);

O2A1O1Ixp5_ASAP7_75t_L g1093 ( 
.A1(n_851),
.A2(n_932),
.B(n_781),
.C(n_808),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_824),
.A2(n_813),
.B(n_837),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_936),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_836),
.A2(n_864),
.B(n_871),
.Y(n_1096)
);

INVx3_ASAP7_75t_SL g1097 ( 
.A(n_936),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_931),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_863),
.B(n_879),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_921),
.B(n_942),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_967),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_959),
.A2(n_924),
.B(n_929),
.C(n_934),
.Y(n_1102)
);

INVx3_ASAP7_75t_SL g1103 ( 
.A(n_965),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_961),
.A2(n_1076),
.B(n_963),
.C(n_1052),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_976),
.B(n_943),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1015),
.B(n_944),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1016),
.B(n_893),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_980),
.A2(n_920),
.B(n_866),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_970),
.A2(n_907),
.B(n_818),
.C(n_916),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_1003),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_966),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1023),
.A2(n_1065),
.B(n_1085),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_972),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_1003),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1023),
.A2(n_820),
.B(n_901),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_960),
.B(n_893),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_981),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_987),
.B(n_820),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_975),
.A2(n_933),
.B(n_885),
.C(n_894),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_980),
.A2(n_858),
.B(n_856),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_SL g1121 ( 
.A1(n_1059),
.A2(n_898),
.B(n_895),
.C(n_904),
.Y(n_1121)
);

OAI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_998),
.A2(n_912),
.B(n_903),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1084),
.A2(n_846),
.B(n_883),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_985),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1096),
.A2(n_881),
.B(n_946),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_993),
.B(n_898),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_1032),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1028),
.B(n_792),
.Y(n_1128)
);

AOI221x1_ASAP7_75t_L g1129 ( 
.A1(n_1038),
.A2(n_884),
.B1(n_875),
.B2(n_900),
.C(n_792),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1065),
.A2(n_774),
.B(n_792),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1096),
.A2(n_840),
.B(n_774),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_990),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_SL g1133 ( 
.A1(n_975),
.A2(n_774),
.B1(n_1008),
.B2(n_983),
.C(n_1038),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_1067),
.A2(n_1017),
.B(n_1019),
.C(n_1086),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1085),
.A2(n_1066),
.B(n_958),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1075),
.B(n_988),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1069),
.B(n_1001),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1099),
.A2(n_1041),
.B(n_1051),
.C(n_1078),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1036),
.A2(n_1063),
.B(n_1100),
.C(n_1008),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_SL g1140 ( 
.A1(n_983),
.A2(n_1036),
.B(n_1048),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1024),
.B(n_992),
.Y(n_1141)
);

AO21x2_ASAP7_75t_L g1142 ( 
.A1(n_1066),
.A2(n_986),
.B(n_1094),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1002),
.A2(n_952),
.B1(n_954),
.B2(n_1006),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_958),
.A2(n_968),
.B(n_1094),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1047),
.B(n_1045),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1093),
.A2(n_968),
.B(n_1063),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1011),
.A2(n_953),
.B1(n_995),
.B2(n_1035),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1021),
.A2(n_962),
.B(n_1060),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1053),
.A2(n_962),
.B(n_1034),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1001),
.B(n_1055),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_955),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1062),
.A2(n_986),
.A3(n_1027),
.B(n_1033),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_971),
.A2(n_978),
.B(n_977),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_971),
.A2(n_977),
.B(n_1033),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1058),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1001),
.B(n_1055),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1088),
.A2(n_1074),
.B(n_1072),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1009),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_982),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1022),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_989),
.A2(n_1039),
.B1(n_1029),
.B2(n_1083),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1018),
.Y(n_1162)
);

INVx8_ASAP7_75t_L g1163 ( 
.A(n_1001),
.Y(n_1163)
);

AOI221xp5_ASAP7_75t_L g1164 ( 
.A1(n_991),
.A2(n_979),
.B1(n_1040),
.B2(n_1026),
.C(n_1050),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1042),
.A2(n_957),
.B(n_1056),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1042),
.A2(n_1056),
.B(n_1061),
.Y(n_1166)
);

O2A1O1Ixp5_ASAP7_75t_L g1167 ( 
.A1(n_1037),
.A2(n_1012),
.B(n_1089),
.C(n_1090),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1069),
.B(n_1022),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_964),
.Y(n_1169)
);

AOI222xp33_ASAP7_75t_L g1170 ( 
.A1(n_1043),
.A2(n_997),
.B1(n_1005),
.B2(n_1071),
.C1(n_1095),
.C2(n_1007),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1022),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_994),
.B(n_1022),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1079),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_974),
.A2(n_1081),
.B(n_1082),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_996),
.B(n_1070),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_973),
.Y(n_1176)
);

AOI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_1046),
.A2(n_1080),
.B1(n_1030),
.B2(n_1073),
.C(n_984),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1068),
.Y(n_1178)
);

OA22x2_ASAP7_75t_L g1179 ( 
.A1(n_1097),
.A2(n_999),
.B1(n_1091),
.B2(n_1092),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1044),
.A2(n_1064),
.B1(n_1049),
.B2(n_1098),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_SL g1181 ( 
.A1(n_999),
.A2(n_1000),
.B(n_1010),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1004),
.A2(n_1025),
.B(n_1077),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1004),
.A2(n_1025),
.B(n_1077),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_994),
.A2(n_969),
.B(n_1054),
.C(n_1087),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1087),
.B(n_1079),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_L g1186 ( 
.A1(n_1020),
.A2(n_1079),
.B(n_1057),
.C(n_1013),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_999),
.A2(n_1014),
.B(n_1000),
.C(n_1010),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1000),
.B(n_1010),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1031),
.A2(n_467),
.B1(n_611),
.B2(n_612),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1065),
.A2(n_920),
.A3(n_887),
.B(n_932),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_L g1191 ( 
.A(n_959),
.B(n_403),
.C(n_773),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_966),
.Y(n_1192)
);

NAND2x1p5_ASAP7_75t_L g1193 ( 
.A(n_1003),
.B(n_810),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_959),
.A2(n_779),
.B(n_531),
.C(n_515),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_959),
.A2(n_779),
.B(n_531),
.C(n_515),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_967),
.B(n_611),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1038),
.A2(n_959),
.B1(n_1023),
.B2(n_1036),
.C(n_1065),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_959),
.A2(n_779),
.B(n_531),
.C(n_515),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1024),
.B(n_892),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_SL g1202 ( 
.A(n_955),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_980),
.A2(n_1084),
.B(n_1096),
.Y(n_1203)
);

OR2x6_ASAP7_75t_L g1204 ( 
.A(n_1055),
.B(n_810),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1015),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_959),
.A2(n_773),
.B(n_1027),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1003),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_960),
.B(n_867),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_980),
.A2(n_1084),
.B(n_1096),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_967),
.B(n_611),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_980),
.A2(n_1084),
.B(n_1096),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_982),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_SL g1215 ( 
.A(n_959),
.B(n_822),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1066),
.A2(n_1065),
.B(n_1096),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1023),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_965),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_960),
.B(n_867),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_959),
.A2(n_1023),
.B(n_825),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1221)
);

AO32x2_ASAP7_75t_L g1222 ( 
.A1(n_959),
.A2(n_1027),
.A3(n_956),
.B1(n_825),
.B2(n_952),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_967),
.B(n_611),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_976),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_959),
.A2(n_1023),
.B(n_825),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_976),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1003),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_967),
.B(n_611),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_959),
.A2(n_1023),
.B(n_825),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_959),
.A2(n_1023),
.B(n_825),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_967),
.B(n_611),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1065),
.A2(n_920),
.A3(n_887),
.B(n_932),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_959),
.A2(n_779),
.B(n_531),
.C(n_515),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_967),
.B(n_788),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_959),
.A2(n_489),
.B(n_480),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_966),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_980),
.A2(n_1084),
.B(n_1096),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1111),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1191),
.A2(n_1147),
.B1(n_1170),
.B2(n_1189),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1191),
.A2(n_1147),
.B1(n_1170),
.B2(n_1206),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1207),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1113),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1117),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1208),
.A2(n_1219),
.B1(n_1143),
.B2(n_1231),
.Y(n_1248)
);

BUFx5_ASAP7_75t_L g1249 ( 
.A(n_1172),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1150),
.B(n_1156),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1208),
.A2(n_1219),
.B1(n_1143),
.B2(n_1230),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1124),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1204),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1136),
.A2(n_1232),
.B1(n_1223),
.B2(n_1196),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1215),
.A2(n_1118),
.B1(n_1231),
.B2(n_1220),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1132),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1215),
.A2(n_1220),
.B1(n_1225),
.B2(n_1230),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1210),
.A2(n_1228),
.B1(n_1140),
.B2(n_1194),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1140),
.A2(n_1161),
.B1(n_1164),
.B2(n_1126),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1195),
.A2(n_1237),
.B(n_1199),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1213),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1225),
.A2(n_1205),
.B1(n_1101),
.B2(n_1204),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1101),
.A2(n_1204),
.B1(n_1116),
.B2(n_1162),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1238),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1224),
.Y(n_1265)
);

INVx8_ASAP7_75t_L g1266 ( 
.A(n_1163),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1116),
.A2(n_1158),
.B1(n_1192),
.B2(n_1240),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1179),
.A2(n_1222),
.B1(n_1150),
.B2(n_1156),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1151),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1226),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1145),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1139),
.A2(n_1198),
.B(n_1104),
.Y(n_1272)
);

BUFx4f_ASAP7_75t_SL g1273 ( 
.A(n_1103),
.Y(n_1273)
);

INVx5_ASAP7_75t_L g1274 ( 
.A(n_1163),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1178),
.A2(n_1179),
.B1(n_1146),
.B2(n_1107),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1146),
.A2(n_1155),
.B1(n_1127),
.B2(n_1122),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1110),
.Y(n_1277)
);

BUFx4_ASAP7_75t_R g1278 ( 
.A(n_1222),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1173),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1169),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1207),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1127),
.A2(n_1177),
.B1(n_1115),
.B2(n_1128),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1141),
.Y(n_1283)
);

INVx6_ASAP7_75t_L g1284 ( 
.A(n_1207),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1175),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1105),
.A2(n_1109),
.B(n_1112),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1110),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1201),
.B(n_1114),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1201),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1222),
.A2(n_1106),
.B1(n_1115),
.B2(n_1227),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1157),
.A2(n_1102),
.B(n_1135),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1185),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1163),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1227),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1114),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1188),
.B(n_1137),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1202),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1180),
.A2(n_1217),
.B1(n_1202),
.B2(n_1149),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1119),
.A2(n_1168),
.B1(n_1239),
.B2(n_1197),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1193),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1193),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1134),
.B(n_1172),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1174),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1176),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1133),
.A2(n_1149),
.B1(n_1130),
.B2(n_1214),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1217),
.A2(n_1133),
.B1(n_1142),
.B2(n_1216),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1187),
.B(n_1181),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1200),
.A2(n_1211),
.B1(n_1236),
.B2(n_1233),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1186),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1138),
.B(n_1183),
.Y(n_1311)
);

BUFx2_ASAP7_75t_SL g1312 ( 
.A(n_1160),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1184),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1221),
.A2(n_1229),
.B1(n_1234),
.B2(n_1129),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1167),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1216),
.B(n_1171),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1190),
.B(n_1235),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1144),
.A2(n_1154),
.B1(n_1153),
.B2(n_1121),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1142),
.A2(n_1166),
.B1(n_1165),
.B2(n_1108),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1125),
.A2(n_1131),
.B1(n_1148),
.B2(n_1123),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1120),
.A2(n_1209),
.B1(n_1212),
.B2(n_1203),
.Y(n_1321)
);

BUFx4f_ASAP7_75t_SL g1322 ( 
.A(n_1190),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1235),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1241),
.A2(n_1152),
.B1(n_1189),
.B2(n_467),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1111),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1159),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1111),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1328)
);

BUFx8_ASAP7_75t_L g1329 ( 
.A(n_1202),
.Y(n_1329)
);

INVx6_ASAP7_75t_L g1330 ( 
.A(n_1207),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1159),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1218),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1159),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1147),
.A2(n_674),
.B1(n_586),
.B2(n_318),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1202),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1196),
.B(n_1223),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1111),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1147),
.A2(n_674),
.B1(n_586),
.B2(n_318),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1189),
.A2(n_779),
.B1(n_1191),
.B2(n_1147),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1189),
.A2(n_467),
.B1(n_615),
.B2(n_612),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1111),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_R g1346 ( 
.A1(n_1136),
.A2(n_611),
.B1(n_542),
.B2(n_481),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1224),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1189),
.A2(n_531),
.B(n_515),
.Y(n_1349)
);

OAI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1189),
.A2(n_1191),
.B1(n_1147),
.B2(n_674),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1189),
.A2(n_1191),
.B1(n_1147),
.B2(n_674),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1145),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1189),
.A2(n_467),
.B1(n_615),
.B2(n_612),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1159),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1207),
.Y(n_1355)
);

CKINVDCx6p67_ASAP7_75t_R g1356 ( 
.A(n_1103),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1191),
.A2(n_674),
.B1(n_659),
.B2(n_751),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1110),
.Y(n_1358)
);

BUFx8_ASAP7_75t_SL g1359 ( 
.A(n_1224),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1196),
.B(n_1223),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1150),
.B(n_1001),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1218),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1189),
.A2(n_1191),
.B1(n_1147),
.B2(n_674),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1145),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1196),
.B(n_1223),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1242),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1264),
.B(n_1317),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1246),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1306),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1318),
.A2(n_1319),
.B(n_1321),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1303),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1283),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1280),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1342),
.A2(n_1278),
.B1(n_1341),
.B2(n_1334),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1303),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1299),
.A2(n_1316),
.A3(n_1311),
.B(n_1258),
.Y(n_1377)
);

CKINVDCx16_ASAP7_75t_R g1378 ( 
.A(n_1265),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1319),
.A2(n_1321),
.B(n_1320),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1247),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1252),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1256),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1322),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1325),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1327),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1293),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1340),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1345),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1323),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1243),
.A2(n_1346),
.B1(n_1244),
.B2(n_1363),
.Y(n_1390)
);

NOR2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1356),
.B(n_1271),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1365),
.B(n_1248),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1337),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1394)
);

BUFx2_ASAP7_75t_SL g1395 ( 
.A(n_1274),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1360),
.B(n_1259),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1359),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1292),
.B(n_1267),
.Y(n_1398)
);

AOI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1313),
.A2(n_1302),
.B(n_1296),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1290),
.B(n_1267),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1322),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1290),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1305),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1291),
.A2(n_1272),
.B(n_1307),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1278),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1261),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1326),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1331),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1333),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1354),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1279),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1307),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1304),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1347),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1286),
.A2(n_1320),
.B(n_1260),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1310),
.B(n_1253),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1310),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1310),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1275),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1309),
.A2(n_1349),
.B(n_1351),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1350),
.A2(n_1351),
.B1(n_1328),
.B2(n_1357),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1343),
.A2(n_1353),
.B1(n_1344),
.B2(n_1357),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1324),
.B(n_1282),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_SL g1424 ( 
.A(n_1335),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1275),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1298),
.Y(n_1426)
);

INVxp33_ASAP7_75t_L g1427 ( 
.A(n_1254),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1298),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1282),
.A2(n_1262),
.B(n_1276),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1249),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1262),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1285),
.B(n_1364),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1312),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1314),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1328),
.A2(n_1344),
.B1(n_1338),
.B2(n_1339),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1314),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1263),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1336),
.A2(n_1338),
.B1(n_1348),
.B2(n_1339),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1263),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1308),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1352),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1309),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1276),
.B(n_1315),
.C(n_1336),
.Y(n_1443)
);

BUFx2_ASAP7_75t_SL g1444 ( 
.A(n_1274),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1352),
.B(n_1289),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1295),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1348),
.A2(n_1268),
.B1(n_1358),
.B2(n_1277),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1288),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1249),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1249),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1392),
.B(n_1249),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1373),
.A2(n_1390),
.B(n_1422),
.C(n_1420),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1411),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1411),
.B(n_1269),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1421),
.A2(n_1287),
.B1(n_1294),
.B2(n_1277),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1438),
.A2(n_1287),
.B1(n_1273),
.B2(n_1250),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1372),
.B(n_1335),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1373),
.A2(n_1270),
.B(n_1361),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1440),
.B(n_1273),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1435),
.A2(n_1245),
.B1(n_1355),
.B2(n_1330),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1440),
.B(n_1329),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1394),
.B(n_1297),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1375),
.A2(n_1245),
.B1(n_1330),
.B2(n_1355),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1446),
.B(n_1329),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1443),
.A2(n_1245),
.B1(n_1355),
.B2(n_1281),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1415),
.A2(n_1300),
.B(n_1301),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1377),
.B(n_1404),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1381),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1415),
.B(n_1403),
.C(n_1404),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1367),
.B(n_1332),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1393),
.B(n_1362),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1423),
.A2(n_1266),
.B1(n_1284),
.B2(n_1402),
.C(n_1425),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_SL g1473 ( 
.A1(n_1415),
.A2(n_1284),
.B(n_1398),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1383),
.B(n_1401),
.Y(n_1474)
);

OAI211xp5_ASAP7_75t_L g1475 ( 
.A1(n_1403),
.A2(n_1415),
.B(n_1404),
.C(n_1436),
.Y(n_1475)
);

INVx5_ASAP7_75t_L g1476 ( 
.A(n_1416),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1377),
.B(n_1404),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1432),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1400),
.A2(n_1427),
.B1(n_1396),
.B2(n_1429),
.Y(n_1479)
);

OAI21xp33_ASAP7_75t_L g1480 ( 
.A1(n_1434),
.A2(n_1436),
.B(n_1402),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1448),
.B(n_1380),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1419),
.A2(n_1425),
.B(n_1447),
.C(n_1434),
.Y(n_1482)
);

O2A1O1Ixp5_ASAP7_75t_SL g1483 ( 
.A1(n_1433),
.A2(n_1413),
.B(n_1442),
.C(n_1412),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1389),
.B(n_1430),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1370),
.A2(n_1379),
.B(n_1442),
.Y(n_1485)
);

NAND4xp25_ASAP7_75t_SL g1486 ( 
.A(n_1397),
.B(n_1419),
.C(n_1405),
.D(n_1426),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1399),
.B(n_1417),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_SL g1488 ( 
.A1(n_1441),
.A2(n_1414),
.B(n_1417),
.C(n_1418),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1429),
.A2(n_1391),
.B1(n_1378),
.B2(n_1428),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1429),
.A2(n_1418),
.B1(n_1431),
.B2(n_1439),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1491)
);

CKINVDCx14_ASAP7_75t_R g1492 ( 
.A(n_1414),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1376),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_1384),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1376),
.Y(n_1495)
);

CKINVDCx14_ASAP7_75t_R g1496 ( 
.A(n_1386),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1413),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1429),
.A2(n_1424),
.B1(n_1395),
.B2(n_1444),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1453),
.Y(n_1499)
);

OAI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1452),
.A2(n_1439),
.B1(n_1437),
.B2(n_1399),
.C(n_1389),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1493),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_1450),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1467),
.B(n_1450),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1477),
.B(n_1451),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1451),
.B(n_1377),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1494),
.B(n_1377),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1497),
.B(n_1377),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1485),
.B(n_1369),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1484),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1468),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1489),
.B(n_1371),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1475),
.B(n_1385),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1469),
.A2(n_1424),
.B1(n_1416),
.B2(n_1387),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1491),
.B(n_1385),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1452),
.A2(n_1382),
.B1(n_1387),
.B2(n_1388),
.C(n_1369),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1481),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1453),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1483),
.B(n_1382),
.C(n_1388),
.Y(n_1518)
);

NAND2x1_ASAP7_75t_L g1519 ( 
.A(n_1493),
.B(n_1430),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1376),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1479),
.A2(n_1408),
.B1(n_1410),
.B2(n_1406),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1478),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1485),
.B(n_1449),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1485),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1487),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1480),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1484),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1473),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1479),
.A2(n_1406),
.B1(n_1407),
.B2(n_1409),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1500),
.A2(n_1462),
.B1(n_1486),
.B2(n_1455),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1500),
.A2(n_1462),
.B1(n_1463),
.B2(n_1490),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1507),
.Y(n_1532)
);

AO21x2_ASAP7_75t_L g1533 ( 
.A1(n_1524),
.A2(n_1482),
.B(n_1466),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1505),
.B(n_1495),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1524),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1524),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1508),
.B(n_1505),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1513),
.A2(n_1492),
.B1(n_1498),
.B2(n_1496),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1508),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1523),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1512),
.A2(n_1458),
.B1(n_1456),
.B2(n_1482),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1508),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1505),
.B(n_1504),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1523),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1510),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1519),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1502),
.Y(n_1549)
);

NAND4xp25_ASAP7_75t_SL g1550 ( 
.A(n_1513),
.B(n_1492),
.C(n_1464),
.D(n_1471),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1502),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1504),
.B(n_1506),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1374),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1502),
.B(n_1474),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1528),
.B(n_1459),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1518),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1512),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1515),
.B(n_1459),
.C(n_1472),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_L g1559 ( 
.A1(n_1515),
.A2(n_1461),
.B(n_1460),
.C(n_1457),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1543),
.B(n_1503),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1557),
.B(n_1526),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1545),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1543),
.B(n_1503),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1557),
.B(n_1528),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1543),
.B(n_1503),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1557),
.B(n_1556),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1545),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1509),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1556),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1548),
.B(n_1476),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1557),
.B(n_1525),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1576)
);

NOR2xp67_ASAP7_75t_L g1577 ( 
.A(n_1548),
.B(n_1527),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1556),
.B(n_1525),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1545),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1556),
.B(n_1522),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1581)
);

INVxp33_ASAP7_75t_SL g1582 ( 
.A(n_1555),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1538),
.B(n_1499),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1501),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1545),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1540),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1546),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1548),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1548),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1570),
.B(n_1549),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1579),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1570),
.B(n_1532),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1579),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1580),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1586),
.B(n_1554),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1584),
.B(n_1499),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1570),
.B(n_1530),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1580),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1562),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1584),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1583),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1562),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1586),
.B(n_1554),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1582),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1553),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1567),
.A2(n_1558),
.B1(n_1537),
.B2(n_1511),
.Y(n_1612)
);

OAI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1567),
.A2(n_1559),
.B(n_1530),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1578),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1568),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1561),
.B(n_1553),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1577),
.B(n_1586),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1561),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1587),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1592),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1564),
.B(n_1553),
.Y(n_1623)
);

INVxp67_ASAP7_75t_SL g1624 ( 
.A(n_1583),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_SL g1625 ( 
.A(n_1571),
.B(n_1550),
.Y(n_1625)
);

OAI32xp33_ASAP7_75t_L g1626 ( 
.A1(n_1581),
.A2(n_1558),
.A3(n_1530),
.B1(n_1542),
.B2(n_1539),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1593),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1593),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1564),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1573),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1573),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1560),
.B(n_1554),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1555),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1574),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1589),
.B(n_1546),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1581),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1571),
.B(n_1538),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1613),
.B(n_1589),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1610),
.B(n_1604),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1603),
.B(n_1589),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1605),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1600),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1611),
.B(n_1590),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1635),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1619),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1635),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1625),
.A2(n_1558),
.B1(n_1577),
.B2(n_1542),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1615),
.B(n_1590),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1638),
.B(n_1571),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1606),
.B(n_1590),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1608),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1634),
.B(n_1585),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1602),
.Y(n_1657)
);

AND3x2_ASAP7_75t_L g1658 ( 
.A(n_1634),
.B(n_1595),
.C(n_1555),
.Y(n_1658)
);

OAI32xp33_ASAP7_75t_L g1659 ( 
.A1(n_1602),
.A2(n_1539),
.A3(n_1542),
.B1(n_1531),
.B2(n_1591),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1612),
.B(n_1585),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1614),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1618),
.B(n_1560),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1638),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1637),
.B(n_1585),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1616),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1595),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1631),
.B(n_1539),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1626),
.A2(n_1538),
.B(n_1550),
.Y(n_1669)
);

NAND2x1p5_ASAP7_75t_L g1670 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1607),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1632),
.B(n_1572),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1620),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1638),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1655),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1669),
.B(n_1607),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1624),
.Y(n_1677)
);

AOI222xp33_ASAP7_75t_L g1678 ( 
.A1(n_1639),
.A2(n_1626),
.B1(n_1598),
.B2(n_1531),
.C1(n_1559),
.C2(n_1617),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1670),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1652),
.A2(n_1541),
.B1(n_1618),
.B2(n_1531),
.Y(n_1680)
);

OAI211xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1666),
.A2(n_1636),
.B(n_1594),
.C(n_1559),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1659),
.A2(n_1541),
.B(n_1550),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1662),
.B(n_1601),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1643),
.A2(n_1541),
.B1(n_1623),
.B2(n_1521),
.C(n_1529),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1645),
.B(n_1572),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1659),
.A2(n_1645),
.B(n_1650),
.Y(n_1687)
);

AOI311xp33_ASAP7_75t_L g1688 ( 
.A1(n_1660),
.A2(n_1621),
.A3(n_1629),
.B(n_1628),
.C(n_1627),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1665),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1665),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1654),
.B(n_1622),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1572),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1663),
.A2(n_1674),
.B1(n_1533),
.B2(n_1652),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1652),
.A2(n_1574),
.B1(n_1588),
.B2(n_1571),
.C(n_1536),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1657),
.A2(n_1596),
.B(n_1540),
.C(n_1544),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1671),
.B(n_1576),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1644),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1642),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1652),
.A2(n_1574),
.B1(n_1588),
.B2(n_1536),
.C(n_1535),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1671),
.B(n_1576),
.Y(n_1700)
);

OAI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1681),
.A2(n_1651),
.B(n_1656),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1675),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1685),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1689),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1690),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1680),
.A2(n_1647),
.B1(n_1649),
.B2(n_1658),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1676),
.B(n_1670),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1687),
.B(n_1641),
.C(n_1640),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1679),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1697),
.Y(n_1712)
);

AOI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1678),
.A2(n_1649),
.B(n_1647),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1677),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1670),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1679),
.B(n_1653),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1686),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1683),
.B(n_1688),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1692),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1705),
.A2(n_1682),
.B1(n_1684),
.B2(n_1696),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1700),
.Y(n_1721)
);

AOI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1713),
.A2(n_1699),
.B1(n_1693),
.B2(n_1694),
.C(n_1695),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1683),
.Y(n_1723)
);

OAI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1709),
.A2(n_1716),
.B1(n_1708),
.B2(n_1718),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1707),
.A2(n_1695),
.B(n_1667),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1710),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1711),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1707),
.A2(n_1653),
.B(n_1664),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1712),
.B(n_1662),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1717),
.B(n_1718),
.Y(n_1730)
);

NOR4xp25_ASAP7_75t_L g1731 ( 
.A(n_1724),
.B(n_1714),
.C(n_1702),
.D(n_1703),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1730),
.B(n_1715),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1725),
.A2(n_1701),
.B1(n_1708),
.B2(n_1719),
.C(n_1704),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_SL g1734 ( 
.A(n_1722),
.B(n_1706),
.C(n_1646),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1726),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1723),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1721),
.B(n_1646),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1729),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1729),
.B(n_1661),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1727),
.B(n_1720),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1737),
.B(n_1728),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1738),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1732),
.A2(n_1673),
.B(n_1596),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1732),
.B(n_1596),
.Y(n_1744)
);

AO221x1_ASAP7_75t_L g1745 ( 
.A1(n_1736),
.A2(n_1551),
.B1(n_1547),
.B2(n_1588),
.C(n_1540),
.Y(n_1745)
);

NOR4xp25_ASAP7_75t_L g1746 ( 
.A(n_1741),
.B(n_1740),
.C(n_1734),
.D(n_1733),
.Y(n_1746)
);

XNOR2xp5_ASAP7_75t_L g1747 ( 
.A(n_1742),
.B(n_1731),
.Y(n_1747)
);

NAND4xp25_ASAP7_75t_SL g1748 ( 
.A(n_1743),
.B(n_1739),
.C(n_1735),
.D(n_1745),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1744),
.A2(n_1668),
.B1(n_1672),
.B2(n_1470),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1741),
.A2(n_1594),
.B1(n_1536),
.B2(n_1535),
.C(n_1540),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1742),
.Y(n_1751)
);

XNOR2xp5_ASAP7_75t_L g1752 ( 
.A(n_1747),
.B(n_1465),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1751),
.B(n_1594),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1749),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1748),
.B(n_1454),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1750),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1753),
.B(n_1601),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1753),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1754),
.A2(n_1746),
.B1(n_1609),
.B2(n_1565),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1757),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1760),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1756),
.B1(n_1755),
.B2(n_1759),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1758),
.B1(n_1752),
.B2(n_1609),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

AOI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1762),
.A2(n_1633),
.B(n_1563),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1764),
.B(n_1535),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1765),
.A2(n_1633),
.B1(n_1565),
.B2(n_1575),
.Y(n_1767)
);

OAI211xp5_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1517),
.B(n_1549),
.C(n_1569),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1767),
.B(n_1566),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1769),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1536),
.B1(n_1535),
.B2(n_1575),
.C(n_1565),
.Y(n_1771)
);

AOI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1517),
.B(n_1488),
.C(n_1575),
.Y(n_1772)
);


endmodule