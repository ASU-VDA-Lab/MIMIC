module fake_jpeg_25433_n_408 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_408);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_50),
.Y(n_82)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_59),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_77),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_62),
.Y(n_113)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_69),
.Y(n_93)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_75),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_35),
.B(n_1),
.CON(n_73),
.SN(n_73)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_38),
.B1(n_31),
.B2(n_37),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_1),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_81),
.Y(n_107)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_95),
.A2(n_53),
.B1(n_6),
.B2(n_7),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_31),
.B1(n_37),
.B2(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_100),
.A2(n_119),
.B1(n_120),
.B2(n_55),
.Y(n_167)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_34),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_1),
.B(n_2),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_1),
.B(n_2),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_31),
.B1(n_37),
.B2(n_42),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_49),
.B1(n_43),
.B2(n_47),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_62),
.C(n_51),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_62),
.C(n_79),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_48),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_51),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_78),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_72),
.A2(n_29),
.B1(n_40),
.B2(n_18),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_40),
.B1(n_25),
.B2(n_22),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_128),
.B(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_28),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_134),
.B1(n_141),
.B2(n_153),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_131),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_132),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_134)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_135),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_136),
.B(n_139),
.Y(n_185)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_34),
.B(n_33),
.C(n_41),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_140),
.B(n_143),
.C(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_28),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_28),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_24),
.B1(n_33),
.B2(n_41),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_82),
.B(n_28),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_28),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_154),
.Y(n_173)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_144),
.Y(n_187)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_148),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_2),
.B(n_6),
.Y(n_193)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_41),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_41),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_160),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_89),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_98),
.A2(n_33),
.B1(n_6),
.B2(n_7),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_125),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_41),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_125),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_53),
.C(n_56),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_97),
.B1(n_118),
.B2(n_99),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_113),
.B1(n_87),
.B2(n_102),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_109),
.A2(n_61),
.B1(n_58),
.B2(n_7),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_2),
.B(n_10),
.C(n_11),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_172),
.A2(n_15),
.B1(n_187),
.B2(n_186),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_97),
.B1(n_118),
.B2(n_99),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_188),
.B1(n_201),
.B2(n_130),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_190),
.B1(n_192),
.B2(n_204),
.Y(n_210)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_88),
.C(n_6),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_184),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_193),
.B(n_164),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_154),
.C(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_122),
.B1(n_105),
.B2(n_114),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_128),
.A2(n_87),
.B1(n_111),
.B2(n_94),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_111),
.B1(n_113),
.B2(n_102),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_204),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_116),
.B1(n_7),
.B2(n_9),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_116),
.B1(n_10),
.B2(n_11),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_14),
.B(n_15),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_152),
.B1(n_162),
.B2(n_157),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_176),
.A2(n_145),
.B1(n_151),
.B2(n_158),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_213),
.A2(n_238),
.B1(n_197),
.B2(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_221),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_209),
.C(n_170),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_198),
.C(n_171),
.Y(n_256)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_232),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_219),
.B1(n_220),
.B2(n_226),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_165),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_188),
.A2(n_160),
.B1(n_127),
.B2(n_147),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_144),
.B1(n_137),
.B2(n_135),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_222),
.B(n_224),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_182),
.B(n_132),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_223),
.A2(n_235),
.B(n_237),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_185),
.B(n_149),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_225),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_172),
.A2(n_152),
.B1(n_159),
.B2(n_131),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_166),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_228),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_148),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_13),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_230),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_185),
.B(n_13),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_205),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_237),
.B1(n_240),
.B2(n_246),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_14),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_241),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_201),
.A2(n_15),
.B1(n_173),
.B2(n_199),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_173),
.B(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_178),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_244),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_206),
.B(n_195),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_223),
.B1(n_234),
.B2(n_219),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_194),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_191),
.A2(n_206),
.B1(n_190),
.B2(n_194),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_247),
.B(n_256),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_253),
.A2(n_272),
.B(n_276),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_245),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_254),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_198),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_265),
.C(n_247),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_212),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_258),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_210),
.A2(n_228),
.B1(n_221),
.B2(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_270),
.B1(n_223),
.B2(n_217),
.Y(n_283)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_216),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_196),
.C(n_202),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_268),
.C(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_207),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_273),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_207),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_228),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_203),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_203),
.Y(n_273)
);

OAI32xp33_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_205),
.A3(n_227),
.B1(n_210),
.B2(n_211),
.Y(n_275)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_275),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_235),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_289),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_283),
.A2(n_296),
.B1(n_297),
.B2(n_255),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_244),
.C(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_268),
.C(n_271),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_225),
.B1(n_240),
.B2(n_226),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_299),
.B1(n_250),
.B2(n_258),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_222),
.B(n_211),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_230),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_224),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_300),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_260),
.A2(n_262),
.B1(n_248),
.B2(n_269),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_238),
.B1(n_231),
.B2(n_232),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_255),
.A2(n_238),
.B1(n_231),
.B2(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_301),
.B(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_250),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_249),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_306),
.A2(n_282),
.B1(n_287),
.B2(n_299),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_329),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_327),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_251),
.Y(n_310)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_313),
.C(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_256),
.C(n_249),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_316),
.A2(n_301),
.B1(n_286),
.B2(n_285),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_322),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_261),
.B1(n_251),
.B2(n_275),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_SL g335 ( 
.A(n_320),
.B(n_283),
.C(n_291),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_261),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_263),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_324),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_263),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_259),
.C(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_259),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_329),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_294),
.B(n_259),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_340),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_284),
.C(n_302),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_344),
.C(n_322),
.Y(n_352)
);

OAI321xp33_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_343),
.A3(n_317),
.B1(n_295),
.B2(n_292),
.C(n_285),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_296),
.B1(n_293),
.B2(n_283),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_341),
.B1(n_347),
.B2(n_348),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_326),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_339),
.Y(n_354)
);

AO22x1_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_296),
.B1(n_293),
.B2(n_297),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_321),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_279),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_284),
.C(n_291),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_318),
.Y(n_364)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_315),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_345),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_351),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_342),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_314),
.B(n_281),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_353),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_324),
.C(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_361),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_335),
.A2(n_317),
.B(n_312),
.Y(n_356)
);

OAI21x1_ASAP7_75t_SL g376 ( 
.A1(n_356),
.A2(n_358),
.B(n_362),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_319),
.C(n_313),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_332),
.C(n_334),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_360),
.Y(n_369)
);

BUFx12_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

A2O1A1O1Ixp25_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_307),
.B(n_311),
.C(n_318),
.D(n_298),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_330),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_346),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_366),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_342),
.C(n_359),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_333),
.C(n_364),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_374),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_331),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_363),
.A2(n_300),
.B1(n_308),
.B2(n_304),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_298),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_356),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_381),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_365),
.C(n_369),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_373),
.A2(n_351),
.B1(n_350),
.B2(n_357),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_354),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_386),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_383),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_370),
.A2(n_360),
.B(n_362),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_385),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_376),
.A2(n_361),
.B1(n_339),
.B2(n_297),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_361),
.Y(n_386)
);

NAND2x1_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_392),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_369),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_393),
.Y(n_395)
);

OA21x2_ASAP7_75t_SL g392 ( 
.A1(n_380),
.A2(n_288),
.B(n_289),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_367),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_390),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_396),
.A2(n_397),
.B(n_399),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_371),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_297),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_398),
.A2(n_394),
.B(n_387),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_402),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_395),
.A2(n_379),
.B(n_386),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_400),
.B(n_399),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_404),
.A2(n_297),
.B(n_377),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_405),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_403),
.Y(n_408)
);


endmodule