module real_jpeg_7496_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_0),
.A2(n_54),
.B1(n_108),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_1),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_32),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_1),
.A2(n_96),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_1),
.A2(n_248),
.B(n_251),
.C(n_254),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_262),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_1),
.B(n_81),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_1),
.B(n_105),
.C(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_1),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_1),
.B(n_142),
.C(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_1),
.B(n_25),
.Y(n_323)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_78),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_78),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_6),
.Y(n_262)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_7),
.Y(n_250)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_117),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_9),
.A2(n_46),
.B1(n_122),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_122),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_9),
.A2(n_61),
.B1(n_122),
.B2(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_11),
.Y(n_368)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_13),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_366),
.B(n_369),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_205),
.B1(n_364),
.B2(n_365),
.Y(n_15)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_16),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_203),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_180),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_18),
.B(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.C(n_150),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_19),
.A2(n_20),
.B1(n_110),
.B2(n_111),
.Y(n_234)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_50),
.B2(n_68),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_23),
.A2(n_50),
.B(n_69),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B(n_45),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_24),
.A2(n_44),
.B1(n_45),
.B2(n_154),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_24),
.A2(n_44),
.B1(n_45),
.B2(n_154),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_27),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_27),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_27),
.Y(n_148)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_32),
.Y(n_253)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_50),
.A2(n_68),
.B1(n_70),
.B2(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_51),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_53),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_58),
.B(n_223),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_59),
.A2(n_171),
.B1(n_176),
.B2(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_59),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_60),
.A2(n_223),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_60),
.A2(n_223),
.B1(n_259),
.B2(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_61),
.Y(n_274)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_64),
.Y(n_226)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_66),
.Y(n_277)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_81),
.B(n_91),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_81),
.B1(n_101),
.B2(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_76),
.Y(n_286)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_81),
.B(n_162),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_92),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.Y(n_92)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_93),
.B(n_198),
.Y(n_334)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B(n_149),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_115),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_113),
.B(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_115),
.B(n_153),
.C(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_115),
.A2(n_320),
.B1(n_321),
.B2(n_324),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_115),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_115),
.A2(n_153),
.B1(n_213),
.B2(n_324),
.Y(n_347)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_126),
.B1(n_137),
.B2(n_146),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_126),
.B1(n_137),
.B2(n_146),
.Y(n_152)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_126),
.B(n_137),
.Y(n_231)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_133),
.Y(n_306)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_188),
.B(n_193),
.Y(n_187)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_137),
.Y(n_296)
);

AOI22x1_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_144),
.Y(n_137)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_147),
.A2(n_249),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_182),
.B1(n_183),
.B2(n_201),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_150),
.A2(n_151),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_152),
.A2(n_153),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_152),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_152),
.A2(n_212),
.B1(n_228),
.B2(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_152),
.A2(n_212),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_152),
.B(n_184),
.C(n_334),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_153),
.Y(n_213)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_170),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_159),
.A2(n_160),
.B1(n_170),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_159),
.A2(n_160),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_159),
.A2(n_160),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_160),
.B(n_258),
.C(n_295),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_160),
.B(n_316),
.C(n_318),
.Y(n_329)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_168),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_202),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_200),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_217),
.C(n_230),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_184),
.A2(n_200),
.B1(n_230),
.B2(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_184),
.A2(n_200),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_231),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_205),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI211xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_263),
.B(n_358),
.C(n_363),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_235),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_208),
.A2(n_235),
.B(n_359),
.C(n_362),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_232),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_209),
.B(n_232),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.C(n_216),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_214),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_212),
.B(n_284),
.C(n_303),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_228),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_219),
.A2(n_228),
.B1(n_284),
.B2(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_219),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_228),
.A2(n_284),
.B1(n_285),
.B2(n_289),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_236),
.B(n_238),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.C(n_245),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_240),
.B(n_243),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_245),
.B(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_246),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_257),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_247),
.A2(n_257),
.B1(n_258),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_257),
.A2(n_258),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_258),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_279),
.Y(n_280)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_343),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_328),
.B(n_342),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_313),
.B(n_327),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_300),
.B(n_312),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_291),
.B(n_299),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_281),
.B(n_290),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_278),
.B(n_280),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_282),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_322),
.C(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_289),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_298),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_298),
.Y(n_299)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_302),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_311),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_309),
.B2(n_310),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_310),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_326),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_318),
.B1(n_319),
.B2(n_325),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_330),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_338),
.C(n_339),
.Y(n_352)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_353),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_352),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_352),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_351),
.C(n_355),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_353),
.A2(n_360),
.B(n_361),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_356),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_368),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);


endmodule