module real_jpeg_6458_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_0),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_0),
.Y(n_298)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_0),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_0),
.Y(n_349)
);

INVx8_ASAP7_75t_L g448 ( 
.A(n_0),
.Y(n_448)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_1),
.A2(n_50),
.B1(n_101),
.B2(n_234),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_1),
.A2(n_50),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_1),
.A2(n_50),
.B1(n_252),
.B2(n_283),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_2),
.Y(n_145)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g405 ( 
.A(n_2),
.Y(n_405)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_2),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_3),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_4),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_4),
.A2(n_126),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_4),
.A2(n_83),
.B1(n_126),
.B2(n_222),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_5),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_61),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_61),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_6),
.A2(n_61),
.B1(n_378),
.B2(n_381),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_7),
.A2(n_157),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_7),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_7),
.B(n_80),
.C(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_7),
.B(n_106),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_7),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_7),
.B(n_158),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_7),
.B(n_137),
.Y(n_336)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_8),
.Y(n_497)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_11),
.A2(n_67),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_92),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_11),
.A2(n_92),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_12),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_12),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_12),
.A2(n_187),
.B1(n_284),
.B2(n_303),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_12),
.A2(n_137),
.B1(n_284),
.B2(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_12),
.A2(n_57),
.B1(n_201),
.B2(n_284),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_13),
.Y(n_177)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_13),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_14),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_14),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_14),
.A2(n_67),
.B1(n_200),
.B2(n_257),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_14),
.A2(n_200),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_14),
.A2(n_200),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_16),
.A2(n_60),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_16),
.A2(n_222),
.B1(n_237),
.B2(n_270),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_16),
.A2(n_237),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_16),
.A2(n_237),
.B1(n_369),
.B2(n_425),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_17),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_17),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_17),
.A2(n_116),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_17),
.A2(n_91),
.B1(n_116),
.B2(n_193),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_17),
.A2(n_116),
.B1(n_263),
.B2(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_496),
.B(n_498),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_206),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_205),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_147),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_24),
.B(n_147),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_127),
.B2(n_128),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.C(n_93),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_27),
.A2(n_129),
.B1(n_130),
.B2(n_146),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_27),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_27),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_48),
.B1(n_54),
.B2(n_56),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_28),
.A2(n_54),
.B1(n_56),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_28),
.A2(n_236),
.B(n_240),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_28),
.A2(n_38),
.B1(n_236),
.B2(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_29),
.B(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_29),
.A2(n_418),
.B(n_421),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_36),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_38),
.B(n_254),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

OAI32xp33_ASAP7_75t_L g391 ( 
.A1(n_39),
.A2(n_392),
.A3(n_395),
.B1(n_397),
.B2(n_402),
.Y(n_391)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_43),
.Y(n_138)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_43),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_43),
.Y(n_342)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_45),
.Y(n_139)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_46),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_49),
.B(n_55),
.Y(n_197)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_51),
.Y(n_202)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_54),
.A2(n_198),
.B(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_55),
.B(n_199),
.Y(n_240)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_63),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_62),
.A2(n_63),
.B1(n_93),
.B2(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_79),
.B(n_90),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_64),
.A2(n_251),
.B(n_255),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_64),
.A2(n_281),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_64),
.A2(n_255),
.B(n_327),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_64),
.A2(n_326),
.B1(n_429),
.B2(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_65),
.A2(n_153),
.B1(n_158),
.B2(n_159),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_65),
.A2(n_153),
.B1(n_158),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_65),
.A2(n_158),
.B1(n_192),
.B2(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_65),
.B(n_256),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_79),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_68),
.Y(n_257)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_69),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_69),
.Y(n_283)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_70),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_70),
.Y(n_286)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_76),
.Y(n_260)
);

INVx5_ASAP7_75t_SL g330 ( 
.A(n_76),
.Y(n_330)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_79),
.A2(n_281),
.B(n_287),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_79),
.A2(n_287),
.B(n_429),
.Y(n_428)
);

AOI22x1_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_84),
.Y(n_277)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_91),
.Y(n_328)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_112),
.B1(n_119),
.B2(n_120),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_119),
.B1(n_120),
.B2(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_95),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_95),
.A2(n_119),
.B1(n_163),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_95),
.A2(n_119),
.B1(n_368),
.B2(n_424),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_106),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_96)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_97),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_100),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_105),
.Y(n_334)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_105),
.Y(n_394)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_105),
.Y(n_401)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_106),
.A2(n_113),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_106),
.A2(n_161),
.B1(n_373),
.B2(n_453),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_106)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_118),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_119),
.B(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_119),
.A2(n_368),
.B(n_372),
.Y(n_367)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_138),
.Y(n_371)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_169),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_148),
.B(n_151),
.CI(n_169),
.CON(n_208),
.SN(n_208)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_151),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_160),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g356 ( 
.A(n_157),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_158),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_158),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_161),
.A2(n_333),
.B(n_337),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_161),
.B(n_373),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_161),
.A2(n_337),
.B(n_469),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g350 ( 
.A1(n_168),
.A2(n_336),
.A3(n_351),
.B1(n_352),
.B2(n_356),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B(n_196),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_191),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_196),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_171),
.A2(n_191),
.B1(n_214),
.B2(n_438),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_178),
.B(n_181),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_172),
.A2(n_181),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_172),
.A2(n_269),
.B(n_273),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_172),
.A2(n_254),
.B(n_273),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_172),
.A2(n_296),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_173),
.B(n_274),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_173),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_173),
.A2(n_179),
.B1(n_346),
.B2(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_173),
.A2(n_410),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_175),
.Y(n_348)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_177),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g305 ( 
.A(n_177),
.Y(n_305)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_184),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_191),
.Y(n_438)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_202),
.Y(n_396)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_241),
.B(n_495),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_208),
.B(n_209),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_208),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.C(n_218),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_215),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_218),
.B(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_232),
.C(n_235),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_219),
.B(n_436),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_220),
.B(n_225),
.Y(n_463)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_221),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_223),
.Y(n_315)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_226),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g351 ( 
.A(n_228),
.Y(n_351)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_232),
.B(n_235),
.Y(n_436)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_233),
.Y(n_453)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_240),
.Y(n_421)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI311xp33_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_432),
.A3(n_471),
.B1(n_489),
.C1(n_494),
.Y(n_243)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_385),
.B(n_431),
.Y(n_244)
);

AO21x1_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_359),
.B(n_384),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_320),
.B(n_358),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_290),
.B(n_319),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_267),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_249),
.B(n_267),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_258),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_250),
.A2(n_258),
.B1(n_259),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_SL g333 ( 
.A1(n_254),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_254),
.B(n_403),
.Y(n_402)
);

OAI21xp33_ASAP7_75t_SL g418 ( 
.A1(n_254),
.A2(n_402),
.B(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_279),
.C(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_272),
.Y(n_382)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_288),
.B2(n_289),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_311),
.B(n_318),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_300),
.B(n_310),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_299),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_309),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_309),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_306),
.B(n_308),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_308),
.A2(n_345),
.B(n_349),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_316),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_322),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_343),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_332),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_331),
.C(n_343),
.Y(n_360)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx6_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_350),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_360),
.B(n_361),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_366),
.B2(n_383),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_365),
.C(n_383),
.Y(n_386)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_374),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_375),
.C(n_376),
.Y(n_412)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_377),
.Y(n_408)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_386),
.B(n_387),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_415),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_406),
.B2(n_407),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_412),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_412),
.B(n_413),
.C(n_415),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_422),
.B2(n_430),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_423),
.C(n_428),
.Y(n_480)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_428),
.Y(n_422)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_457),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_433),
.A2(n_457),
.B(n_490),
.C(n_493),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_454),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_434),
.B(n_454),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_437),
.C(n_439),
.Y(n_434)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_435),
.B(n_437),
.CI(n_439),
.CON(n_470),
.SN(n_470)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_449),
.C(n_452),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_443),
.Y(n_479)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx8_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_450),
.B1(n_452),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_452),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_470),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_470),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.C(n_464),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_460),
.B1(n_463),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_463),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.C(n_468),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_470),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_491),
.B(n_492),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_481),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_481),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.C(n_480),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_487),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_486),
.Y(n_491)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx13_ASAP7_75t_L g500 ( 
.A(n_497),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);


endmodule