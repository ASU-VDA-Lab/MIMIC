module fake_jpeg_11022_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_28),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_11),
.B(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_20),
.C(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_0),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_1),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_45),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_9),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_98),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_50),
.A3(n_67),
.B1(n_63),
.B2(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_55),
.B1(n_67),
.B2(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_101),
.B1(n_104),
.B2(n_12),
.Y(n_117)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_5),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_22),
.C(n_38),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_9),
.C(n_10),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_3),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_114),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_117),
.B1(n_44),
.B2(n_33),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_110),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_10),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_95),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_116),
.B(n_120),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_100),
.C(n_92),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_14),
.C(n_19),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_32),
.C(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_21),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_111),
.B1(n_116),
.B2(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_126),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_127),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_125),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_132),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_128),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_122),
.Y(n_137)
);


endmodule