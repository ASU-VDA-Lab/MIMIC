module fake_netlist_1_9366_n_1041 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1041);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1041;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_947;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_991;
wire n_843;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g266 ( .A(n_28), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_40), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_196), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_2), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_151), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_134), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_56), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_247), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_87), .B(n_63), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_38), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_114), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_64), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_97), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_197), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_58), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_202), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_109), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_3), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_211), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_172), .Y(n_288) );
INVxp67_ASAP7_75t_L g289 ( .A(n_26), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_36), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_91), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_126), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_16), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_239), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_66), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_156), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_96), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
INVx4_ASAP7_75t_R g299 ( .A(n_68), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_5), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_222), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_248), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_89), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_241), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_73), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_143), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_175), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_117), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_93), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_84), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_131), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_244), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_37), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_171), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_1), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_178), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_111), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_13), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_120), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_169), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_82), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_22), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_261), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_57), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_221), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_76), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_65), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_127), .Y(n_329) );
INVxp33_ASAP7_75t_SL g330 ( .A(n_112), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_179), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_207), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_11), .Y(n_333) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_16), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_260), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_150), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_115), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_149), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_94), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_26), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_245), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_24), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_170), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_9), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_148), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_61), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_176), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_92), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_249), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_259), .Y(n_350) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_168), .B(n_215), .Y(n_351) );
BUFx2_ASAP7_75t_SL g352 ( .A(n_236), .Y(n_352) );
INVxp33_ASAP7_75t_L g353 ( .A(n_98), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_174), .Y(n_354) );
NOR2xp67_ASAP7_75t_L g355 ( .A(n_122), .B(n_141), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_159), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_69), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_152), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_19), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_11), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_234), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_9), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_184), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_79), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_165), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_164), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_17), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_51), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_177), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_95), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_206), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_216), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_238), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_166), .Y(n_374) );
INVx4_ASAP7_75t_R g375 ( .A(n_257), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_100), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_71), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_7), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_23), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_185), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_121), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_83), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_142), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_90), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_124), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_128), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_173), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_72), .B(n_256), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_189), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_183), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_140), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_20), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_180), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_67), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_80), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_217), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_266), .Y(n_397) );
BUFx8_ASAP7_75t_L g398 ( .A(n_308), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_277), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_277), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_376), .B(n_0), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_272), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_392), .B(n_0), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_270), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_327), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_392), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_275), .B(n_1), .Y(n_409) );
AOI22x1_ASAP7_75t_SL g410 ( .A1(n_319), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_290), .B(n_4), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_285), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_395), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_395), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_300), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_316), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_273), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_281), .Y(n_418) );
CKINVDCx6p67_ASAP7_75t_R g419 ( .A(n_279), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_334), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_342), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_272), .Y(n_422) );
OAI22xp5_ASAP7_75t_SL g423 ( .A1(n_289), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_289), .Y(n_424) );
AND2x2_ASAP7_75t_SL g425 ( .A(n_291), .B(n_29), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_353), .B(n_8), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_359), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_424), .B(n_362), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_402), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_426), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_397), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_424), .B(n_353), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_422), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_422), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_403), .B(n_382), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_426), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_397), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_422), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_409), .B(n_411), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_408), .B(n_367), .Y(n_444) );
AND2x6_ASAP7_75t_L g445 ( .A(n_401), .B(n_298), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_422), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_406), .Y(n_447) );
INVx5_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_419), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_406), .B(n_309), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_399), .Y(n_451) );
OR2x6_ASAP7_75t_L g452 ( .A(n_423), .B(n_352), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_399), .B(n_361), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_412), .B(n_293), .Y(n_454) );
NAND2xp33_ASAP7_75t_R g455 ( .A(n_410), .B(n_330), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_419), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_398), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_444), .B(n_425), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_432), .A2(n_425), .B1(n_404), .B2(n_416), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_435), .A2(n_398), .B1(n_420), .B2(n_292), .Y(n_461) );
OR2x6_ASAP7_75t_L g462 ( .A(n_458), .B(n_398), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_444), .A2(n_303), .B1(n_321), .B2(n_284), .Y(n_463) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_428), .B(n_324), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_440), .A2(n_374), .B1(n_380), .B2(n_356), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_454), .A2(n_421), .B1(n_415), .B2(n_427), .C(n_378), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_449), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_429), .B(n_418), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_443), .B(n_439), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_433), .B(n_417), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_443), .B(n_333), .C(n_323), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_457), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_439), .B(n_417), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_433), .B(n_337), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_441), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_441), .B(n_337), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_452), .A2(n_340), .B1(n_360), .B2(n_344), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_456), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_447), .B(n_341), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_448), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_452), .B(n_379), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_450), .B(n_341), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_448), .B(n_349), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_450), .B(n_329), .Y(n_484) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_448), .B(n_349), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_451), .A2(n_400), .B(n_407), .C(n_405), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_456), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_445), .B(n_282), .Y(n_489) );
AO22x1_ASAP7_75t_L g490 ( .A1(n_445), .A2(n_329), .B1(n_455), .B2(n_286), .Y(n_490) );
NOR2xp33_ASAP7_75t_R g491 ( .A(n_455), .B(n_288), .Y(n_491) );
NOR2xp67_ASAP7_75t_L g492 ( .A(n_451), .B(n_413), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_445), .B(n_294), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_445), .B(n_297), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_453), .B(n_413), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_453), .B(n_268), .C(n_267), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_469), .A2(n_414), .B(n_271), .C(n_274), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_474), .A2(n_278), .B(n_269), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_468), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_459), .A2(n_283), .B1(n_287), .B2(n_280), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_470), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_460), .A2(n_296), .B1(n_304), .B2(n_302), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_462), .A2(n_306), .B1(n_312), .B2(n_305), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_489), .A2(n_494), .B(n_493), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_472), .B(n_295), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_485), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_485), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_487), .A2(n_320), .B(n_314), .Y(n_509) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_466), .A2(n_307), .B(n_301), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_462), .A2(n_328), .B1(n_335), .B2(n_325), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_462), .A2(n_339), .B1(n_343), .B2(n_338), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_481), .A2(n_354), .B(n_357), .C(n_348), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_467), .B(n_313), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_484), .B(n_315), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_484), .B(n_317), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_464), .B(n_298), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_463), .A2(n_365), .B1(n_366), .B2(n_364), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_465), .B(n_10), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_461), .B(n_311), .Y(n_520) );
BUFx4f_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_473), .B(n_318), .Y(n_522) );
OAI21xp33_ASAP7_75t_SL g523 ( .A1(n_476), .A2(n_369), .B(n_368), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_477), .B(n_10), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_497), .Y(n_525) );
BUFx8_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_471), .B(n_331), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_478), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_483), .A2(n_384), .B(n_385), .C(n_370), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_491), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_475), .A2(n_372), .B(n_371), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_479), .B(n_322), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_SL g533 ( .A1(n_482), .A2(n_276), .B(n_442), .C(n_438), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_478), .B(n_326), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_496), .B(n_332), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_486), .A2(n_390), .B1(n_377), .B2(n_383), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_490), .B(n_480), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_492), .B(n_336), .Y(n_539) );
NOR2xp67_ASAP7_75t_R g540 ( .A(n_462), .B(n_386), .Y(n_540) );
OAI22x1_ASAP7_75t_L g541 ( .A1(n_517), .A2(n_504), .B1(n_512), .B2(n_519), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_505), .A2(n_391), .B(n_389), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_521), .B(n_345), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_521), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_509), .A2(n_396), .B(n_393), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_533), .A2(n_387), .B(n_430), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_526), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_536), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_501), .B(n_346), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_511), .A2(n_345), .B1(n_394), .B2(n_350), .Y(n_550) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_507), .A2(n_355), .B(n_351), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_498), .A2(n_363), .B(n_276), .C(n_388), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_513), .B(n_347), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_520), .B(n_358), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_524), .B(n_12), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_530), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_525), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_525), .B(n_373), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_500), .A2(n_446), .B(n_437), .C(n_436), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_526), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_507), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_502), .B(n_381), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_503), .B(n_12), .Y(n_563) );
BUFx4_ASAP7_75t_SL g564 ( .A(n_540), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_518), .B(n_13), .Y(n_565) );
NAND2x1_ASAP7_75t_L g566 ( .A(n_508), .B(n_299), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_523), .B(n_14), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_528), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
CKINVDCx8_ASAP7_75t_R g571 ( .A(n_538), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_527), .Y(n_572) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_508), .A2(n_431), .B(n_430), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_529), .B(n_310), .C(n_272), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_506), .B(n_14), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_532), .A2(n_437), .B(n_434), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_499), .A2(n_310), .B(n_272), .C(n_431), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_515), .B(n_516), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_534), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_537), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_531), .B(n_15), .Y(n_581) );
NOR4xp25_ASAP7_75t_L g582 ( .A(n_510), .B(n_15), .C(n_17), .D(n_18), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_522), .B(n_18), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_514), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_539), .A2(n_436), .B(n_434), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_535), .B(n_19), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_517), .B(n_20), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_588), .A2(n_310), .B(n_375), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_580), .B(n_21), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_555), .B(n_23), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_544), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_548), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_542), .A2(n_310), .B(n_31), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_547), .Y(n_595) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_573), .A2(n_32), .B(n_30), .Y(n_596) );
AO31x2_ASAP7_75t_L g597 ( .A1(n_546), .A2(n_24), .A3(n_25), .B(n_27), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_567), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_557), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_541), .B(n_25), .Y(n_600) );
NOR2xp67_ASAP7_75t_L g601 ( .A(n_560), .B(n_27), .Y(n_601) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_545), .A2(n_586), .B(n_576), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_565), .Y(n_603) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_551), .A2(n_146), .B(n_33), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_579), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_581), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_544), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_569), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_572), .B(n_28), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_544), .B(n_265), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_554), .B(n_34), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_557), .Y(n_612) );
AOI21x1_ASAP7_75t_L g613 ( .A1(n_574), .A2(n_35), .B(n_39), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_575), .B(n_264), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_563), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_571), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_557), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_584), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_587), .Y(n_619) );
AO31x2_ASAP7_75t_L g620 ( .A1(n_577), .A2(n_47), .A3(n_48), .B(n_49), .Y(n_620) );
OAI21x1_ASAP7_75t_L g621 ( .A1(n_566), .A2(n_50), .B(n_52), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_559), .A2(n_53), .B(n_54), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_584), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_583), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_584), .Y(n_625) );
OA21x2_ASAP7_75t_L g626 ( .A1(n_574), .A2(n_55), .B(n_59), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_585), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_568), .B(n_60), .Y(n_628) );
CKINVDCx6p67_ASAP7_75t_R g629 ( .A(n_564), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_553), .B(n_62), .Y(n_630) );
AOI21xp33_ASAP7_75t_SL g631 ( .A1(n_556), .A2(n_70), .B(n_74), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_562), .B(n_75), .Y(n_632) );
INVx6_ASAP7_75t_L g633 ( .A(n_558), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_552), .A2(n_77), .B(n_78), .C(n_81), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_570), .Y(n_635) );
AO31x2_ASAP7_75t_L g636 ( .A1(n_582), .A2(n_85), .A3(n_86), .B(n_88), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_550), .B(n_549), .Y(n_637) );
INVx6_ASAP7_75t_L g638 ( .A(n_558), .Y(n_638) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_543), .A2(n_99), .B(n_101), .Y(n_639) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_561), .A2(n_102), .B(n_103), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_580), .B(n_104), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_558), .B(n_105), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_580), .B(n_106), .Y(n_643) );
NOR2x1_ASAP7_75t_SL g644 ( .A(n_557), .B(n_107), .Y(n_644) );
OAI21x1_ASAP7_75t_SL g645 ( .A1(n_567), .A2(n_108), .B(n_110), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_580), .B(n_113), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_548), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_578), .A2(n_116), .B(n_118), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_578), .A2(n_119), .B(n_123), .Y(n_649) );
INVx3_ASAP7_75t_L g650 ( .A(n_544), .Y(n_650) );
BUFx8_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_625), .Y(n_652) );
OA21x2_ASAP7_75t_L g653 ( .A1(n_602), .A2(n_125), .B(n_129), .Y(n_653) );
AOI21xp5_ASAP7_75t_SL g654 ( .A1(n_616), .A2(n_130), .B(n_132), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_633), .Y(n_655) );
BUFx3_ASAP7_75t_L g656 ( .A(n_651), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_647), .B(n_263), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_596), .A2(n_622), .B(n_640), .Y(n_658) );
BUFx3_ASAP7_75t_L g659 ( .A(n_651), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_593), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_605), .Y(n_661) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_625), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_625), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_590), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_600), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_633), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_608), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_608), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_627), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_606), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_591), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_599), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_609), .B(n_133), .Y(n_673) );
AO21x2_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_135), .B(n_136), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_603), .B(n_262), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_612), .B(n_137), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_597), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_604), .Y(n_678) );
AO21x2_ASAP7_75t_L g679 ( .A1(n_641), .A2(n_138), .B(n_139), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_597), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_601), .B(n_144), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_595), .B(n_145), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_604), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_597), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_617), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_618), .Y(n_686) );
AO21x2_ASAP7_75t_L g687 ( .A1(n_643), .A2(n_147), .B(n_153), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_598), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_619), .B(n_154), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_624), .B(n_155), .Y(n_690) );
AO21x2_ASAP7_75t_L g691 ( .A1(n_646), .A2(n_157), .B(n_158), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_628), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_628), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_638), .Y(n_694) );
OAI21x1_ASAP7_75t_L g695 ( .A1(n_613), .A2(n_160), .B(n_161), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_589), .B(n_258), .Y(n_696) );
BUFx2_ASAP7_75t_SL g697 ( .A(n_629), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_637), .B(n_162), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_638), .Y(n_699) );
AO21x2_ASAP7_75t_L g700 ( .A1(n_634), .A2(n_163), .B(n_167), .Y(n_700) );
BUFx3_ASAP7_75t_L g701 ( .A(n_607), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_607), .B(n_181), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_592), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_623), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_592), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_650), .Y(n_706) );
INVx3_ASAP7_75t_L g707 ( .A(n_650), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_635), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_611), .B(n_630), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_639), .Y(n_710) );
OR2x6_ASAP7_75t_L g711 ( .A(n_610), .B(n_182), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_635), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_621), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_635), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_636), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_632), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_636), .Y(n_717) );
NOR2x1_ASAP7_75t_SL g718 ( .A(n_642), .B(n_186), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_614), .B(n_187), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_615), .Y(n_720) );
INVx2_ASAP7_75t_SL g721 ( .A(n_620), .Y(n_721) );
NOR2x1p5_ASAP7_75t_L g722 ( .A(n_631), .B(n_188), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_644), .B(n_191), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_620), .Y(n_724) );
BUFx2_ASAP7_75t_R g725 ( .A(n_644), .Y(n_725) );
AOI21x1_ASAP7_75t_L g726 ( .A1(n_626), .A2(n_254), .B(n_194), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_648), .B(n_193), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_649), .A2(n_195), .B1(n_198), .B2(n_199), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_620), .B(n_253), .Y(n_729) );
AOI33xp33_ASAP7_75t_L g730 ( .A1(n_594), .A2(n_200), .A3(n_203), .B1(n_204), .B2(n_205), .B3(n_208), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_626), .Y(n_731) );
INVxp67_ASAP7_75t_SL g732 ( .A(n_625), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_593), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_633), .Y(n_734) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_625), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_591), .B(n_209), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_605), .B(n_210), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_591), .B(n_212), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_605), .B(n_213), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_605), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_606), .B(n_214), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_605), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_665), .B(n_218), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_661), .B(n_252), .Y(n_744) );
BUFx2_ASAP7_75t_L g745 ( .A(n_701), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_671), .B(n_219), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_740), .B(n_250), .Y(n_747) );
AND2x4_ASAP7_75t_SL g748 ( .A(n_711), .B(n_220), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_664), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_742), .B(n_673), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_667), .B(n_226), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_660), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_733), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_663), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_733), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_663), .Y(n_756) );
INVx2_ASAP7_75t_SL g757 ( .A(n_701), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_669), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_688), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_672), .Y(n_760) );
AO21x2_ASAP7_75t_L g761 ( .A1(n_713), .A2(n_227), .B(n_228), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_734), .B(n_229), .Y(n_762) );
INVx5_ASAP7_75t_L g763 ( .A(n_656), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_668), .Y(n_764) );
INVx4_ASAP7_75t_L g765 ( .A(n_711), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_655), .B(n_230), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_670), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_668), .B(n_231), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_677), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_736), .B(n_738), .Y(n_770) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_672), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_704), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_694), .B(n_232), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_699), .B(n_233), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_656), .Y(n_775) );
OR2x2_ASAP7_75t_L g776 ( .A(n_704), .B(n_235), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_692), .B(n_246), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_680), .Y(n_778) );
BUFx3_ASAP7_75t_L g779 ( .A(n_659), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_684), .B(n_237), .Y(n_780) );
INVx4_ASAP7_75t_L g781 ( .A(n_711), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_678), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_678), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_662), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_693), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_657), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_685), .B(n_240), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_683), .Y(n_788) );
AO21x2_ASAP7_75t_L g789 ( .A1(n_683), .A2(n_242), .B(n_243), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_666), .B(n_682), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_685), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_666), .B(n_659), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_706), .B(n_698), .Y(n_793) );
INVx5_ASAP7_75t_L g794 ( .A(n_662), .Y(n_794) );
INVx5_ASAP7_75t_L g795 ( .A(n_662), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_689), .B(n_690), .Y(n_796) );
OR2x2_ASAP7_75t_L g797 ( .A(n_703), .B(n_686), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_686), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_708), .B(n_652), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_708), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_741), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_652), .B(n_732), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_741), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_732), .Y(n_804) );
BUFx3_ASAP7_75t_L g805 ( .A(n_662), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_681), .B(n_702), .Y(n_806) );
AND2x4_ASAP7_75t_L g807 ( .A(n_712), .B(n_714), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_716), .B(n_709), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_712), .B(n_735), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_741), .Y(n_810) );
INVx5_ASAP7_75t_L g811 ( .A(n_735), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_735), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_735), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_737), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_739), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_705), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_731), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_723), .B(n_729), .Y(n_818) );
NOR2x1_ASAP7_75t_SL g819 ( .A(n_697), .B(n_696), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_705), .B(n_707), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_731), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_707), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_675), .B(n_676), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_720), .B(n_676), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_724), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_725), .Y(n_826) );
INVx2_ASAP7_75t_SL g827 ( .A(n_676), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_723), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_715), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_719), .B(n_727), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_719), .B(n_723), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_717), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_722), .B(n_730), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_710), .B(n_721), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_760), .B(n_674), .Y(n_835) );
INVx3_ASAP7_75t_L g836 ( .A(n_765), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_759), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_750), .B(n_691), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_745), .B(n_691), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_757), .B(n_687), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_771), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_752), .B(n_730), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_757), .B(n_687), .Y(n_843) );
AND2x4_ASAP7_75t_SL g844 ( .A(n_765), .B(n_728), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_790), .B(n_679), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_758), .Y(n_846) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_804), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_804), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_765), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_770), .B(n_679), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_753), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_755), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_793), .B(n_653), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_767), .B(n_700), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_772), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_792), .B(n_658), .Y(n_856) );
AND2x4_ASAP7_75t_L g857 ( .A(n_781), .B(n_718), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_806), .B(n_728), .Y(n_858) );
OR2x2_ASAP7_75t_L g859 ( .A(n_764), .B(n_654), .Y(n_859) );
AND2x4_ASAP7_75t_SL g860 ( .A(n_781), .B(n_754), .Y(n_860) );
BUFx2_ASAP7_75t_L g861 ( .A(n_779), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_781), .B(n_695), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_754), .Y(n_863) );
INVx3_ASAP7_75t_L g864 ( .A(n_794), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_756), .B(n_726), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_756), .B(n_808), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_797), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_800), .B(n_786), .Y(n_868) );
OR2x2_ASAP7_75t_L g869 ( .A(n_799), .B(n_802), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_800), .B(n_785), .Y(n_870) );
INVx4_ASAP7_75t_L g871 ( .A(n_763), .Y(n_871) );
OR2x2_ASAP7_75t_L g872 ( .A(n_791), .B(n_798), .Y(n_872) );
NOR2x1_ASAP7_75t_L g873 ( .A(n_779), .B(n_775), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_820), .B(n_831), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_769), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_807), .B(n_796), .Y(n_876) );
AND2x4_ASAP7_75t_L g877 ( .A(n_828), .B(n_763), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_807), .B(n_823), .Y(n_878) );
OR2x2_ASAP7_75t_L g879 ( .A(n_826), .B(n_824), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_829), .Y(n_880) );
INVx6_ASAP7_75t_L g881 ( .A(n_763), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_801), .B(n_810), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_778), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_816), .Y(n_884) );
BUFx2_ASAP7_75t_L g885 ( .A(n_763), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_803), .B(n_807), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_822), .B(n_768), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_776), .Y(n_888) );
NAND2x1_ASAP7_75t_L g889 ( .A(n_827), .B(n_834), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_814), .B(n_815), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_751), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_780), .Y(n_892) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_782), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_830), .B(n_780), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_827), .B(n_818), .Y(n_895) );
INVx1_ASAP7_75t_SL g896 ( .A(n_805), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_819), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_746), .B(n_809), .Y(n_898) );
OR2x2_ASAP7_75t_L g899 ( .A(n_818), .B(n_829), .Y(n_899) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_832), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_832), .B(n_813), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_809), .B(n_787), .Y(n_902) );
NOR2xp67_ASAP7_75t_L g903 ( .A(n_871), .B(n_795), .Y(n_903) );
NAND2x1_ASAP7_75t_L g904 ( .A(n_881), .B(n_834), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_837), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_846), .Y(n_906) );
AND3x1_ASAP7_75t_L g907 ( .A(n_873), .B(n_833), .C(n_743), .Y(n_907) );
INVx2_ASAP7_75t_SL g908 ( .A(n_861), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_869), .B(n_788), .Y(n_909) );
NAND2x1p5_ASAP7_75t_L g910 ( .A(n_871), .B(n_795), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_876), .B(n_809), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_874), .B(n_834), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_866), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_855), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_878), .B(n_813), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_867), .B(n_812), .Y(n_916) );
CKINVDCx16_ASAP7_75t_R g917 ( .A(n_879), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_894), .B(n_812), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_870), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_870), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_847), .B(n_788), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_868), .B(n_812), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_902), .B(n_784), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_856), .B(n_784), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_847), .Y(n_925) );
AND3x1_ASAP7_75t_L g926 ( .A(n_836), .B(n_743), .C(n_762), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_841), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_841), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_884), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_851), .B(n_821), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_852), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_872), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_890), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_863), .B(n_821), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_848), .Y(n_935) );
NAND2x1p5_ASAP7_75t_L g936 ( .A(n_885), .B(n_794), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_863), .B(n_817), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_850), .B(n_783), .Y(n_938) );
NAND2xp5_ASAP7_75t_SL g939 ( .A(n_862), .B(n_748), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_890), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_897), .B(n_836), .Y(n_941) );
AND2x4_ASAP7_75t_L g942 ( .A(n_860), .B(n_825), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_858), .A2(n_748), .B1(n_773), .B2(n_774), .Y(n_943) );
NAND2xp5_ASAP7_75t_SL g944 ( .A(n_862), .B(n_795), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_848), .Y(n_945) );
BUFx3_ASAP7_75t_L g946 ( .A(n_881), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_880), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_898), .B(n_784), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_882), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_838), .B(n_825), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_882), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_875), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_935), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_919), .B(n_845), .Y(n_954) );
OR2x2_ASAP7_75t_L g955 ( .A(n_909), .B(n_899), .Y(n_955) );
NAND2x1p5_ASAP7_75t_L g956 ( .A(n_903), .B(n_864), .Y(n_956) );
NAND2x1_ASAP7_75t_L g957 ( .A(n_908), .B(n_881), .Y(n_957) );
NAND4xp25_ASAP7_75t_L g958 ( .A(n_943), .B(n_849), .C(n_853), .D(n_895), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_920), .B(n_888), .Y(n_959) );
AOI21xp33_ASAP7_75t_SL g960 ( .A1(n_939), .A2(n_849), .B(n_857), .Y(n_960) );
OR2x6_ASAP7_75t_L g961 ( .A(n_939), .B(n_857), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_921), .Y(n_962) );
NAND2xp33_ASAP7_75t_SL g963 ( .A(n_904), .B(n_889), .Y(n_963) );
NOR5xp2_ASAP7_75t_L g964 ( .A(n_935), .B(n_900), .C(n_880), .D(n_893), .E(n_883), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_927), .B(n_839), .C(n_835), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_947), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_933), .B(n_900), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_905), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_917), .A2(n_864), .B1(n_892), .B2(n_896), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_912), .B(n_860), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_906), .Y(n_971) );
OR2x2_ASAP7_75t_L g972 ( .A(n_913), .B(n_893), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_925), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_911), .B(n_896), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_945), .Y(n_975) );
O2A1O1Ixp33_ASAP7_75t_L g976 ( .A1(n_940), .A2(n_842), .B(n_747), .C(n_744), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_934), .Y(n_977) );
OR2x2_ASAP7_75t_L g978 ( .A(n_938), .B(n_886), .Y(n_978) );
NAND2x1p5_ASAP7_75t_L g979 ( .A(n_946), .B(n_811), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_949), .B(n_886), .Y(n_980) );
INVxp67_ASAP7_75t_L g981 ( .A(n_941), .Y(n_981) );
AOI21xp33_ASAP7_75t_L g982 ( .A1(n_976), .A2(n_941), .B(n_928), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_967), .Y(n_983) );
INVx3_ASAP7_75t_L g984 ( .A(n_957), .Y(n_984) );
INVx1_ASAP7_75t_SL g985 ( .A(n_974), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_975), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_978), .B(n_938), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_956), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_975), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_977), .B(n_951), .Y(n_990) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_964), .B(n_907), .C(n_914), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g992 ( .A1(n_958), .A2(n_926), .B1(n_918), .B2(n_915), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_977), .Y(n_993) );
NAND2xp5_ASAP7_75t_SL g994 ( .A(n_963), .B(n_936), .Y(n_994) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_961), .A2(n_936), .B1(n_944), .B2(n_910), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_969), .A2(n_932), .B1(n_929), .B2(n_931), .C(n_950), .Y(n_996) );
OAI21xp5_ASAP7_75t_L g997 ( .A1(n_981), .A2(n_944), .B(n_910), .Y(n_997) );
OR2x2_ASAP7_75t_L g998 ( .A(n_955), .B(n_950), .Y(n_998) );
A2O1A1Ixp33_ASAP7_75t_L g999 ( .A1(n_960), .A2(n_844), .B(n_970), .C(n_965), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_986), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_996), .B(n_953), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g1002 ( .A1(n_992), .A2(n_961), .B1(n_954), .B2(n_980), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_999), .A2(n_995), .B1(n_988), .B2(n_994), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1004 ( .A1(n_982), .A2(n_959), .B1(n_968), .B2(n_971), .C(n_953), .Y(n_1004) );
NAND2xp5_ASAP7_75t_SL g1005 ( .A(n_984), .B(n_979), .Y(n_1005) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_991), .A2(n_962), .B1(n_973), .B2(n_966), .C(n_972), .Y(n_1006) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_988), .Y(n_1007) );
AOI211xp5_ASAP7_75t_L g1008 ( .A1(n_997), .A2(n_877), .B(n_948), .C(n_922), .Y(n_1008) );
NOR3xp33_ASAP7_75t_L g1009 ( .A(n_984), .B(n_766), .C(n_777), .Y(n_1009) );
AOI322xp5_ASAP7_75t_L g1010 ( .A1(n_985), .A2(n_983), .A3(n_993), .B1(n_990), .B2(n_989), .C1(n_923), .C2(n_924), .Y(n_1010) );
O2A1O1Ixp5_ASAP7_75t_L g1011 ( .A1(n_987), .A2(n_937), .B(n_934), .C(n_952), .Y(n_1011) );
NOR3xp33_ASAP7_75t_L g1012 ( .A(n_998), .B(n_842), .C(n_937), .Y(n_1012) );
NAND3xp33_ASAP7_75t_SL g1013 ( .A(n_994), .B(n_749), .C(n_859), .Y(n_1013) );
OAI21xp33_ASAP7_75t_SL g1014 ( .A1(n_994), .A2(n_930), .B(n_840), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_982), .A2(n_916), .B1(n_930), .B2(n_887), .C(n_844), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_982), .A2(n_891), .B1(n_843), .B2(n_865), .C(n_942), .Y(n_1016) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_994), .A2(n_942), .B(n_877), .Y(n_1017) );
NAND3xp33_ASAP7_75t_L g1018 ( .A(n_991), .B(n_749), .C(n_854), .Y(n_1018) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_1003), .A2(n_1004), .B1(n_1006), .B2(n_1001), .C(n_1007), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1000), .Y(n_1020) );
INVxp33_ASAP7_75t_L g1021 ( .A(n_1005), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1011), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1012), .Y(n_1023) );
NOR2x1_ASAP7_75t_L g1024 ( .A(n_1023), .B(n_1013), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_1022), .Y(n_1025) );
NOR3xp33_ASAP7_75t_L g1026 ( .A(n_1019), .B(n_1014), .C(n_1018), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1020), .B(n_1010), .Y(n_1027) );
AND3x4_ASAP7_75t_L g1028 ( .A(n_1026), .B(n_1009), .C(n_1021), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1025), .Y(n_1029) );
NAND4xp25_ASAP7_75t_L g1030 ( .A(n_1024), .B(n_1002), .C(n_1015), .D(n_1008), .Y(n_1030) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_1029), .B(n_1027), .C(n_1016), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1028), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1030), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1033), .Y(n_1034) );
NOR2xp67_ASAP7_75t_L g1035 ( .A(n_1032), .B(n_1017), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_1035), .A2(n_1031), .B1(n_761), .B2(n_811), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1034), .Y(n_1037) );
XOR2x2_ASAP7_75t_L g1038 ( .A(n_1037), .B(n_1036), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_1038), .A2(n_805), .B1(n_811), .B2(n_795), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_1039), .A2(n_811), .B1(n_794), .B2(n_901), .Y(n_1040) );
AOI21xp33_ASAP7_75t_L g1041 ( .A1(n_1040), .A2(n_789), .B(n_794), .Y(n_1041) );
endmodule