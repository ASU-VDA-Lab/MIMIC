module fake_netlist_6_4641_n_1615 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1615);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1615;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_20),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_29),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_59),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_61),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_84),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_3),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_35),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_56),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_15),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_43),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_116),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_98),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_95),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_91),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_13),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_9),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_60),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_25),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_11),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_11),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_65),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_29),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_24),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_58),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_66),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_19),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_111),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_8),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_25),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_37),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_108),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_83),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_6),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_38),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_105),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_64),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_12),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_54),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_41),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_146),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_143),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_77),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_10),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_89),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_50),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_90),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_21),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_145),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_86),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_41),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_87),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_28),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_68),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_28),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_80),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_30),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_26),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_121),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_99),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_48),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_96),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_46),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_100),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_26),
.Y(n_250)
);

INVxp33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_63),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_43),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_0),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_48),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_85),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_92),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_33),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_107),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_31),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_37),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_70),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_6),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_94),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_31),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_30),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_49),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_24),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_101),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_22),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_103),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_136),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_18),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_15),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_82),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_140),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_34),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_13),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_46),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_23),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_40),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_45),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_88),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_19),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_159),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_235),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_192),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_194),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_174),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_153),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_193),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_252),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_167),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_188),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_194),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_200),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_194),
.Y(n_311)
);

BUFx6f_ASAP7_75t_SL g312 ( 
.A(n_238),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_194),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_209),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_194),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_225),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_196),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_151),
.Y(n_322)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_233),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_262),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_149),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_220),
.B(n_163),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_157),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_296),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_197),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_271),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_151),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_199),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_201),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_162),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_205),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_207),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_208),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_160),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_161),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_195),
.B(n_3),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_177),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_214),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_179),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_212),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_153),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_217),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_219),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_221),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_223),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_226),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_228),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_230),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_227),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_232),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_162),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_239),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_242),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_245),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_248),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_158),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_189),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_254),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_263),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_191),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_273),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_152),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_323),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_148),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_299),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_301),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_305),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_152),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_321),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_309),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_344),
.B(n_238),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_R g385 ( 
.A(n_365),
.B(n_154),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_172),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_335),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_368),
.B(n_154),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_337),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_338),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_333),
.B(n_172),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_331),
.B(n_183),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_175),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g413 ( 
.A(n_307),
.B(n_195),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_347),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_303),
.B(n_236),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_346),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_347),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_308),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_355),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_341),
.A2(n_283),
.B(n_281),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_325),
.B(n_155),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_327),
.B(n_155),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_352),
.B(n_156),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_356),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_175),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_323),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_415),
.B(n_358),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_430),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_392),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_430),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_415),
.B(n_359),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_306),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_390),
.B(n_313),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_376),
.B(n_334),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_376),
.B(n_185),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_390),
.B(n_185),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_413),
.B(n_255),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_413),
.B(n_340),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_407),
.B(n_186),
.Y(n_460)
);

BUFx6f_ASAP7_75t_SL g461 ( 
.A(n_386),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_186),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_383),
.A2(n_187),
.B1(n_293),
.B2(n_287),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_255),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_379),
.B(n_300),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_383),
.B(n_278),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_373),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_413),
.B(n_278),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_382),
.B(n_286),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_379),
.B(n_229),
.Y(n_471)
);

BUFx4f_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_380),
.B(n_381),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_373),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_382),
.A2(n_187),
.B1(n_290),
.B2(n_292),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_374),
.B(n_353),
.Y(n_481)
);

NAND2x1p5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_150),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_385),
.B(n_370),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_392),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_385),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_400),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_408),
.B(n_270),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g492 ( 
.A(n_420),
.B(n_218),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_441),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_384),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_387),
.B(n_286),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_372),
.B(n_169),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_375),
.B(n_329),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_441),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_400),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_441),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_411),
.A2(n_362),
.B(n_361),
.Y(n_510)
);

AND3x2_ASAP7_75t_L g511 ( 
.A(n_420),
.B(n_267),
.C(n_184),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_411),
.B(n_181),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_386),
.B(n_238),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_425),
.B(n_310),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_382),
.A2(n_297),
.B1(n_190),
.B2(n_279),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_382),
.B(n_183),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_393),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_382),
.A2(n_190),
.B1(n_279),
.B2(n_222),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_382),
.A2(n_190),
.B1(n_279),
.B2(n_222),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_411),
.B(n_362),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_393),
.B(n_206),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_403),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_393),
.B(n_210),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_382),
.A2(n_279),
.B1(n_215),
.B2(n_190),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_409),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_377),
.B(n_312),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_403),
.B(n_216),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_429),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_410),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_399),
.B(n_401),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_391),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_394),
.B(n_363),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_431),
.B(n_240),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_391),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_437),
.A2(n_269),
.B1(n_266),
.B2(n_289),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_431),
.B(n_363),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_397),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_432),
.A2(n_295),
.B1(n_158),
.B2(n_257),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_410),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_404),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_436),
.B(n_244),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_391),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_436),
.A2(n_198),
.B1(n_298),
.B2(n_237),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_386),
.B(n_156),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_410),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_386),
.B(n_164),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_395),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_396),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_396),
.B(n_366),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_402),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_402),
.B(n_369),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_391),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_405),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_405),
.B(n_246),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_391),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_397),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_398),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_398),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_391),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_398),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_412),
.B(n_414),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_412),
.B(n_249),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_386),
.B(n_164),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_414),
.B(n_261),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_416),
.B(n_165),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_423),
.B(n_369),
.Y(n_579)
);

AND2x2_ASAP7_75t_SL g580 ( 
.A(n_423),
.B(n_183),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_424),
.B(n_367),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_424),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_427),
.B(n_268),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_458),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_L g585 ( 
.A(n_538),
.B(n_422),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_458),
.A2(n_190),
.B1(n_222),
.B2(n_215),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_539),
.B(n_371),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_453),
.B(n_428),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_539),
.B(n_371),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_467),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

AND2x6_ASAP7_75t_SL g592 ( 
.A(n_505),
.B(n_251),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_458),
.A2(n_442),
.B1(n_438),
.B2(n_316),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_498),
.B(n_442),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_498),
.B(n_406),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_539),
.B(n_183),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

AND2x2_ASAP7_75t_SL g598 ( 
.A(n_580),
.B(n_215),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_500),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_466),
.A2(n_247),
.B1(n_170),
.B2(n_291),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_580),
.B(n_215),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_506),
.B(n_417),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_509),
.B(n_417),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_539),
.B(n_222),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_554),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_445),
.B(n_165),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_544),
.A2(n_318),
.B1(n_328),
.B2(n_324),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_451),
.B(n_427),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_580),
.B(n_418),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

NAND2x1_ASAP7_75t_L g612 ( 
.A(n_542),
.B(n_410),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_454),
.B(n_418),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_500),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_561),
.B(n_419),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_545),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_561),
.B(n_419),
.Y(n_617)
);

AOI22x1_ASAP7_75t_L g618 ( 
.A1(n_535),
.A2(n_439),
.B1(n_435),
.B2(n_434),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_566),
.B(n_419),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_568),
.B(n_166),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_566),
.B(n_421),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_559),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_549),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_582),
.B(n_421),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_568),
.B(n_168),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_582),
.B(n_464),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_565),
.A2(n_426),
.B(n_421),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_536),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_563),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_472),
.B(n_173),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_451),
.B(n_426),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_545),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_452),
.B(n_426),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_452),
.B(n_517),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_529),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_565),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_544),
.B(n_176),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_574),
.B(n_433),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_488),
.B(n_367),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_574),
.B(n_433),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_531),
.B(n_434),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_541),
.B(n_176),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_461),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_472),
.B(n_180),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_472),
.B(n_180),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_551),
.B(n_224),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_523),
.B(n_224),
.Y(n_651)
);

OAI221xp5_ASAP7_75t_L g652 ( 
.A1(n_463),
.A2(n_202),
.B1(n_234),
.B2(n_231),
.C(n_213),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_459),
.B(n_203),
.C(n_204),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_540),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_507),
.B(n_425),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_544),
.A2(n_259),
.B1(n_243),
.B2(n_253),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_534),
.A2(n_272),
.B1(n_170),
.B2(n_291),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_502),
.B(n_243),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_544),
.A2(n_265),
.B1(n_259),
.B2(n_285),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_572),
.B(n_258),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_471),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_502),
.B(n_265),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_502),
.B(n_534),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_488),
.B(n_162),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_534),
.B(n_285),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_450),
.B(n_312),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_521),
.B(n_410),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_522),
.B(n_410),
.Y(n_668)
);

OAI221xp5_ASAP7_75t_L g669 ( 
.A1(n_510),
.A2(n_546),
.B1(n_457),
.B2(n_460),
.C(n_462),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_528),
.B(n_410),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_312),
.Y(n_671)
);

AOI221xp5_ASAP7_75t_L g672 ( 
.A1(n_546),
.A2(n_288),
.B1(n_282),
.B2(n_280),
.C(n_277),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_535),
.B(n_211),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_523),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_564),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_447),
.B(n_470),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_490),
.B(n_275),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_492),
.B(n_507),
.C(n_486),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_549),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_578),
.B(n_553),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_570),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_478),
.A2(n_275),
.B1(n_274),
.B2(n_272),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_579),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_490),
.B(n_264),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_579),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_523),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_470),
.B(n_260),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_474),
.B(n_260),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_581),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_443),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_555),
.B(n_257),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_474),
.B(n_256),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_489),
.B(n_256),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_581),
.Y(n_695)
);

OAI221xp5_ASAP7_75t_L g696 ( 
.A1(n_510),
.A2(n_250),
.B1(n_247),
.B2(n_182),
.C(n_178),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_489),
.B(n_250),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_562),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_443),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_558),
.A2(n_576),
.B1(n_512),
.B2(n_469),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_471),
.B(n_182),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_518),
.B(n_178),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_171),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_518),
.B(n_171),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_495),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_562),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_491),
.B(n_4),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_461),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_491),
.B(n_4),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_482),
.B(n_147),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_481),
.B(n_8),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_465),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_482),
.A2(n_134),
.B1(n_132),
.B2(n_131),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_518),
.B(n_126),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_518),
.B(n_117),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_543),
.B(n_10),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_503),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_476),
.B(n_12),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_461),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_515),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_482),
.B(n_109),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_547),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_492),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_567),
.B(n_14),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_599),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_613),
.A2(n_496),
.B(n_446),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_586),
.B(n_537),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_586),
.B(n_469),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_722),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_633),
.B(n_469),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_674),
.A2(n_469),
.B(n_525),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_597),
.B(n_537),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_674),
.A2(n_469),
.B(n_525),
.Y(n_733)
);

OAI321xp33_ASAP7_75t_L g734 ( 
.A1(n_657),
.A2(n_543),
.A3(n_465),
.B1(n_575),
.B2(n_583),
.C(n_577),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_628),
.A2(n_449),
.B(n_479),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_608),
.B(n_477),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_L g737 ( 
.A1(n_701),
.A2(n_501),
.B(n_515),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_SL g738 ( 
.A(n_672),
.B(n_511),
.C(n_533),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_584),
.B(n_519),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_636),
.B(n_469),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_614),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_681),
.A2(n_560),
.B(n_557),
.C(n_548),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_661),
.B(n_588),
.Y(n_743)
);

OR2x6_ASAP7_75t_SL g744 ( 
.A(n_720),
.B(n_504),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_665),
.A2(n_513),
.B(n_508),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_598),
.B(n_560),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_597),
.B(n_537),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_687),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_701),
.B(n_557),
.Y(n_749)
);

OAI21xp33_ASAP7_75t_L g750 ( 
.A1(n_707),
.A2(n_548),
.B(n_524),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_597),
.B(n_556),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_588),
.B(n_449),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_640),
.A2(n_479),
.B(n_532),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_681),
.A2(n_573),
.B(n_571),
.C(n_526),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_700),
.A2(n_547),
.B1(n_556),
.B2(n_571),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_669),
.A2(n_473),
.B(n_475),
.C(n_480),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_640),
.A2(n_485),
.B(n_530),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_601),
.B(n_493),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_723),
.B(n_594),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_639),
.A2(n_547),
.B1(n_448),
.B2(n_456),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_595),
.A2(n_485),
.B(n_530),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_677),
.B(n_493),
.Y(n_762)
);

AO21x1_ASAP7_75t_L g763 ( 
.A1(n_710),
.A2(n_473),
.B(n_475),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_717),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_638),
.B(n_456),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_602),
.A2(n_485),
.B(n_530),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_712),
.B(n_448),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_642),
.B(n_493),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_644),
.B(n_654),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_678),
.B(n_480),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_603),
.A2(n_530),
.B(n_520),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_707),
.A2(n_497),
.B(n_494),
.C(n_487),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_685),
.B(n_448),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_665),
.A2(n_494),
.B(n_497),
.C(n_499),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_620),
.A2(n_516),
.B(n_499),
.C(n_487),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_721),
.A2(n_520),
.B(n_444),
.Y(n_776)
);

AO21x1_ASAP7_75t_L g777 ( 
.A1(n_721),
.A2(n_14),
.B(n_16),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_698),
.B(n_483),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_610),
.A2(n_520),
.B(n_444),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_L g780 ( 
.A(n_692),
.B(n_516),
.C(n_484),
.Y(n_780)
);

AOI31xp33_ASAP7_75t_L g781 ( 
.A1(n_657),
.A2(n_16),
.A3(n_17),
.B(n_22),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_609),
.A2(n_547),
.B1(n_484),
.B2(n_483),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_611),
.A2(n_527),
.B(n_455),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_716),
.A2(n_718),
.B1(n_724),
.B2(n_709),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_632),
.A2(n_527),
.B(n_455),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_647),
.B(n_27),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_632),
.A2(n_527),
.B(n_455),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_718),
.A2(n_527),
.B(n_455),
.C(n_36),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_606),
.A2(n_81),
.B1(n_79),
.B2(n_78),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_687),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_648),
.A2(n_74),
.B(n_73),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_606),
.B(n_32),
.C(n_34),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_624),
.B(n_72),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_676),
.B(n_32),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_623),
.B(n_71),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_616),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_684),
.B(n_38),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_686),
.B(n_39),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_649),
.A2(n_55),
.B(n_40),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_722),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_660),
.A2(n_39),
.B(n_42),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_616),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_635),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_649),
.A2(n_658),
.B(n_662),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_690),
.B(n_44),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_675),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_724),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_53),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_596),
.A2(n_54),
.B(n_604),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_615),
.A2(n_625),
.B(n_621),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_646),
.B(n_650),
.Y(n_811)
);

CKINVDCx8_ASAP7_75t_R g812 ( 
.A(n_592),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_617),
.A2(n_619),
.B(n_587),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_706),
.B(n_630),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_627),
.A2(n_722),
.B(n_629),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_591),
.B(n_605),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_589),
.A2(n_631),
.B1(n_634),
.B2(n_626),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_692),
.A2(n_679),
.B1(n_653),
.B2(n_641),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_664),
.B(n_705),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_643),
.B(n_711),
.Y(n_820)
);

INVx11_ASAP7_75t_L g821 ( 
.A(n_680),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_722),
.B(n_593),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_622),
.B(n_645),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_641),
.A2(n_643),
.B1(n_656),
.B2(n_659),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_618),
.A2(n_704),
.B(n_702),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_655),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_688),
.B(n_689),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_693),
.B(n_694),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_697),
.B(n_673),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_714),
.A2(n_715),
.B(n_612),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_590),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_682),
.A2(n_699),
.B(n_691),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_651),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_667),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_668),
.A2(n_670),
.B(n_713),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_703),
.A2(n_666),
.B(n_671),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_600),
.B(n_607),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_647),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_643),
.B(n_683),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_652),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_696),
.A2(n_647),
.B(n_708),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_719),
.B(n_708),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_719),
.B(n_708),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_719),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_655),
.B(n_584),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_584),
.B(n_661),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_586),
.A2(n_681),
.B(n_709),
.C(n_707),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_586),
.B(n_539),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_681),
.A2(n_584),
.B1(n_458),
.B2(n_669),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_669),
.A2(n_584),
.B(n_637),
.C(n_468),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_586),
.B(n_539),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_643),
.Y(n_857)
);

AOI22x1_ASAP7_75t_SL g858 ( 
.A1(n_720),
.A2(n_425),
.B1(n_373),
.B2(n_266),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_586),
.B(n_539),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_586),
.B(n_550),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_586),
.A2(n_681),
.B(n_709),
.C(n_707),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_SL g863 ( 
.A(n_609),
.B(n_539),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_669),
.A2(n_584),
.B(n_637),
.C(n_468),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_599),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_608),
.B(n_451),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_584),
.B(n_661),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_663),
.A2(n_568),
.B(n_552),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_802),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_848),
.A2(n_861),
.B(n_854),
.Y(n_871)
);

INVx4_ASAP7_75t_SL g872 ( 
.A(n_838),
.Y(n_872)
);

OAI21x1_ASAP7_75t_SL g873 ( 
.A1(n_777),
.A2(n_799),
.B(n_791),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_848),
.A2(n_861),
.B1(n_784),
.B2(n_860),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_800),
.B(n_863),
.Y(n_875)
);

AO31x2_ASAP7_75t_L g876 ( 
.A1(n_742),
.A2(n_772),
.A3(n_763),
.B(n_754),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_866),
.B(n_846),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_846),
.B(n_868),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_725),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_736),
.B(n_819),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_784),
.A2(n_849),
.B1(n_807),
.B2(n_727),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_857),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_741),
.Y(n_883)
);

OA21x2_ASAP7_75t_L g884 ( 
.A1(n_742),
.A2(n_745),
.B(n_772),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_838),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_868),
.B(n_811),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_856),
.A2(n_859),
.B(n_727),
.Y(n_887)
);

OAI22xp33_ASAP7_75t_L g888 ( 
.A1(n_818),
.A2(n_781),
.B1(n_734),
.B2(n_839),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_833),
.B(n_838),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_827),
.B(n_828),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_855),
.A2(n_864),
.B(n_835),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_749),
.B(n_759),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_761),
.A2(n_771),
.B(n_766),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_743),
.B(n_820),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_752),
.B(n_770),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_849),
.A2(n_850),
.B(n_847),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_851),
.A2(n_853),
.B(n_852),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_840),
.A2(n_836),
.B(n_743),
.C(n_845),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_800),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_769),
.B(n_829),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_862),
.A2(n_869),
.B(n_867),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_845),
.B(n_773),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_754),
.A2(n_740),
.B(n_730),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_824),
.B(n_737),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_810),
.A2(n_813),
.B(n_735),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_814),
.A2(n_807),
.B(n_831),
.Y(n_906)
);

AO22x1_ASAP7_75t_L g907 ( 
.A1(n_814),
.A2(n_841),
.B1(n_826),
.B2(n_748),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_728),
.A2(n_746),
.B1(n_797),
.B2(n_794),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_739),
.A2(n_733),
.B(n_731),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_823),
.B(n_748),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_796),
.Y(n_911)
);

AO31x2_ASAP7_75t_L g912 ( 
.A1(n_788),
.A2(n_739),
.A3(n_817),
.B(n_760),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_773),
.B(n_765),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_834),
.A2(n_825),
.B(n_755),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_732),
.A2(n_747),
.B(n_751),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_753),
.A2(n_726),
.B(n_762),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_768),
.A2(n_779),
.B(n_782),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_738),
.A2(n_798),
.B(n_805),
.C(n_808),
.Y(n_918)
);

AO21x1_ASAP7_75t_L g919 ( 
.A1(n_795),
.A2(n_822),
.B(n_780),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_858),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_834),
.B(n_778),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_756),
.A2(n_758),
.B(n_788),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_774),
.A2(n_775),
.B(n_750),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_792),
.A2(n_837),
.B1(n_806),
.B2(n_789),
.Y(n_924)
);

BUFx8_ASAP7_75t_L g925 ( 
.A(n_838),
.Y(n_925)
);

AO21x2_ASAP7_75t_L g926 ( 
.A1(n_795),
.A2(n_757),
.B(n_776),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_778),
.B(n_865),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_844),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_729),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_803),
.Y(n_930)
);

OAI21x1_ASAP7_75t_L g931 ( 
.A1(n_785),
.A2(n_787),
.B(n_783),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_744),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_764),
.A2(n_816),
.B(n_765),
.Y(n_933)
);

CKINVDCx11_ASAP7_75t_R g934 ( 
.A(n_812),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_767),
.B(n_790),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_809),
.A2(n_767),
.B(n_801),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_729),
.A2(n_842),
.B(n_843),
.Y(n_937)
);

NOR2x1_ASAP7_75t_SL g938 ( 
.A(n_844),
.B(n_786),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_793),
.A2(n_786),
.B(n_821),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_786),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_866),
.B(n_846),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_725),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_848),
.A2(n_861),
.B(n_734),
.C(n_781),
.Y(n_943)
);

AO31x2_ASAP7_75t_L g944 ( 
.A1(n_742),
.A2(n_772),
.A3(n_763),
.B(n_848),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_866),
.B(n_846),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_848),
.A2(n_681),
.B(n_861),
.C(n_854),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_848),
.A2(n_861),
.B(n_854),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_725),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_845),
.A2(n_681),
.B1(n_588),
.B2(n_453),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_800),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_848),
.A2(n_681),
.B(n_861),
.C(n_854),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_856),
.A2(n_568),
.B(n_552),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_866),
.B(n_854),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_848),
.A2(n_861),
.B(n_854),
.Y(n_954)
);

AO31x2_ASAP7_75t_L g955 ( 
.A1(n_742),
.A2(n_772),
.A3(n_763),
.B(n_848),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_848),
.A2(n_681),
.B(n_861),
.C(n_854),
.Y(n_956)
);

NOR2x1_ASAP7_75t_L g957 ( 
.A(n_842),
.B(n_585),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_833),
.B(n_687),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_800),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_866),
.B(n_846),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_832),
.A2(n_830),
.B(n_815),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_866),
.B(n_854),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_866),
.B(n_846),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_848),
.A2(n_681),
.B(n_861),
.C(n_854),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_848),
.A2(n_681),
.B(n_861),
.C(n_854),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_866),
.B(n_846),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_854),
.A2(n_586),
.B1(n_861),
.B2(n_848),
.Y(n_967)
);

NAND2x1_ASAP7_75t_L g968 ( 
.A(n_800),
.B(n_597),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_866),
.B(n_854),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_854),
.A2(n_586),
.B1(n_861),
.B2(n_848),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_736),
.B(n_467),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_814),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_831),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_866),
.B(n_854),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_800),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_736),
.B(n_866),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_866),
.B(n_854),
.Y(n_977)
);

OAI21x1_ASAP7_75t_SL g978 ( 
.A1(n_777),
.A2(n_799),
.B(n_791),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_736),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_725),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_848),
.A2(n_861),
.B(n_854),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_866),
.B(n_846),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_838),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_736),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_725),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_725),
.Y(n_986)
);

AO21x1_ASAP7_75t_L g987 ( 
.A1(n_856),
.A2(n_859),
.B(n_804),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_866),
.B(n_854),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_870),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_973),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_878),
.B(n_949),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_879),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_905),
.A2(n_887),
.B(n_952),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_886),
.A2(n_890),
.B1(n_892),
.B2(n_895),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_883),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_886),
.B(n_890),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_942),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_885),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_880),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_979),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_889),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_877),
.B(n_941),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_948),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_899),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_885),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_894),
.B(n_892),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_945),
.B(n_960),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_939),
.B(n_885),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_963),
.B(n_966),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_971),
.B(n_984),
.Y(n_1010)
);

CKINVDCx6p67_ASAP7_75t_R g1011 ( 
.A(n_934),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_943),
.A2(n_946),
.B(n_951),
.C(n_956),
.Y(n_1012)
);

INVx3_ASAP7_75t_SL g1013 ( 
.A(n_872),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_976),
.B(n_972),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_983),
.B(n_940),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_982),
.B(n_888),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_925),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_906),
.B(n_958),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_958),
.B(n_882),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_904),
.B(n_900),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_925),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_953),
.B(n_962),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_967),
.A2(n_970),
.B1(n_981),
.B2(n_871),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_924),
.A2(n_964),
.B(n_965),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_L g1025 ( 
.A(n_983),
.B(n_918),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_911),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_975),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_921),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_889),
.B(n_920),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_924),
.A2(n_977),
.B1(n_974),
.B2(n_969),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_928),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_932),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_953),
.B(n_962),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_967),
.A2(n_970),
.B(n_981),
.C(n_947),
.Y(n_1034)
);

BUFx10_ASAP7_75t_L g1035 ( 
.A(n_983),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_940),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_872),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_881),
.A2(n_902),
.B1(n_898),
.B2(n_974),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_975),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_969),
.B(n_988),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_929),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_930),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_891),
.A2(n_916),
.B(n_901),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_897),
.A2(n_917),
.B(n_896),
.Y(n_1044)
);

CKINVDCx8_ASAP7_75t_R g1045 ( 
.A(n_872),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_910),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_881),
.B(n_921),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_980),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_975),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_985),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_986),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_907),
.B(n_933),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_874),
.A2(n_871),
.B(n_947),
.C(n_954),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_908),
.A2(n_909),
.B(n_914),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_938),
.B(n_957),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_913),
.A2(n_874),
.B1(n_954),
.B2(n_927),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_935),
.B(n_929),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_975),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_908),
.B(n_927),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_919),
.B(n_987),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_922),
.B(n_914),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_937),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_922),
.B(n_912),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_899),
.B(n_959),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_912),
.B(n_903),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_875),
.A2(n_959),
.B1(n_950),
.B2(n_923),
.Y(n_1066)
);

BUFx4f_ASAP7_75t_SL g1067 ( 
.A(n_968),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_873),
.A2(n_978),
.B(n_936),
.C(n_923),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_936),
.A2(n_903),
.B1(n_926),
.B2(n_915),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_875),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_926),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_944),
.B(n_955),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_876),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_876),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_944),
.B(n_884),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_961),
.A2(n_893),
.B(n_931),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_934),
.Y(n_1077)
);

CKINVDCx6p67_ASAP7_75t_R g1078 ( 
.A(n_934),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_894),
.B(n_880),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_973),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_943),
.A2(n_586),
.B(n_951),
.C(n_946),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_973),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_889),
.B(n_872),
.Y(n_1083)
);

INVx3_ASAP7_75t_SL g1084 ( 
.A(n_971),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_949),
.A2(n_886),
.B1(n_784),
.B2(n_890),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_925),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_975),
.B(n_899),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_870),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_886),
.B(n_890),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_889),
.B(n_872),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_973),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_973),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_681),
.B(n_943),
.C(n_861),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_885),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_943),
.A2(n_586),
.B(n_951),
.C(n_946),
.Y(n_1095)
);

CKINVDCx8_ASAP7_75t_R g1096 ( 
.A(n_872),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_878),
.B(n_949),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_979),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_943),
.A2(n_586),
.B(n_951),
.C(n_946),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_886),
.B(n_890),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_899),
.Y(n_1101)
);

OA22x2_ASAP7_75t_L g1102 ( 
.A1(n_949),
.A2(n_543),
.B1(n_716),
.B2(n_546),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_973),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_888),
.A2(n_781),
.B1(n_784),
.B2(n_943),
.C(n_967),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_L g1105 ( 
.A(n_886),
.B(n_586),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_889),
.B(n_872),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_894),
.B(n_880),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_949),
.A2(n_886),
.B1(n_784),
.B2(n_890),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_925),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_886),
.B(n_890),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_879),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_973),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_894),
.B(n_880),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_1011),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1048),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1104),
.A2(n_1016),
.B1(n_1102),
.B2(n_1024),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1020),
.B(n_1016),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_991),
.B(n_1097),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_992),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1093),
.A2(n_1097),
.B(n_991),
.Y(n_1120)
);

INVxp33_ASAP7_75t_L g1121 ( 
.A(n_1010),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_995),
.Y(n_1122)
);

CKINVDCx6p67_ASAP7_75t_R g1123 ( 
.A(n_1078),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_997),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1018),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1003),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1035),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1077),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1008),
.B(n_1083),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_1089),
.B1(n_1110),
.B2(n_1100),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_990),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1102),
.A2(n_1006),
.B1(n_1007),
.B2(n_1032),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1091),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1017),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1073),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1039),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1104),
.A2(n_1023),
.B1(n_1108),
.B2(n_1085),
.Y(n_1137)
);

CKINVDCx6p67_ASAP7_75t_R g1138 ( 
.A(n_1013),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1103),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1039),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1074),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1088),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_1021),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1112),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1072),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1007),
.B(n_1002),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1023),
.A2(n_1084),
.B1(n_1006),
.B2(n_1040),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1013),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1072),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1031),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_1084),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1022),
.B(n_1030),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1075),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1009),
.B(n_1079),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1000),
.Y(n_1155)
);

BUFx2_ASAP7_75t_R g1156 ( 
.A(n_1086),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1107),
.B(n_1113),
.Y(n_1157)
);

INVx6_ASAP7_75t_L g1158 ( 
.A(n_1039),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1008),
.B(n_1083),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1050),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1051),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1049),
.B(n_1040),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1111),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1000),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1098),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1081),
.A2(n_1095),
.B1(n_1099),
.B2(n_999),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1081),
.A2(n_1095),
.B1(n_1099),
.B2(n_999),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1014),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1109),
.Y(n_1169)
);

CKINVDCx6p67_ASAP7_75t_R g1170 ( 
.A(n_1058),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1026),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1098),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_994),
.B(n_1033),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1042),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1057),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_1043),
.A2(n_1076),
.B(n_1044),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1028),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1063),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1065),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1012),
.B(n_1034),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1025),
.A2(n_1061),
.B1(n_1038),
.B2(n_1054),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1105),
.A2(n_1052),
.B1(n_1056),
.B2(n_1046),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1068),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1035),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1034),
.A2(n_1012),
.B1(n_1028),
.B2(n_1082),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1047),
.A2(n_1019),
.B1(n_1029),
.B2(n_1055),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1036),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1044),
.A2(n_993),
.B(n_1060),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1049),
.B(n_1060),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1053),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1071),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1008),
.B(n_1090),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1053),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1082),
.A2(n_1055),
.B1(n_1080),
.B2(n_1092),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1059),
.A2(n_1066),
.B1(n_1069),
.B2(n_1070),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1070),
.A2(n_1015),
.B1(n_1067),
.B2(n_1041),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1062),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1004),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1045),
.A2(n_1096),
.B1(n_1015),
.B2(n_1067),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1027),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1062),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1015),
.Y(n_1202)
);

OAI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1058),
.A2(n_1037),
.B1(n_1087),
.B2(n_1106),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1004),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1064),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1101),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1001),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1106),
.B(n_1101),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_998),
.B(n_1094),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1087),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1005),
.A2(n_949),
.B1(n_1089),
.B2(n_996),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1005),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_998),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_998),
.A2(n_1104),
.B1(n_888),
.B2(n_1016),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_998),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1094),
.B(n_1020),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1094),
.A2(n_588),
.B1(n_949),
.B2(n_308),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1035),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_996),
.A2(n_949),
.B1(n_1100),
.B2(n_1089),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_989),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_SL g1221 ( 
.A1(n_991),
.A2(n_588),
.B1(n_743),
.B2(n_425),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_990),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1102),
.A2(n_588),
.B1(n_824),
.B2(n_991),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_990),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1104),
.A2(n_888),
.B1(n_1016),
.B2(n_1102),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1135),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1135),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1155),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1141),
.Y(n_1229)
);

BUFx2_ASAP7_75t_SL g1230 ( 
.A(n_1187),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1173),
.B(n_1118),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1118),
.B(n_1117),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1197),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1201),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1201),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1155),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1165),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1133),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1165),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1173),
.B(n_1152),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1179),
.B(n_1178),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1172),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1183),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1114),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1117),
.B(n_1120),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1153),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1191),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1125),
.B(n_1152),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1221),
.B(n_1157),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1180),
.B(n_1125),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1177),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1145),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1145),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1149),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1180),
.B(n_1216),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1188),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1176),
.A2(n_1193),
.B(n_1190),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1172),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1185),
.B(n_1166),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1195),
.A2(n_1181),
.B(n_1137),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1219),
.B(n_1146),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1164),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1216),
.B(n_1116),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1189),
.A2(n_1162),
.B(n_1190),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1167),
.B(n_1182),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1200),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1175),
.B(n_1225),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1189),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1162),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1144),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1132),
.B(n_1205),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1119),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1122),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1124),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1211),
.A2(n_1161),
.B(n_1126),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1224),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1160),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1163),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1130),
.B(n_1147),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1223),
.B(n_1214),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1154),
.B(n_1168),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1203),
.Y(n_1283)
);

AO21x1_ASAP7_75t_SL g1284 ( 
.A1(n_1202),
.A2(n_1186),
.B(n_1215),
.Y(n_1284)
);

INVx4_ASAP7_75t_SL g1285 ( 
.A(n_1158),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1158),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1158),
.B(n_1140),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1258),
.B(n_1227),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1249),
.B(n_1121),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1270),
.B(n_1192),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1260),
.A2(n_1217),
.B1(n_1194),
.B2(n_1187),
.Y(n_1291)
);

AOI33xp33_ASAP7_75t_R g1292 ( 
.A1(n_1271),
.A2(n_1151),
.A3(n_1222),
.B1(n_1139),
.B2(n_1131),
.B3(n_1156),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1249),
.B(n_1115),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1258),
.B(n_1220),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1270),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1258),
.B(n_1229),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1265),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1270),
.B(n_1159),
.Y(n_1298)
);

OAI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1266),
.A2(n_1196),
.B1(n_1199),
.B2(n_1150),
.C(n_1171),
.Y(n_1299)
);

INVx6_ASAP7_75t_L g1300 ( 
.A(n_1285),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1276),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1276),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1240),
.B(n_1150),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1258),
.B(n_1220),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1276),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_L g1307 ( 
.A(n_1262),
.B(n_1210),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1260),
.A2(n_1174),
.B(n_1142),
.Y(n_1308)
);

INVxp33_ASAP7_75t_L g1309 ( 
.A(n_1282),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1262),
.B(n_1198),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1283),
.Y(n_1311)
);

INVx3_ASAP7_75t_SL g1312 ( 
.A(n_1285),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1283),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1283),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1240),
.B(n_1198),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1276),
.B(n_1204),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1231),
.B(n_1204),
.Y(n_1317)
);

AOI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1281),
.A2(n_1192),
.B1(n_1159),
.B2(n_1129),
.C(n_1143),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1281),
.A2(n_1159),
.B1(n_1129),
.B2(n_1192),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1231),
.B(n_1206),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1246),
.B(n_1206),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1257),
.B(n_1213),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1246),
.B(n_1213),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1228),
.B(n_1129),
.Y(n_1324)
);

AOI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1280),
.A2(n_1143),
.B1(n_1169),
.B2(n_1208),
.C(n_1148),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1257),
.B(n_1209),
.Y(n_1326)
);

AOI322xp5_ASAP7_75t_L g1327 ( 
.A1(n_1250),
.A2(n_1169),
.A3(n_1114),
.B1(n_1134),
.B2(n_1212),
.C1(n_1128),
.C2(n_1184),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1236),
.B(n_1170),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1269),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1266),
.A2(n_1261),
.B1(n_1280),
.B2(n_1272),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1291),
.A2(n_1272),
.B(n_1268),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1326),
.B(n_1251),
.Y(n_1332)
);

OAI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1330),
.A2(n_1268),
.B(n_1264),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1309),
.B(n_1289),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1289),
.B(n_1237),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1323),
.B(n_1242),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1323),
.B(n_1263),
.Y(n_1337)
);

OA211x2_ASAP7_75t_L g1338 ( 
.A1(n_1292),
.A2(n_1238),
.B(n_1285),
.C(n_1284),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1291),
.A2(n_1261),
.B1(n_1282),
.B2(n_1230),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1303),
.B(n_1277),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1325),
.A2(n_1261),
.B1(n_1264),
.B2(n_1230),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1292),
.A2(n_1232),
.B1(n_1239),
.B2(n_1259),
.C(n_1256),
.Y(n_1342)
);

OAI221xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1327),
.A2(n_1232),
.B1(n_1138),
.B2(n_1123),
.C(n_1256),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1321),
.B(n_1259),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1325),
.B(n_1286),
.Y(n_1345)
);

OAI221xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1327),
.A2(n_1318),
.B1(n_1299),
.B2(n_1319),
.C(n_1328),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1321),
.B(n_1315),
.Y(n_1347)
);

NAND4xp25_ASAP7_75t_L g1348 ( 
.A(n_1299),
.B(n_1279),
.C(n_1273),
.D(n_1274),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1311),
.B(n_1255),
.Y(n_1349)
);

OAI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1318),
.A2(n_1261),
.B1(n_1286),
.B2(n_1269),
.C(n_1184),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1311),
.B(n_1233),
.Y(n_1351)
);

AOI221xp5_ASAP7_75t_L g1352 ( 
.A1(n_1310),
.A2(n_1274),
.B1(n_1273),
.B2(n_1278),
.C(n_1279),
.Y(n_1352)
);

OAI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1328),
.A2(n_1308),
.B1(n_1307),
.B2(n_1310),
.C(n_1320),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1315),
.B(n_1267),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1320),
.B(n_1317),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1293),
.B(n_1324),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_SL g1357 ( 
.A(n_1312),
.B(n_1287),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1312),
.A2(n_1212),
.B1(n_1138),
.B2(n_1287),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1313),
.B(n_1233),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1307),
.A2(n_1269),
.B(n_1208),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1301),
.B(n_1278),
.C(n_1243),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1313),
.B(n_1234),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1314),
.B(n_1234),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1324),
.B(n_1244),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1293),
.B(n_1275),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1290),
.A2(n_1284),
.B1(n_1269),
.B2(n_1123),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1306),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1322),
.B(n_1235),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1300),
.A2(n_1245),
.B1(n_1241),
.B2(n_1247),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1301),
.B(n_1252),
.C(n_1248),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1322),
.B(n_1253),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1322),
.B(n_1253),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1290),
.B(n_1285),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1329),
.B(n_1254),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1367),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1347),
.B(n_1288),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1367),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1332),
.B(n_1288),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1371),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1355),
.B(n_1288),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1371),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1353),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1332),
.B(n_1296),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1374),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1372),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1356),
.B(n_1316),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1361),
.A2(n_1305),
.B(n_1302),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1334),
.B(n_1316),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1349),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1372),
.B(n_1297),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1368),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1336),
.B(n_1296),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1337),
.B(n_1294),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1349),
.Y(n_1394)
);

NOR2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1348),
.B(n_1170),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1351),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1354),
.B(n_1294),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1359),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1340),
.B(n_1295),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1362),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1363),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1335),
.B(n_1128),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1333),
.A2(n_1298),
.B1(n_1290),
.B2(n_1300),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1377),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1377),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1382),
.B(n_1352),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1390),
.B(n_1297),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1398),
.B(n_1364),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1390),
.B(n_1297),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1375),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1390),
.B(n_1297),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1390),
.B(n_1297),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1375),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1375),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1379),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1379),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1382),
.B(n_1331),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1381),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1396),
.Y(n_1420)
);

NOR3xp33_ASAP7_75t_L g1421 ( 
.A(n_1387),
.B(n_1331),
.C(n_1346),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1388),
.B(n_1344),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1387),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1381),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1398),
.B(n_1290),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1390),
.B(n_1297),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1385),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_1297),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1384),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1403),
.B(n_1361),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1385),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1391),
.Y(n_1432)
);

NOR2x1_ASAP7_75t_L g1433 ( 
.A(n_1395),
.B(n_1370),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1391),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1384),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1403),
.B(n_1370),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1376),
.B(n_1304),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1396),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1376),
.B(n_1304),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1418),
.B(n_1402),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1407),
.B(n_1392),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1405),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1430),
.B(n_1388),
.Y(n_1444)
);

AOI32xp33_ASAP7_75t_L g1445 ( 
.A1(n_1421),
.A2(n_1339),
.A3(n_1333),
.B1(n_1398),
.B2(n_1404),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1406),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1425),
.B(n_1398),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1421),
.B(n_1339),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1407),
.B(n_1392),
.Y(n_1449)
);

NAND2x1p5_ASAP7_75t_L g1450 ( 
.A(n_1433),
.B(n_1395),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1425),
.B(n_1389),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1428),
.B(n_1408),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1433),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1428),
.B(n_1389),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1416),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1409),
.B(n_1134),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1409),
.A2(n_1338),
.B1(n_1357),
.B2(n_1345),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_R g1459 ( 
.A(n_1408),
.B(n_1410),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1423),
.B(n_1380),
.Y(n_1460)
);

AO21x1_ASAP7_75t_L g1461 ( 
.A1(n_1423),
.A2(n_1360),
.B(n_1369),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1414),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1435),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1422),
.B(n_1380),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1416),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1417),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1417),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1422),
.B(n_1397),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1414),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1429),
.A2(n_1343),
.B(n_1348),
.C(n_1350),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1428),
.B(n_1408),
.Y(n_1471)
);

NAND2x1_ASAP7_75t_L g1472 ( 
.A(n_1435),
.B(n_1400),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1430),
.B(n_1397),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1436),
.B(n_1399),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1410),
.A2(n_1338),
.B1(n_1357),
.B2(n_1358),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1419),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1410),
.B(n_1383),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1436),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1419),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1437),
.B(n_1393),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1414),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1437),
.B(n_1393),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1442),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1450),
.Y(n_1484)
);

XNOR2xp5_ASAP7_75t_L g1485 ( 
.A(n_1448),
.B(n_1341),
.Y(n_1485)
);

OR2x6_ASAP7_75t_L g1486 ( 
.A(n_1450),
.B(n_1148),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1472),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1453),
.B(n_1412),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1443),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1446),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1440),
.B(n_1386),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1450),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1454),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1448),
.A2(n_1366),
.B1(n_1360),
.B2(n_1429),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1457),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1472),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1463),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1444),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1456),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1444),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1465),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1441),
.B(n_1424),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1449),
.B(n_1424),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1478),
.B(n_1427),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1466),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1470),
.A2(n_1300),
.B1(n_1394),
.B2(n_1342),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1467),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1460),
.B(n_1420),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1476),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1455),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1462),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1455),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1451),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1471),
.B(n_1413),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1487),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1483),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1485),
.B(n_1445),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1484),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1485),
.B(n_1473),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1506),
.A2(n_1458),
.B1(n_1475),
.B2(n_1461),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1516),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1492),
.A2(n_1469),
.B(n_1462),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1483),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1498),
.B(n_1451),
.Y(n_1530)
);

OAI31xp33_ASAP7_75t_L g1531 ( 
.A1(n_1494),
.A2(n_1459),
.A3(n_1471),
.B(n_1369),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1512),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1500),
.B(n_1468),
.Y(n_1533)
);

AOI21xp33_ASAP7_75t_L g1534 ( 
.A1(n_1486),
.A2(n_1481),
.B(n_1469),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1487),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1496),
.Y(n_1536)
);

AOI211xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1497),
.A2(n_1459),
.B(n_1447),
.C(n_1477),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1515),
.B(n_1464),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1488),
.B(n_1447),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1489),
.Y(n_1540)
);

AOI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1486),
.A2(n_1481),
.B(n_1480),
.Y(n_1541)
);

OAI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1518),
.A2(n_1482),
.B1(n_1477),
.B2(n_1439),
.C(n_1413),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1488),
.B(n_1413),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1522),
.B(n_1502),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1527),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1520),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1532),
.B(n_1503),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1519),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1523),
.B(n_1508),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1537),
.B(n_1486),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1520),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1521),
.B(n_1508),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1513),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1543),
.B(n_1486),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1530),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1538),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1536),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1531),
.A2(n_1496),
.B(n_1501),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1539),
.B(n_1513),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1561),
.A2(n_1525),
.B(n_1531),
.Y(n_1563)
);

NOR4xp25_ASAP7_75t_L g1564 ( 
.A(n_1556),
.B(n_1529),
.C(n_1540),
.D(n_1528),
.Y(n_1564)
);

AOI211xp5_ASAP7_75t_L g1565 ( 
.A1(n_1550),
.A2(n_1541),
.B(n_1534),
.C(n_1542),
.Y(n_1565)
);

OAI32xp33_ASAP7_75t_L g1566 ( 
.A1(n_1550),
.A2(n_1538),
.A3(n_1519),
.B1(n_1540),
.B2(n_1535),
.Y(n_1566)
);

OAI21xp33_ASAP7_75t_L g1567 ( 
.A1(n_1558),
.A2(n_1543),
.B(n_1535),
.Y(n_1567)
);

NOR4xp25_ASAP7_75t_L g1568 ( 
.A(n_1559),
.B(n_1519),
.C(n_1505),
.D(n_1493),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_L g1569 ( 
.A(n_1548),
.B(n_1489),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1545),
.A2(n_1505),
.B1(n_1511),
.B2(n_1490),
.C(n_1507),
.Y(n_1570)
);

OAI32xp33_ASAP7_75t_L g1571 ( 
.A1(n_1562),
.A2(n_1507),
.A3(n_1493),
.B1(n_1511),
.B2(n_1490),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1555),
.B(n_1510),
.Y(n_1572)
);

OAI222xp33_ASAP7_75t_L g1573 ( 
.A1(n_1557),
.A2(n_1509),
.B1(n_1517),
.B2(n_1514),
.C1(n_1426),
.C2(n_1373),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1569),
.Y(n_1574)
);

NOR2xp67_ASAP7_75t_L g1575 ( 
.A(n_1572),
.B(n_1548),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1563),
.B(n_1557),
.Y(n_1576)
);

NOR2x1_ASAP7_75t_L g1577 ( 
.A(n_1573),
.B(n_1545),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1571),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1567),
.B(n_1553),
.Y(n_1579)
);

AOI211x1_ASAP7_75t_L g1580 ( 
.A1(n_1566),
.A2(n_1552),
.B(n_1549),
.C(n_1544),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1564),
.B(n_1547),
.C(n_1551),
.Y(n_1581)
);

OAI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1568),
.A2(n_1560),
.B1(n_1546),
.B2(n_1509),
.Y(n_1582)
);

NAND4xp25_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1554),
.C(n_1560),
.D(n_1546),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1574),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1575),
.B(n_1570),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1580),
.B(n_1517),
.Y(n_1587)
);

NAND4xp75_ASAP7_75t_L g1588 ( 
.A(n_1577),
.B(n_1127),
.C(n_1218),
.D(n_1426),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1582),
.B(n_1420),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1587),
.B(n_1578),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1585),
.Y(n_1591)
);

NOR2xp67_ASAP7_75t_L g1592 ( 
.A(n_1586),
.B(n_1583),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1584),
.B(n_1581),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1588),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1589),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1591),
.B(n_1579),
.Y(n_1596)
);

NAND4xp75_ASAP7_75t_L g1597 ( 
.A(n_1593),
.B(n_1592),
.C(n_1590),
.D(n_1595),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1594),
.Y(n_1598)
);

AND3x4_ASAP7_75t_L g1599 ( 
.A(n_1590),
.B(n_1394),
.C(n_1401),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1593),
.B(n_1420),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1596),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1598),
.B(n_1438),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1597),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1603),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1604),
.B(n_1601),
.C(n_1603),
.Y(n_1605)
);

AO221x1_ASAP7_75t_L g1606 ( 
.A1(n_1605),
.A2(n_1603),
.B1(n_1599),
.B2(n_1602),
.C(n_1600),
.Y(n_1606)
);

AOI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1605),
.A2(n_1602),
.B(n_1207),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1606),
.Y(n_1608)
);

AOI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1607),
.A2(n_1602),
.B1(n_1127),
.B2(n_1218),
.C(n_1431),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1608),
.A2(n_1148),
.B(n_1431),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_1434),
.B(n_1432),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1610),
.B(n_1411),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1612),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_1611),
.B1(n_1411),
.B2(n_1415),
.C(n_1434),
.Y(n_1614)
);

AOI211xp5_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_1136),
.B(n_1140),
.C(n_1426),
.Y(n_1615)
);


endmodule