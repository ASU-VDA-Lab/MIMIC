module fake_jpeg_8111_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_55),
.B(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_0),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_18),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_1),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_45),
.B(n_56),
.C(n_54),
.Y(n_71)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_52),
.B(n_5),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_47),
.B1(n_1),
.B2(n_9),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_76),
.B1(n_30),
.B2(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_84),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

AOI211xp5_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_93),
.B(n_87),
.C(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_86),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_74),
.C(n_82),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_32),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_33),
.C(n_34),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_36),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_83),
.C(n_40),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_39),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_41),
.Y(n_107)
);


endmodule