module fake_jpeg_3230_n_117 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_50),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_34),
.B1(n_39),
.B2(n_32),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_33),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_58),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_41),
.B(n_37),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_47),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_39),
.B1(n_41),
.B2(n_33),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_63),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_29),
.B1(n_45),
.B2(n_42),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_47),
.B(n_1),
.C(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_6),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_5),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_5),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_14),
.A3(n_25),
.B1(n_23),
.B2(n_22),
.C1(n_11),
.C2(n_12),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_71),
.C(n_15),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_95),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_17),
.B1(n_27),
.B2(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_82),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_105),
.C(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_82),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_97),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_86),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_108),
.Y(n_109)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_100),
.B1(n_102),
.B2(n_97),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_103),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_7),
.C(n_8),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_10),
.B(n_58),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_116),
.Y(n_117)
);


endmodule