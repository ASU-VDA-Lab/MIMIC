module real_jpeg_4016_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_1),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_1),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_1),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_1),
.B(n_123),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_1),
.B(n_213),
.Y(n_348)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_2),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_3),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_4),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_4),
.B(n_100),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_4),
.B(n_182),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_4),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_4),
.B(n_50),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_5),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_5),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_5),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_5),
.B(n_371),
.Y(n_370)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_7),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_7),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_7),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_8),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_8),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_8),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_8),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_8),
.B(n_267),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_8),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_9),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_9),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_9),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_9),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_9),
.B(n_179),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_9),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_9),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_9),
.B(n_360),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_10),
.Y(n_353)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_12),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_12),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_12),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_12),
.B(n_179),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_12),
.B(n_100),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_14),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_14),
.B(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_15),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_16),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_16),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_16),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_16),
.B(n_100),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_16),
.B(n_88),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_16),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_16),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_17),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_17),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_17),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_17),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_17),
.B(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_192),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_191),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_149),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_22),
.B(n_149),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g441 ( 
.A(n_22),
.Y(n_441)
);

FAx1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_95),
.CI(n_124),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_61),
.C(n_74),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_24),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.C(n_48),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_25),
.B(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_32),
.C(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_28),
.B1(n_44),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_42),
.C(n_44),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_31),
.A2(n_32),
.B1(n_101),
.B2(n_105),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_101),
.C(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_35),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_39),
.Y(n_161)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_41),
.B(n_48),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_42),
.B(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_44),
.Y(n_170)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_49),
.B(n_53),
.C(n_57),
.Y(n_146)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_50),
.Y(n_318)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_55),
.Y(n_167)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_56),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_60),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_74),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_67),
.C(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_67),
.A2(n_68),
.B1(n_90),
.B2(n_91),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_75),
.C(n_90),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_71),
.Y(n_215)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_72),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_76),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.C(n_87),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_77),
.B(n_87),
.Y(n_157)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_82),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_86),
.Y(n_303)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_105),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_104),
.Y(n_271)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_120),
.Y(n_148)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_143),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_142),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_147),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_147),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

FAx1_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_152),
.CI(n_154),
.CON(n_195),
.SN(n_195)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_171),
.C(n_173),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_155),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_168),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_156),
.B(n_425),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_158),
.A2(n_159),
.B1(n_168),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_160),
.B(n_166),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_162),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_168),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_173),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.C(n_187),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_181),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_175),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_181),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_180),
.Y(n_369)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_184),
.Y(n_283)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_184),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_187),
.Y(n_233)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_251),
.B(n_439),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_195),
.B(n_196),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_195),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_203),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_198),
.B(n_201),
.Y(n_435)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_203),
.B(n_435),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_231),
.C(n_234),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_205),
.B(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_216),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_206),
.A2(n_207),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_209),
.A2(n_210),
.B(n_212),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_209),
.B(n_216),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_226),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_226),
.B(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_227),
.B(n_318),
.Y(n_317)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_230),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_234),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.C(n_248),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_236),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.C(n_244),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_237),
.B(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_241),
.A2(n_244),
.B1(n_245),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_241),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_246),
.B(n_248),
.Y(n_417)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_433),
.B(n_438),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_420),
.B(n_432),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_402),
.B(n_419),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_376),
.B(n_401),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_343),
.B(n_375),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_310),
.B(n_342),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_293),
.B(n_309),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_276),
.B(n_292),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_272),
.B(n_275),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_268),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_266),
.Y(n_277)
);

INVx4_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_284),
.B2(n_285),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_287),
.C(n_290),
.Y(n_308)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_290),
.B2(n_291),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_308),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_308),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_299),
.C(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_298),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_328),
.C(n_329),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_313),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_327),
.C(n_330),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_317),
.C(n_319),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_322),
.B2(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_325),
.Y(n_354)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_339),
.C(n_340),
.Y(n_373)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_336),
.Y(n_340)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_339),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_374),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_374),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_356),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_355),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_355),
.C(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_349),
.Y(n_391)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_390),
.C(n_391),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_364),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_366),
.C(n_372),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_363),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_362),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_362),
.C(n_363),
.Y(n_387)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_372),
.B2(n_373),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_370),
.Y(n_386)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_399),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_399),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_388),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_380),
.C(n_388),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_411),
.C(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_386),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_393),
.C(n_398),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_397),
.B2(n_398),
.Y(n_392)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_418),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_418),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_409),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_408),
.C(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_414),
.C(n_416),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_430),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_430),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_427),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_427),
.C(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_436),
.Y(n_438)
);


endmodule