module fake_jpeg_2780_n_76 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_76);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_35),
.B1(n_18),
.B2(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_27),
.B1(n_19),
.B2(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_24),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_0),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_5),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_9),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_10),
.C(n_11),
.Y(n_58)
);

XOR2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_12),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_67),
.C(n_65),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g76 ( 
.A(n_75),
.Y(n_76)
);


endmodule