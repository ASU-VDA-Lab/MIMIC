module fake_ibex_1028_n_210 (n_7, n_20, n_40, n_17, n_25, n_36, n_41, n_43, n_18, n_3, n_22, n_28, n_32, n_39, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_38, n_42, n_15, n_37, n_24, n_31, n_44, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_210);

input n_7;
input n_20;
input n_40;
input n_17;
input n_25;
input n_36;
input n_41;
input n_43;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_38;
input n_42;
input n_15;
input n_37;
input n_24;
input n_31;
input n_44;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_210;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_208;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_171;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_205;
wire n_204;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_177;
wire n_203;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_67;
wire n_209;
wire n_164;
wire n_198;
wire n_124;
wire n_110;
wire n_193;
wire n_47;
wire n_169;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_121;
wire n_109;
wire n_127;
wire n_175;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_191;
wire n_178;
wire n_62;
wire n_71;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_180;
wire n_194;
wire n_122;
wire n_116;
wire n_61;
wire n_201;
wire n_94;
wire n_134;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_172;
wire n_49;
wire n_66;
wire n_74;
wire n_90;
wire n_176;
wire n_58;
wire n_192;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_72;
wire n_206;
wire n_166;
wire n_195;
wire n_163;
wire n_188;
wire n_200;
wire n_114;
wire n_199;
wire n_97;
wire n_102;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_52;
wire n_189;
wire n_99;
wire n_156;
wire n_105;
wire n_135;
wire n_126;
wire n_187;
wire n_154;
wire n_182;
wire n_111;
wire n_196;
wire n_104;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_149;
wire n_54;
wire n_186;
wire n_50;
wire n_92;
wire n_144;
wire n_170;
wire n_101;
wire n_190;
wire n_113;
wire n_138;
wire n_96;
wire n_185;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_202;
wire n_158;
wire n_132;
wire n_174;
wire n_157;
wire n_160;
wire n_184;
wire n_56;
wire n_146;
wire n_91;
wire n_207;
wire n_45;

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp67_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_5),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_33),
.B(n_38),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_69),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_53),
.B(n_3),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_3),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_8),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

OR2x6_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_29),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_17),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_18),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_72),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_65),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_61),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_66),
.B(n_71),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

O2A1O1Ixp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_75),
.B(n_98),
.C(n_110),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_100),
.B(n_90),
.C(n_95),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_111),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_101),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_102),
.B(n_107),
.Y(n_137)
);

CKINVDCx10_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_100),
.C(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_126),
.B1(n_122),
.B2(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_96),
.B(n_101),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_93),
.B(n_104),
.C(n_97),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_117),
.B(n_119),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_112),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_114),
.C(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_109),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_128),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_108),
.B(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_103),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_92),
.A2(n_125),
.B(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_121),
.B(n_89),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_129),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_127),
.B(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_127),
.B1(n_139),
.B2(n_136),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_136),
.Y(n_166)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_140),
.B1(n_130),
.B2(n_133),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_134),
.B(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_145),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_158),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_137),
.B(n_142),
.C(n_161),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_150),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_150),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_152),
.B(n_135),
.Y(n_178)
);

OR2x6_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_154),
.B(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_158),
.B(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_170),
.C(n_165),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_174),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_172),
.B(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_167),
.Y(n_195)
);

AOI222xp33_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_166),
.B1(n_167),
.B2(n_131),
.C1(n_144),
.C2(n_179),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_175),
.B1(n_179),
.B2(n_185),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_184),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_198),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_201),
.Y(n_202)
);

NAND5xp2_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_196),
.C(n_197),
.D(n_195),
.E(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

NAND2x1p5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_204),
.Y(n_206)
);

OAI221xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_205),
.B1(n_192),
.B2(n_195),
.C(n_199),
.Y(n_207)
);

OAI21x1_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_189),
.B(n_186),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_188),
.B(n_191),
.Y(n_209)
);

OAI221xp5_ASAP7_75t_R g210 ( 
.A1(n_209),
.A2(n_184),
.B1(n_189),
.B2(n_186),
.C(n_188),
.Y(n_210)
);


endmodule