module real_jpeg_18316_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_1),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_1),
.A2(n_82),
.A3(n_283),
.B1(n_284),
.B2(n_287),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_1),
.A2(n_184),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_1),
.B(n_112),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_1),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_1),
.B(n_374),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_17),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_3),
.A2(n_33),
.B1(n_75),
.B2(n_176),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_3),
.A2(n_33),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_3),
.A2(n_33),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_5),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_5),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_5),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_67),
.B1(n_69),
.B2(n_74),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_7),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_9),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_9),
.A2(n_103),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_103),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_9),
.A2(n_32),
.B1(n_103),
.B2(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

BUFx4f_ASAP7_75t_L g198 ( 
.A(n_12),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_467),
.B(n_470),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_274),
.B(n_461),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_248),
.C(n_268),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_215),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_22),
.A2(n_463),
.B(n_464),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_157),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_23),
.B(n_157),
.Y(n_464)
);

XOR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_147),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_145),
.B2(n_146),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_25),
.B(n_146),
.C(n_147),
.Y(n_249)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_63),
.B2(n_64),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_27),
.A2(n_28),
.B1(n_218),
.B2(n_299),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_27),
.A2(n_28),
.B1(n_174),
.B2(n_375),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_28),
.B(n_218),
.C(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_28),
.B(n_65),
.C(n_113),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_28),
.B(n_174),
.C(n_435),
.Y(n_434)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_47),
.B2(n_55),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_29),
.A2(n_34),
.B1(n_47),
.B2(n_55),
.Y(n_145)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_34),
.B(n_47),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_34),
.Y(n_266)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_42),
.B(n_47),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_35),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_37),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_44),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_46),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g405 ( 
.A(n_46),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_47),
.A2(n_255),
.B(n_264),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_47),
.A2(n_255),
.B1(n_266),
.B2(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_47),
.Y(n_374)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_53),
.Y(n_156)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_55),
.Y(n_213)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_58),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_59),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_59),
.B(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_113),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_79),
.B1(n_102),
.B2(n_112),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_66),
.A2(n_79),
.B1(n_112),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_67),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_68),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_68),
.A2(n_170),
.B1(n_229),
.B2(n_233),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_69),
.A2(n_393),
.B1(n_402),
.B2(n_406),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_73),
.Y(n_401)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_77),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_80),
.A2(n_92),
.B1(n_151),
.B2(n_175),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_80),
.A2(n_92),
.B1(n_151),
.B2(n_175),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_80),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g427 ( 
.A1(n_80),
.A2(n_92),
.B(n_151),
.Y(n_427)
);

NAND2x1p5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_92),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_92),
.B(n_253),
.Y(n_252)
);

OA22x2_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_97),
.Y(n_322)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_102),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_149),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_136),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_115),
.A2(n_164),
.B(n_182),
.Y(n_181)
);

AOI21x1_ASAP7_75t_SL g385 ( 
.A1(n_115),
.A2(n_386),
.B(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_126),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g220 ( 
.A1(n_116),
.A2(n_125),
.B1(n_183),
.B2(n_221),
.Y(n_220)
);

AO22x2_ASAP7_75t_L g298 ( 
.A1(n_116),
.A2(n_125),
.B1(n_183),
.B2(n_221),
.Y(n_298)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_123),
.Y(n_116)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_122),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B1(n_132),
.B2(n_135),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_135),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_163),
.B1(n_172),
.B2(n_173),
.Y(n_162)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_145),
.B(n_427),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_148),
.C(n_149),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_146),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_146),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_146),
.B(n_299),
.C(n_385),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_155),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_155),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_178),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_162),
.B(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_174),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_169),
.A2(n_170),
.B1(n_256),
.B2(n_260),
.Y(n_255)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_171),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_173),
.B(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_174),
.A2(n_370),
.B1(n_371),
.B2(n_375),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_174),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_174),
.B(n_348),
.C(n_373),
.Y(n_389)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_193),
.B(n_211),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_192),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_181),
.A2(n_192),
.B1(n_193),
.B2(n_418),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_181),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_183),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B(n_189),
.Y(n_183)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_189),
.A2(n_205),
.A3(n_319),
.B1(n_323),
.B2(n_327),
.Y(n_318)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_191),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_193),
.B1(n_211),
.B2(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_228),
.B1(n_235),
.B2(n_236),
.Y(n_227)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_200),
.Y(n_293)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_200),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_201),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_202),
.B(n_291),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_207),
.Y(n_347)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_214),
.B(n_469),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_245),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_216),
.B(n_245),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_241),
.C(n_242),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_217),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_218),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_297)
);

INVx3_ASAP7_75t_SL g299 ( 
.A(n_218),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_218),
.A2(n_299),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_219),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_227),
.Y(n_219)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_220),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_220),
.B(n_314),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_220),
.A2(n_302),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_220),
.A2(n_227),
.B1(n_302),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_227),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_228),
.A2(n_351),
.B(n_422),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_232),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g303 ( 
.A1(n_235),
.A2(n_290),
.B1(n_304),
.B2(n_310),
.Y(n_303)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_240),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_241),
.B(n_243),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g461 ( 
.A1(n_248),
.A2(n_268),
.B(n_462),
.C(n_465),
.D(n_466),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_249),
.B(n_250),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g473 ( 
.A(n_250),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.CI(n_267),
.CON(n_250),
.SN(n_250)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_254),
.C(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_269),
.B(n_273),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_269),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_269),
.B(n_468),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_270),
.Y(n_469)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

AO221x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_408),
.B1(n_410),
.B2(n_454),
.C(n_460),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_379),
.B(n_407),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_363),
.B(n_378),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_315),
.B(n_362),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_301),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_280),
.B(n_301),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_297),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_281),
.B(n_298),
.C(n_299),
.Y(n_377)
);

XOR2x2_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_289),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_282),
.B(n_289),
.Y(n_366)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_298),
.A2(n_300),
.B1(n_318),
.B2(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_298),
.B(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_298),
.A2(n_300),
.B1(n_421),
.B2(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.C(n_314),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_302),
.B(n_366),
.C(n_368),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_303),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_353),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_303),
.A2(n_334),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_349),
.B(n_351),
.Y(n_348)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

AOI21x1_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_337),
.B(n_361),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_333),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g361 ( 
.A(n_317),
.B(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_334),
.B(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_356),
.B(n_360),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_352),
.B(n_355),
.Y(n_338)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_357),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_357),
.B(n_358),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_377),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_377),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_368),
.B1(n_369),
.B2(n_376),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_365),
.Y(n_376)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_366),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_381),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_388),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_382),
.B(n_389),
.C(n_390),
.Y(n_440)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_438),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_428),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_R g460 ( 
.A(n_411),
.B(n_413),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.C(n_419),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_417),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.C(n_426),
.Y(n_419)
);

XNOR2x1_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_431),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_436),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_436),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.C(n_434),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_432),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_450),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_441),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_446),
.C(n_448),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_453),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_456),
.B(n_458),
.C(n_459),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_471),
.Y(n_470)
);


endmodule