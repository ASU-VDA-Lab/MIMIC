module real_aes_18148_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_0), .Y(n_522) );
AND2x4_ASAP7_75t_L g110 ( .A(n_1), .B(n_111), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_2), .A2(n_4), .B1(n_192), .B2(n_193), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_3), .A2(n_21), .B1(n_143), .B2(n_145), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_5), .A2(n_51), .B1(n_210), .B2(n_211), .Y(n_209) );
BUFx3_ASAP7_75t_L g552 ( .A(n_6), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_7), .A2(n_14), .B1(n_150), .B2(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_9), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_10), .A2(n_100), .B1(n_116), .B2(n_843), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_11), .B(n_190), .Y(n_558) );
BUFx2_ASAP7_75t_L g104 ( .A(n_12), .Y(n_104) );
OR2x2_ASAP7_75t_L g124 ( .A(n_12), .B(n_30), .Y(n_124) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_15), .B(n_207), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_16), .B(n_228), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_17), .A2(n_83), .B1(n_143), .B2(n_207), .Y(n_529) );
OAI22xp33_ASAP7_75t_L g131 ( .A1(n_18), .A2(n_132), .B1(n_497), .B2(n_498), .Y(n_131) );
INVx1_ASAP7_75t_L g497 ( .A(n_18), .Y(n_497) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_19), .A2(n_47), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_20), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_22), .B(n_145), .Y(n_572) );
INVx4_ASAP7_75t_R g236 ( .A(n_23), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_24), .B(n_148), .Y(n_173) );
AO32x1_ASAP7_75t_L g526 ( .A1(n_25), .A2(n_156), .A3(n_157), .B1(n_527), .B2(n_530), .Y(n_526) );
AO32x2_ASAP7_75t_L g623 ( .A1(n_25), .A2(n_156), .A3(n_157), .B1(n_527), .B2(n_530), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_26), .B(n_145), .Y(n_182) );
INVx1_ASAP7_75t_L g200 ( .A(n_27), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_SL g278 ( .A1(n_28), .A2(n_147), .B(n_150), .C(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_29), .A2(n_44), .B1(n_150), .B2(n_151), .Y(n_149) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_31), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_32), .A2(n_50), .B1(n_145), .B2(n_237), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_33), .A2(n_89), .B1(n_143), .B2(n_151), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_34), .B(n_560), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_35), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_36), .B(n_581), .Y(n_601) );
INVx1_ASAP7_75t_L g179 ( .A(n_37), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_38), .B(n_150), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_39), .A2(n_66), .B1(n_151), .B2(n_535), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_40), .Y(n_259) );
INVx2_ASAP7_75t_L g501 ( .A(n_41), .Y(n_501) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
BUFx3_ASAP7_75t_L g827 ( .A(n_42), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_43), .B(n_603), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_45), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_46), .A2(n_82), .B1(n_150), .B2(n_151), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_48), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_49), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_52), .A2(n_76), .B1(n_175), .B2(n_581), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_53), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_54), .A2(n_80), .B1(n_143), .B2(n_207), .Y(n_548) );
INVx1_ASAP7_75t_L g159 ( .A(n_55), .Y(n_159) );
AND2x4_ASAP7_75t_L g161 ( .A(n_56), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_57), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_58), .A2(n_88), .B1(n_151), .B2(n_189), .Y(n_188) );
AO22x1_ASAP7_75t_L g205 ( .A1(n_59), .A2(n_71), .B1(n_174), .B2(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_60), .B(n_143), .Y(n_557) );
INVx1_ASAP7_75t_L g162 ( .A(n_61), .Y(n_162) );
AND2x2_ASAP7_75t_L g281 ( .A(n_62), .B(n_156), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_63), .B(n_156), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_64), .A2(n_153), .B(n_210), .C(n_521), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_65), .B(n_143), .C(n_562), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_67), .B(n_210), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_68), .Y(n_274) );
AND2x2_ASAP7_75t_L g523 ( .A(n_69), .B(n_241), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_70), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_72), .B(n_145), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_73), .A2(n_94), .B1(n_175), .B2(n_207), .Y(n_583) );
INVx2_ASAP7_75t_L g148 ( .A(n_74), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_75), .B(n_261), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_77), .B(n_156), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_78), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_79), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_81), .B(n_166), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_84), .B(n_562), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g503 ( .A1(n_85), .A2(n_504), .B1(n_820), .B2(n_821), .Y(n_503) );
INVx1_ASAP7_75t_L g820 ( .A(n_85), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_85), .A2(n_498), .B1(n_820), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_86), .A2(n_98), .B1(n_151), .B2(n_237), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_87), .B(n_581), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_90), .B(n_156), .Y(n_256) );
INVx1_ASAP7_75t_L g115 ( .A(n_91), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_91), .B(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_92), .B(n_228), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_93), .A2(n_196), .B(n_210), .C(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g240 ( .A(n_95), .B(n_241), .Y(n_240) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_96), .B(n_190), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_97), .Y(n_571) );
INVx3_ASAP7_75t_L g843 ( .A(n_100), .Y(n_843) );
INVx8_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_107), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .C(n_114), .Y(n_108) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g122 ( .A(n_113), .Y(n_122) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_114), .Y(n_828) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g832 ( .A(n_115), .Y(n_832) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_125), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_117), .A2(n_127), .B(n_131), .Y(n_126) );
NOR2xp67_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
CKINVDCx8_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
INVx4_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
AND2x6_ASAP7_75t_SL g120 ( .A(n_121), .B(n_123), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_123), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR2x1_ASAP7_75t_L g842 ( .A(n_124), .B(n_827), .Y(n_842) );
OAI21xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_499), .B(n_502), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx12f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g498 ( .A(n_132), .Y(n_498) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_132), .Y(n_834) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_374), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_322), .Y(n_133) );
OAI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_201), .B(n_242), .C(n_307), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_137), .A2(n_243), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_167), .Y(n_137) );
INVx2_ASAP7_75t_L g303 ( .A(n_138), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_138), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g414 ( .A(n_139), .B(n_169), .Y(n_414) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_SL g282 ( .A(n_140), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_140), .B(n_185), .Y(n_319) );
AND2x2_ASAP7_75t_L g352 ( .A(n_140), .B(n_269), .Y(n_352) );
OR2x2_ASAP7_75t_L g357 ( .A(n_140), .B(n_185), .Y(n_357) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_155), .A3(n_160), .B(n_163), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B1(n_149), .B2(n_152), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_143), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_SL g581 ( .A(n_143), .Y(n_581) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_144), .Y(n_145) );
INVx3_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
INVx1_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_144), .Y(n_207) );
INVx1_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
INVx1_ASAP7_75t_L g237 ( .A(n_144), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_145), .B(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_145), .A2(n_237), .B1(n_517), .B2(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g535 ( .A(n_145), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_146), .A2(n_188), .B1(n_191), .B2(n_195), .Y(n_187) );
OAI22x1_ASAP7_75t_L g217 ( .A1(n_146), .A2(n_195), .B1(n_218), .B2(n_220), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_146), .A2(n_152), .B1(n_534), .B2(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_146), .A2(n_147), .B1(n_548), .B2(n_549), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_146), .A2(n_580), .B1(n_582), .B2(n_583), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_146), .A2(n_601), .B(n_602), .Y(n_600) );
INVx6_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_147), .A2(n_205), .B(n_208), .C(n_214), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_147), .A2(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_147), .B(n_205), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_147), .A2(n_277), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_147), .A2(n_557), .B(n_558), .Y(n_556) );
BUFx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx1_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
INVx4_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_151), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
INVx2_ASAP7_75t_L g560 ( .A(n_151), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_152), .A2(n_181), .B(n_182), .Y(n_180) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_152), .A2(n_209), .B(n_213), .Y(n_208) );
AOI21x1_ASAP7_75t_L g597 ( .A1(n_152), .A2(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g262 ( .A(n_154), .Y(n_262) );
AOI31xp67_ASAP7_75t_L g546 ( .A1(n_155), .A2(n_160), .A3(n_547), .B(n_550), .Y(n_546) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_156), .B(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g183 ( .A(n_157), .B(n_160), .Y(n_183) );
BUFx3_ASAP7_75t_L g532 ( .A(n_157), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_157), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_157), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g568 ( .A(n_157), .Y(n_568) );
INVx2_ASAP7_75t_SL g595 ( .A(n_157), .Y(n_595) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
INVx1_ASAP7_75t_L g267 ( .A(n_160), .Y(n_267) );
OAI21x1_ASAP7_75t_L g555 ( .A1(n_160), .A2(n_556), .B(n_559), .Y(n_555) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_160), .A2(n_570), .B(n_573), .Y(n_569) );
BUFx10_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
BUFx10_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
AO31x2_ASAP7_75t_L g531 ( .A1(n_161), .A2(n_532), .A3(n_533), .B(n_537), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
BUFx2_ASAP7_75t_L g186 ( .A(n_165), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_165), .B(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_165), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g241 ( .A(n_165), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_165), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI21xp33_ASAP7_75t_L g214 ( .A1(n_166), .A2(n_213), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
INVx2_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g496 ( .A(n_168), .Y(n_496) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_184), .Y(n_168) );
AND2x2_ASAP7_75t_L g297 ( .A(n_169), .B(n_185), .Y(n_297) );
INVx3_ASAP7_75t_L g305 ( .A(n_169), .Y(n_305) );
NAND2x1p5_ASAP7_75t_SL g337 ( .A(n_169), .B(n_321), .Y(n_337) );
INVx1_ASAP7_75t_L g355 ( .A(n_169), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_169), .B(n_300), .Y(n_380) );
BUFx2_ASAP7_75t_L g466 ( .A(n_169), .Y(n_466) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_180), .B(n_183), .Y(n_171) );
OAI21xp33_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_176), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_175), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
BUFx4f_ASAP7_75t_L g277 ( .A(n_178), .Y(n_277) );
INVx1_ASAP7_75t_L g562 ( .A(n_178), .Y(n_562) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g250 ( .A(n_185), .Y(n_250) );
INVx1_ASAP7_75t_L g306 ( .A(n_185), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_185), .B(n_282), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_185), .B(n_269), .Y(n_415) );
AO31x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .A3(n_197), .B(n_199), .Y(n_185) );
AOI21x1_ASAP7_75t_L g270 ( .A1(n_186), .A2(n_271), .B(n_281), .Y(n_270) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_190), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_235) );
O2A1O1Ixp5_ASAP7_75t_L g570 ( .A1(n_193), .A2(n_277), .B(n_571), .C(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_194), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_195), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g519 ( .A(n_196), .Y(n_519) );
INVx1_ASAP7_75t_SL g582 ( .A(n_196), .Y(n_582) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_197), .A2(n_532), .A3(n_579), .B(n_584), .Y(n_578) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_SL g530 ( .A(n_198), .Y(n_530) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_225), .Y(n_201) );
INVx1_ASAP7_75t_L g473 ( .A(n_202), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
OR2x2_ASAP7_75t_L g245 ( .A(n_203), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g310 ( .A(n_203), .Y(n_310) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVxp67_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g603 ( .A(n_207), .Y(n_603) );
INVx1_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_212), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_215), .A2(n_272), .B(n_278), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_215), .A2(n_515), .B(n_520), .Y(n_514) );
INVx2_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
OR2x2_ASAP7_75t_L g311 ( .A(n_216), .B(n_226), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_216), .B(n_226), .Y(n_316) );
INVx2_ASAP7_75t_L g361 ( .A(n_216), .Y(n_361) );
AND2x2_ASAP7_75t_L g402 ( .A(n_216), .B(n_255), .Y(n_402) );
AND2x2_ASAP7_75t_L g436 ( .A(n_216), .B(n_333), .Y(n_436) );
AO31x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_221), .A3(n_222), .B(n_223), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_219), .A2(n_259), .B(n_260), .C(n_261), .Y(n_258) );
INVx2_ASAP7_75t_L g554 ( .A(n_221), .Y(n_554) );
INVx2_ASAP7_75t_L g239 ( .A(n_222), .Y(n_239) );
INVx1_ASAP7_75t_L g247 ( .A(n_225), .Y(n_247) );
INVx1_ASAP7_75t_L g366 ( .A(n_225), .Y(n_366) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g286 ( .A(n_226), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g327 ( .A(n_226), .B(n_288), .Y(n_327) );
INVx2_ASAP7_75t_L g333 ( .A(n_226), .Y(n_333) );
AND2x2_ASAP7_75t_L g388 ( .A(n_226), .B(n_255), .Y(n_388) );
AND2x2_ASAP7_75t_L g445 ( .A(n_226), .B(n_254), .Y(n_445) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_240), .Y(n_226) );
AOI21x1_ASAP7_75t_L g513 ( .A1(n_227), .A2(n_514), .B(n_523), .Y(n_513) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_234), .B(n_239), .Y(n_230) );
INVx1_ASAP7_75t_L g575 ( .A(n_237), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B1(n_283), .B2(n_294), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NAND3xp33_ASAP7_75t_SL g423 ( .A(n_245), .B(n_424), .C(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g342 ( .A(n_246), .Y(n_342) );
AND2x2_ASAP7_75t_L g392 ( .A(n_246), .B(n_254), .Y(n_392) );
INVx1_ASAP7_75t_L g492 ( .A(n_247), .Y(n_492) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_249), .B(n_447), .Y(n_483) );
BUFx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g338 ( .A(n_250), .Y(n_338) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_268), .Y(n_252) );
INVx1_ASAP7_75t_L g326 ( .A(n_253), .Y(n_326) );
BUFx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g406 ( .A(n_254), .B(n_287), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_254), .B(n_332), .Y(n_425) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g293 ( .A(n_255), .Y(n_293) );
BUFx3_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
AND2x2_ASAP7_75t_L g360 ( .A(n_255), .B(n_361), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_263), .B(n_266), .Y(n_257) );
INVx2_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_262), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_573) );
INVx2_ASAP7_75t_L g453 ( .A(n_268), .Y(n_453) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_282), .Y(n_268) );
INVx2_ASAP7_75t_L g321 ( .A(n_269), .Y(n_321) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g300 ( .A(n_270), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_285), .B(n_292), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g340 ( .A(n_286), .B(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g470 ( .A(n_286), .Y(n_470) );
INVx1_ASAP7_75t_L g315 ( .A(n_287), .Y(n_315) );
AND2x2_ASAP7_75t_L g395 ( .A(n_287), .B(n_333), .Y(n_395) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g332 ( .A(n_288), .B(n_333), .Y(n_332) );
AOI21x1_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_293), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g428 ( .A(n_293), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_302), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_295), .A2(n_336), .B1(n_339), .B2(n_343), .Y(n_335) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_296), .A2(n_316), .B1(n_348), .B2(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
BUFx2_ASAP7_75t_SL g334 ( .A(n_297), .Y(n_334) );
AND2x4_ASAP7_75t_L g452 ( .A(n_297), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g461 ( .A(n_297), .Y(n_461) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g373 ( .A(n_299), .Y(n_373) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_300), .B(n_305), .Y(n_431) );
INVxp67_ASAP7_75t_L g460 ( .A(n_300), .Y(n_460) );
AND2x2_ASAP7_75t_L g465 ( .A(n_300), .B(n_331), .Y(n_465) );
OR2x2_ASAP7_75t_L g447 ( .A(n_301), .B(n_321), .Y(n_447) );
INVx1_ASAP7_75t_L g328 ( .A(n_302), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_303), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g367 ( .A(n_304), .B(n_352), .Y(n_367) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_305), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
OR2x2_ASAP7_75t_L g446 ( .A(n_305), .B(n_447), .Y(n_446) );
OAI21xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B(n_317), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g370 ( .A(n_309), .Y(n_370) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g364 ( .A(n_310), .B(n_361), .Y(n_364) );
INVx2_ASAP7_75t_L g488 ( .A(n_310), .Y(n_488) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AND2x2_ASAP7_75t_L g417 ( .A(n_314), .B(n_360), .Y(n_417) );
AND2x2_ASAP7_75t_L g442 ( .A(n_314), .B(n_388), .Y(n_442) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
AND2x2_ASAP7_75t_L g372 ( .A(n_316), .B(n_326), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_316), .B(n_371), .Y(n_384) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g469 ( .A(n_319), .Y(n_469) );
OR2x2_ASAP7_75t_L g485 ( .A(n_319), .B(n_380), .Y(n_485) );
INVx1_ASAP7_75t_L g409 ( .A(n_321), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_346), .C(n_368), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B1(n_329), .B2(n_334), .C(n_335), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g348 ( .A(n_327), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_327), .B(n_392), .Y(n_476) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g371 ( .A(n_331), .Y(n_371) );
AND3x1_ASAP7_75t_L g467 ( .A(n_331), .B(n_468), .C(n_469), .Y(n_467) );
AND2x2_ASAP7_75t_L g454 ( .A(n_332), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g464 ( .A(n_332), .Y(n_464) );
INVxp67_ASAP7_75t_L g478 ( .A(n_334), .Y(n_478) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g433 ( .A(n_337), .B(n_357), .Y(n_433) );
INVx2_ASAP7_75t_L g468 ( .A(n_337), .Y(n_468) );
INVx1_ASAP7_75t_L g386 ( .A(n_338), .Y(n_386) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_340), .A2(n_388), .B(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_341), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g349 ( .A(n_342), .Y(n_349) );
OR2x2_ASAP7_75t_L g443 ( .A(n_342), .B(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g403 ( .A(n_345), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_345), .B(n_402), .Y(n_482) );
AND3x1_ASAP7_75t_L g346 ( .A(n_347), .B(n_353), .C(n_358), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND2x2_ASAP7_75t_L g397 ( .A(n_349), .B(n_388), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_350), .A2(n_417), .B1(n_418), .B2(n_420), .Y(n_416) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OAI321xp33_ASAP7_75t_L g439 ( .A1(n_351), .A2(n_440), .A3(n_441), .B1(n_443), .B2(n_446), .C(n_448), .Y(n_439) );
AND2x2_ASAP7_75t_L g491 ( .A(n_351), .B(n_356), .Y(n_491) );
AND2x2_ASAP7_75t_L g389 ( .A(n_352), .B(n_355), .Y(n_389) );
INVx2_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
AND2x2_ASAP7_75t_L g407 ( .A(n_354), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g419 ( .A(n_357), .B(n_409), .Y(n_419) );
INVx2_ASAP7_75t_L g451 ( .A(n_357), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B(n_367), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g455 ( .A(n_361), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_364), .B(n_371), .Y(n_381) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_373), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_371), .B(n_395), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_371), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g472 ( .A(n_371), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g440 ( .A(n_373), .Y(n_440) );
NOR2xp67_ASAP7_75t_L g374 ( .A(n_375), .B(n_437), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_399), .C(n_422), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_390), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .B1(n_382), .B2(n_385), .C(n_387), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
OR2x2_ASAP7_75t_L g430 ( .A(n_379), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI21xp33_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_396), .B(n_398), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g427 ( .A(n_395), .B(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_SL g410 ( .A1(n_396), .A2(n_411), .B(n_416), .Y(n_410) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_404), .B(n_407), .C(n_410), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_401), .B(n_476), .Y(n_475) );
NAND2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_409), .B(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_412), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_429), .B1(n_432), .B2(n_434), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_431), .Y(n_494) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_474), .C(n_489), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_456), .Y(n_438) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
OAI21xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B(n_454), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_462), .C(n_471), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AOI32xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .A3(n_466), .B1(n_467), .B2(n_470), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g490 ( .A(n_465), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI22x1_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B1(n_484), .B2(n_486), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI21xp33_ASAP7_75t_L g493 ( .A1(n_482), .A2(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_492), .B(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x6_ASAP7_75t_SL g824 ( .A(n_500), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_501), .B(n_840), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_822), .B1(n_829), .B2(n_833), .C(n_835), .Y(n_502) );
INVx1_ASAP7_75t_L g821 ( .A(n_504), .Y(n_821) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND4xp75_ASAP7_75t_L g505 ( .A(n_506), .B(n_694), .C(n_748), .D(n_792), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_647), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_613), .Y(n_507) );
O2A1O1Ixp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_539), .B(n_543), .C(n_586), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_524), .Y(n_509) );
AND2x2_ASAP7_75t_L g664 ( .A(n_510), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g653 ( .A(n_511), .B(n_589), .Y(n_653) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_512), .Y(n_619) );
AND2x2_ASAP7_75t_L g668 ( .A(n_512), .B(n_531), .Y(n_668) );
INVx1_ASAP7_75t_L g680 ( .A(n_512), .Y(n_680) );
INVx1_ASAP7_75t_L g778 ( .A(n_512), .Y(n_778) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g541 ( .A(n_513), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_516), .B(n_519), .Y(n_515) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g606 ( .A(n_525), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_531), .Y(n_525) );
AND2x2_ASAP7_75t_L g542 ( .A(n_526), .B(n_531), .Y(n_542) );
INVx1_ASAP7_75t_L g646 ( .A(n_526), .Y(n_646) );
INVx1_ASAP7_75t_L g757 ( .A(n_526), .Y(n_757) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_530), .A2(n_597), .B(n_600), .Y(n_596) );
INVx3_ASAP7_75t_L g589 ( .A(n_531), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_531), .B(n_593), .Y(n_644) );
AND2x2_ASAP7_75t_L g679 ( .A(n_531), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g719 ( .A(n_540), .Y(n_719) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g588 ( .A(n_541), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_541), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g621 ( .A(n_541), .Y(n_621) );
OR2x2_ASAP7_75t_L g685 ( .A(n_541), .B(n_593), .Y(n_685) );
OR2x2_ASAP7_75t_L g756 ( .A(n_541), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_SL g693 ( .A(n_542), .Y(n_693) );
AND2x2_ASAP7_75t_L g745 ( .A(n_542), .B(n_608), .Y(n_745) );
AND2x2_ASAP7_75t_L g802 ( .A(n_542), .B(n_719), .Y(n_802) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_565), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_544), .B(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g811 ( .A(n_544), .B(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
INVx2_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
AND2x2_ASAP7_75t_L g637 ( .A(n_545), .B(n_616), .Y(n_637) );
AND2x2_ASAP7_75t_L g707 ( .A(n_545), .B(n_578), .Y(n_707) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g661 ( .A(n_546), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g615 ( .A(n_553), .B(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g676 ( .A(n_553), .B(n_567), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_564), .Y(n_553) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_554), .A2(n_555), .B(n_564), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g683 ( .A(n_566), .B(n_660), .Y(n_683) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_578), .Y(n_566) );
INVx2_ASAP7_75t_SL g605 ( .A(n_567), .Y(n_605) );
BUFx2_ASAP7_75t_L g658 ( .A(n_567), .Y(n_658) );
INVx1_ASAP7_75t_L g730 ( .A(n_567), .Y(n_730) );
AND2x2_ASAP7_75t_L g763 ( .A(n_567), .B(n_611), .Y(n_763) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_577), .Y(n_567) );
OA21x2_ASAP7_75t_L g616 ( .A1(n_568), .A2(n_569), .B(n_577), .Y(n_616) );
INVx2_ASAP7_75t_L g591 ( .A(n_578), .Y(n_591) );
INVx1_ASAP7_75t_L g611 ( .A(n_578), .Y(n_611) );
INVx1_ASAP7_75t_L g639 ( .A(n_578), .Y(n_639) );
AND2x2_ASAP7_75t_L g729 ( .A(n_578), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g770 ( .A(n_578), .B(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g786 ( .A(n_578), .B(n_771), .Y(n_786) );
AND2x2_ASAP7_75t_L g812 ( .A(n_578), .B(n_616), .Y(n_812) );
OAI32xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_590), .A3(n_605), .B1(n_606), .B2(n_609), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_588), .B(n_753), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_588), .B(n_791), .Y(n_790) );
AND2x4_ASAP7_75t_L g622 ( .A(n_589), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g724 ( .A(n_589), .Y(n_724) );
INVx1_ASAP7_75t_L g784 ( .A(n_589), .Y(n_784) );
INVx1_ASAP7_75t_L g722 ( .A(n_590), .Y(n_722) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_SL g626 ( .A(n_591), .Y(n_626) );
AND2x2_ASAP7_75t_L g715 ( .A(n_591), .B(n_630), .Y(n_715) );
AND2x2_ASAP7_75t_L g783 ( .A(n_592), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g608 ( .A(n_593), .Y(n_608) );
AND2x2_ASAP7_75t_L g618 ( .A(n_593), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g654 ( .A(n_593), .Y(n_654) );
AND2x2_ASAP7_75t_L g665 ( .A(n_593), .B(n_623), .Y(n_665) );
AND2x2_ASAP7_75t_L g689 ( .A(n_593), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g699 ( .A(n_593), .B(n_690), .Y(n_699) );
INVxp67_ASAP7_75t_L g753 ( .A(n_593), .Y(n_753) );
BUFx2_ASAP7_75t_L g765 ( .A(n_593), .Y(n_765) );
INVx1_ASAP7_75t_L g769 ( .A(n_593), .Y(n_769) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI21x1_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_604), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_605), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g761 ( .A(n_605), .Y(n_761) );
AND2x2_ASAP7_75t_L g669 ( .A(n_608), .B(n_646), .Y(n_669) );
AND2x2_ASAP7_75t_L g798 ( .A(n_608), .B(n_622), .Y(n_798) );
OAI22xp5_ASAP7_75t_SL g686 ( .A1(n_609), .A2(n_687), .B1(n_691), .B2(n_692), .Y(n_686) );
O2A1O1Ixp5_ASAP7_75t_R g760 ( .A1(n_609), .A2(n_761), .B(n_762), .C(n_764), .Y(n_760) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g614 ( .A(n_610), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g628 ( .A(n_612), .Y(n_628) );
INVx1_ASAP7_75t_L g671 ( .A(n_612), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_612), .B(n_641), .Y(n_747) );
AND2x2_ASAP7_75t_L g759 ( .A(n_612), .B(n_630), .Y(n_759) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B1(n_620), .B2(n_624), .C1(n_634), .C2(n_642), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_614), .A2(n_656), .B1(n_734), .B2(n_795), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_614), .A2(n_678), .B1(n_814), .B2(n_816), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_615), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_615), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g789 ( .A(n_615), .Y(n_789) );
INVx1_ASAP7_75t_L g819 ( .A(n_615), .Y(n_819) );
INVx1_ASAP7_75t_L g633 ( .A(n_616), .Y(n_633) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g688 ( .A(n_619), .Y(n_688) );
AOI321xp33_ASAP7_75t_L g766 ( .A1(n_620), .A2(n_664), .A3(n_767), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_766) );
AND2x4_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
OR2x2_ASAP7_75t_L g698 ( .A(n_621), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g718 ( .A(n_622), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g690 ( .A(n_623), .Y(n_690) );
NAND2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
OR2x2_ASAP7_75t_L g691 ( .A(n_626), .B(n_660), .Y(n_691) );
AND2x2_ASAP7_75t_L g711 ( .A(n_626), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g801 ( .A(n_627), .Y(n_801) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g732 ( .A(n_629), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_630), .B(n_633), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g641 ( .A(n_631), .Y(n_641) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g660 ( .A(n_632), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_635), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_637), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g772 ( .A(n_641), .Y(n_772) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_643), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g705 ( .A(n_644), .Y(n_705) );
INVx1_ASAP7_75t_L g655 ( .A(n_645), .Y(n_655) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_646), .Y(n_703) );
INVx2_ASAP7_75t_L g737 ( .A(n_646), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_672), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_656), .B(n_662), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_651), .B(n_655), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_652), .A2(n_739), .B1(n_789), .B2(n_790), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx2_ASAP7_75t_L g754 ( .A(n_653), .Y(n_754) );
AND2x2_ASAP7_75t_L g678 ( .A(n_654), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g692 ( .A(n_654), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g743 ( .A(n_654), .Y(n_743) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g723 ( .A(n_658), .B(n_659), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_658), .B(n_707), .Y(n_739) );
AND2x2_ASAP7_75t_L g785 ( .A(n_658), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_659), .B(n_763), .Y(n_800) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g712 ( .A(n_660), .Y(n_712) );
INVx1_ASAP7_75t_L g771 ( .A(n_661), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_670), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g733 ( .A(n_665), .B(n_688), .Y(n_733) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_668), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g742 ( .A(n_668), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_671), .B(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_686), .Y(n_672) );
OAI21xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B(n_681), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_674), .A2(n_741), .B1(n_744), .B2(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI311xp33_ASAP7_75t_L g774 ( .A1(n_676), .A2(n_775), .A3(n_776), .B(n_779), .C(n_780), .Y(n_774) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g702 ( .A(n_679), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_679), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g773 ( .A(n_683), .Y(n_773) );
INVx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx2_ASAP7_75t_L g779 ( .A(n_689), .Y(n_779) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_693), .Y(n_796) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_720), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .C(n_708), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AO21x1_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AO221x1_ASAP7_75t_L g781 ( .A1(n_702), .A2(n_782), .B1(n_785), .B2(n_787), .C(n_788), .Y(n_781) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g780 ( .A(n_707), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_713), .B(n_716), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .B(n_725), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g775 ( .A(n_724), .Y(n_775) );
AOI221x1_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_733), .B1(n_734), .B2(n_738), .C(n_740), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_731), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g758 ( .A(n_729), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AO22x1_ASAP7_75t_L g805 ( .A1(n_733), .A2(n_806), .B1(n_808), .B2(n_811), .Y(n_805) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g782 ( .A(n_736), .B(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_737), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVxp33_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_781), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_766), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_758), .B(n_760), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .C(n_756), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g791 ( .A(n_753), .Y(n_791) );
AND2x2_ASAP7_75t_L g777 ( .A(n_757), .B(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g787 ( .A(n_763), .B(n_772), .Y(n_787) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
NAND2x1p5_ASAP7_75t_L g815 ( .A(n_769), .B(n_777), .Y(n_815) );
INVx2_ASAP7_75t_L g807 ( .A(n_772), .Y(n_807) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g810 ( .A(n_778), .Y(n_810) );
AND2x2_ASAP7_75t_L g806 ( .A(n_786), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g818 ( .A(n_786), .Y(n_818) );
NOR2x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_803), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_798), .A2(n_799), .B1(n_801), .B2(n_802), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_813), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NOR2x1_ASAP7_75t_R g822 ( .A(n_823), .B(n_828), .Y(n_822) );
NOR2xp67_ASAP7_75t_SL g829 ( .A(n_823), .B(n_830), .Y(n_829) );
INVx5_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx4_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
AND2x2_ASAP7_75t_L g841 ( .A(n_832), .B(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx6_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
BUFx10_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
endmodule