module fake_jpeg_17120_n_376 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_376);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_376;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_42),
.Y(n_88)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_46),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_7),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_26),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_32),
.B1(n_34),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_68),
.A2(n_69),
.B1(n_75),
.B2(n_80),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_32),
.B1(n_30),
.B2(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_30),
.B1(n_34),
.B2(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_39),
.B(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_76),
.B(n_84),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_36),
.B1(n_33),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_78),
.A2(n_110),
.B1(n_111),
.B2(n_9),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_28),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_33),
.C(n_27),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_109),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_29),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_97),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_38),
.B(n_23),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_33),
.B(n_36),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_22),
.B(n_24),
.C(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_11),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_52),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_58),
.A2(n_20),
.B1(n_24),
.B2(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_36),
.B1(n_55),
.B2(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_20),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_36),
.B1(n_33),
.B2(n_27),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_115),
.B(n_116),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_70),
.B(n_41),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_117),
.B(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_121),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_120),
.B(n_132),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g180 ( 
.A(n_133),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_69),
.B(n_75),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_142),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_77),
.A2(n_63),
.B1(n_52),
.B2(n_44),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_154),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_77),
.A2(n_63),
.B1(n_44),
.B2(n_51),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_51),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_6),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_82),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_143),
.A2(n_145),
.B1(n_116),
.B2(n_131),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_8),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_93),
.A2(n_9),
.B1(n_2),
.B2(n_4),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_150),
.Y(n_200)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_9),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_0),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_78),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_67),
.B(n_4),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_159),
.B(n_120),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_68),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_0),
.B1(n_159),
.B2(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_5),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_162),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_83),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_83),
.B(n_11),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_165),
.Y(n_209)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_93),
.A2(n_0),
.A3(n_12),
.B1(n_13),
.B2(n_103),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_174),
.B(n_177),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_90),
.C(n_112),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_191),
.C(n_204),
.Y(n_239)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_178),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_114),
.B1(n_108),
.B2(n_80),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_169),
.A2(n_173),
.B1(n_167),
.B2(n_177),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_135),
.B(n_72),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_173),
.B(n_182),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_0),
.B(n_71),
.Y(n_174)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_130),
.B(n_71),
.Y(n_177)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_197),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_104),
.A3(n_107),
.B1(n_66),
.B2(n_0),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_189),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_66),
.C(n_104),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_150),
.B1(n_141),
.B2(n_155),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

INVx6_ASAP7_75t_SL g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_153),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_149),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_128),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_151),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_147),
.A2(n_148),
.B1(n_164),
.B2(n_115),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_176),
.B(n_172),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_128),
.B(n_160),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_127),
.B(n_133),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_159),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_121),
.B(n_140),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_127),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_246),
.C(n_196),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_213),
.B(n_239),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_216),
.B(n_234),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_248),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_154),
.B1(n_129),
.B2(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_218),
.A2(n_220),
.B1(n_243),
.B2(n_197),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_149),
.B(n_129),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_219),
.A2(n_242),
.B(n_180),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_186),
.A2(n_155),
.B1(n_141),
.B2(n_146),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_244),
.B1(n_183),
.B2(n_178),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_229),
.B(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_119),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_233),
.C(n_214),
.Y(n_284)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_169),
.B1(n_166),
.B2(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_188),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_238),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_190),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_190),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_245),
.B1(n_250),
.B2(n_223),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_169),
.A2(n_170),
.B1(n_199),
.B2(n_193),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_169),
.A2(n_170),
.B1(n_205),
.B2(n_209),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_182),
.B1(n_205),
.B2(n_181),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_181),
.C(n_203),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_185),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_202),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_172),
.A2(n_187),
.B1(n_198),
.B2(n_179),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_171),
.C(n_168),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_207),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_261),
.B(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_214),
.B(n_221),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_263),
.C(n_284),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_258),
.B(n_270),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_273),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_180),
.C(n_228),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_180),
.B1(n_244),
.B2(n_231),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_271),
.B1(n_276),
.B2(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_180),
.B1(n_226),
.B2(n_223),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_217),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_278),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_235),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_222),
.Y(n_274)
);

HAxp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_275),
.CON(n_287),
.SN(n_287)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_224),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_232),
.B1(n_213),
.B2(n_215),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_245),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_233),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_279),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_218),
.A2(n_225),
.B1(n_246),
.B2(n_212),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_220),
.A2(n_242),
.B1(n_229),
.B2(n_240),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_282),
.A2(n_283),
.B1(n_256),
.B2(n_258),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_250),
.A2(n_216),
.B1(n_236),
.B2(n_238),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_293),
.B1(n_297),
.B2(n_308),
.Y(n_329)
);

NOR4xp25_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_249),
.C(n_278),
.D(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_296),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_252),
.B(n_266),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_262),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_260),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_263),
.C(n_284),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_295),
.C(n_303),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_255),
.C(n_281),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_260),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_265),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_304),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_268),
.B(n_254),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_257),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_256),
.A2(n_266),
.B1(n_259),
.B2(n_271),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_308),
.A2(n_311),
.B1(n_261),
.B2(n_280),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_302),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_299),
.B1(n_307),
.B2(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_252),
.A2(n_273),
.B1(n_270),
.B2(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_315),
.A2(n_322),
.B1(n_285),
.B2(n_310),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_269),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_295),
.C(n_303),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_318),
.B(n_292),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_319),
.B(n_321),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_290),
.A2(n_296),
.B1(n_304),
.B2(n_300),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_325),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_309),
.B(n_306),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_289),
.B1(n_286),
.B2(n_287),
.Y(n_342)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

OAI221xp5_ASAP7_75t_L g344 ( 
.A1(n_330),
.A2(n_331),
.B1(n_319),
.B2(n_323),
.C(n_322),
.Y(n_344)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_288),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_338),
.Y(n_357)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_337),
.A2(n_327),
.B(n_347),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_288),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_341),
.C(n_345),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_293),
.C(n_299),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_342),
.B(n_343),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_289),
.A3(n_317),
.B1(n_331),
.B2(n_320),
.C1(n_315),
.C2(n_323),
.Y(n_343)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_312),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_335),
.A2(n_318),
.B(n_346),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_349),
.B(n_347),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_314),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_353),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_313),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_330),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_356),
.Y(n_364)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

AOI221xp5_ASAP7_75t_L g361 ( 
.A1(n_358),
.A2(n_334),
.B1(n_335),
.B2(n_341),
.C(n_340),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_354),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_336),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_360),
.B(n_361),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_339),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_355),
.C(n_357),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_365),
.A2(n_367),
.B1(n_364),
.B2(n_348),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_358),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_368),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_366),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_372),
.C(n_357),
.Y(n_373)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_360),
.A3(n_350),
.B1(n_354),
.B2(n_349),
.C1(n_340),
.C2(n_361),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_333),
.B(n_338),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_353),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);


endmodule