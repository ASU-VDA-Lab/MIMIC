module fake_jpeg_1495_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_73),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_60),
.B1(n_57),
.B2(n_58),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_67),
.B(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_59),
.C(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_56),
.B1(n_60),
.B2(n_48),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_89),
.B1(n_49),
.B2(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_58),
.B1(n_66),
.B2(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_2),
.Y(n_104)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_53),
.B1(n_52),
.B2(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_101),
.B1(n_85),
.B2(n_5),
.Y(n_110)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_107),
.Y(n_111)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_3),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_20),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_105),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_22),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_4),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_6),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_26),
.C(n_45),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_118),
.B1(n_111),
.B2(n_110),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_131),
.B(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_91),
.B1(n_99),
.B2(n_28),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_135),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_99),
.B(n_7),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_12),
.B(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_6),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_29),
.B1(n_43),
.B2(n_42),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_8),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_10),
.C(n_11),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_46),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_11),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_8),
.B(n_9),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_10),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_157),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_37),
.C(n_36),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_166),
.C(n_161),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_32),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_160),
.B(n_140),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.C(n_143),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_15),
.C(n_16),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_171),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_129),
.B1(n_136),
.B2(n_133),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_131),
.B1(n_173),
.B2(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_151),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_142),
.C(n_134),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_136),
.B1(n_165),
.B2(n_153),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_163),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_180),
.B(n_160),
.C(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_179),
.B(n_171),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_183),
.A2(n_185),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_187),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_177),
.C(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_184),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_146),
.Y(n_191)
);


endmodule