module fake_jpeg_17902_n_358 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

CKINVDCx11_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_54),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_40),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_38),
.B1(n_34),
.B2(n_30),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_36),
.B1(n_39),
.B2(n_20),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_30),
.B1(n_38),
.B2(n_34),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_38),
.B1(n_34),
.B2(n_30),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_73),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_29),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_70),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_54),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_71),
.C(n_31),
.Y(n_131)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_19),
.Y(n_92)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_36),
.B1(n_19),
.B2(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_36),
.B1(n_19),
.B2(n_49),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_104),
.B1(n_107),
.B2(n_27),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_55),
.B1(n_53),
.B2(n_44),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_29),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_110),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_0),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_109),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_26),
.CON(n_107),
.SN(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_23),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_27),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_89),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_33),
.B(n_35),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_48),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_131),
.C(n_109),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_83),
.B(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_74),
.B1(n_69),
.B2(n_60),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_93),
.B1(n_112),
.B2(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_83),
.B(n_71),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_88),
.B(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_104),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_74),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_69),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_60),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_95),
.B(n_84),
.C(n_111),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_144),
.A2(n_171),
.B(n_114),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_104),
.B1(n_113),
.B2(n_108),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_133),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_152),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_160),
.Y(n_186)
);

CKINVDCx12_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_156),
.B1(n_115),
.B2(n_137),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_132),
.B(n_130),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_132),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_120),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_113),
.C(n_98),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_63),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_167),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_93),
.C(n_78),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_78),
.C(n_105),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_103),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_78),
.C(n_105),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_169),
.C(n_141),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_101),
.C(n_99),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_33),
.B(n_28),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_72),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_143),
.B(n_139),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_177),
.A2(n_178),
.B(n_182),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_121),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_121),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_198),
.C(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_185),
.B(n_189),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_192),
.C(n_199),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_144),
.A2(n_161),
.B1(n_164),
.B2(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_201),
.B1(n_137),
.B2(n_129),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_120),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_119),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_146),
.A2(n_130),
.B1(n_118),
.B2(n_126),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_138),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_79),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_119),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_150),
.B(n_172),
.C(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_230),
.Y(n_241)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_79),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_130),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_212),
.C(n_218),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_148),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_135),
.C(n_17),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_213),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_127),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_129),
.Y(n_219)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_103),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_177),
.C(n_174),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_173),
.B1(n_99),
.B2(n_32),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_33),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_184),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_25),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_0),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_1),
.B(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_35),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_35),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_232),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_35),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_188),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_236),
.A2(n_255),
.B(n_256),
.Y(n_277)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_204),
.B1(n_182),
.B2(n_199),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_242),
.A2(n_228),
.B1(n_209),
.B2(n_234),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_196),
.B1(n_193),
.B2(n_182),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_249),
.B1(n_250),
.B2(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_208),
.B(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_248),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_173),
.B1(n_176),
.B2(n_101),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_257),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_32),
.B(n_25),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_32),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_230),
.B1(n_210),
.B2(n_216),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_258),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_237),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_215),
.C(n_212),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_273),
.C(n_276),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_215),
.C(n_218),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_220),
.C(n_211),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_217),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_257),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_226),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_283),
.C(n_276),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_282),
.A2(n_241),
.B1(n_252),
.B2(n_250),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_234),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_207),
.B(n_236),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_288),
.A2(n_275),
.B(n_243),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_241),
.B1(n_238),
.B2(n_228),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_255),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_259),
.C(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_252),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_249),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_205),
.B1(n_229),
.B2(n_225),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_259),
.C(n_238),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_280),
.C(n_264),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_240),
.C(n_256),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_299),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_274),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_267),
.B1(n_271),
.B2(n_205),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_309),
.B(n_316),
.Y(n_319)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_278),
.B(n_264),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_285),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_317),
.C(n_285),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_277),
.B(n_274),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_314),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_277),
.B1(n_282),
.B2(n_281),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_298),
.B1(n_286),
.B2(n_293),
.Y(n_320)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_255),
.A3(n_229),
.B1(n_261),
.B2(n_6),
.C(n_7),
.Y(n_316)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_306),
.A2(n_296),
.B(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_322),
.B(n_323),
.Y(n_331)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_306),
.A2(n_11),
.B(n_17),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_313),
.A2(n_312),
.B(n_304),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_10),
.B(n_16),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_311),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_1),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_305),
.B(n_310),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_308),
.B1(n_302),
.B2(n_37),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_328),
.C(n_318),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_308),
.Y(n_333)
);

AOI31xp67_ASAP7_75t_SL g344 ( 
.A1(n_333),
.A2(n_324),
.A3(n_326),
.B(n_6),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_336),
.A2(n_337),
.B(n_338),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_10),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_331),
.B(n_320),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_340),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_342),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_323),
.C(n_322),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_346),
.Y(n_350)
);

AOI211xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_332),
.B(n_5),
.C(n_6),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_37),
.C(n_28),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_347),
.B(n_336),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_345),
.Y(n_351)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_351),
.A2(n_352),
.A3(n_339),
.B1(n_350),
.B2(n_349),
.C1(n_12),
.C2(n_13),
.Y(n_353)
);

OAI311xp33_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_8),
.A3(n_9),
.B1(n_13),
.C1(n_16),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_28),
.C(n_8),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_355),
.A2(n_8),
.B(n_13),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_4),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_4),
.B(n_337),
.Y(n_358)
);


endmodule