module fake_jpeg_30671_n_205 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_31),
.B(n_11),
.Y(n_80)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_16),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_15),
.B1(n_23),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_71),
.B1(n_82),
.B2(n_22),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_0),
.B(n_1),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_19),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_17),
.B1(n_25),
.B2(n_20),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_22),
.B1(n_29),
.B2(n_6),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_32),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_23),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_17),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_75),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_19),
.B1(n_24),
.B2(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_9),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_11),
.A3(n_10),
.B1(n_29),
.B2(n_22),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_85),
.C(n_72),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_22),
.B1(n_29),
.B2(n_8),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_22),
.B1(n_29),
.B2(n_8),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_29),
.C(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_98),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_50),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_48),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_82),
.B1(n_79),
.B2(n_51),
.Y(n_105)
);

AOI22x1_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_78),
.B1(n_64),
.B2(n_50),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_107),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_53),
.B(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_70),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_85),
.B(n_51),
.C(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_90),
.B1(n_92),
.B2(n_103),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_70),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_64),
.B1(n_76),
.B2(n_105),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_93),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_108),
.B1(n_100),
.B2(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_139),
.B1(n_142),
.B2(n_149),
.Y(n_160)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_108),
.B1(n_100),
.B2(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_97),
.B1(n_76),
.B2(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_113),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_156),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_110),
.B(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_162),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_131),
.B(n_123),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_127),
.Y(n_162)
);

NOR4xp25_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_121),
.C(n_119),
.D(n_112),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_135),
.B1(n_112),
.B2(n_138),
.C(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_111),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_139),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_169),
.C(n_172),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_151),
.C(n_146),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_163),
.C(n_122),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_138),
.C(n_150),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_112),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_137),
.C(n_152),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_164),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_122),
.B1(n_140),
.B2(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_157),
.B1(n_172),
.B2(n_169),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_174),
.B1(n_137),
.B2(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_161),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g186 ( 
.A1(n_183),
.A2(n_184),
.B(n_170),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_134),
.B1(n_128),
.B2(n_113),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_182),
.B1(n_180),
.B2(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_179),
.B(n_185),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_202),
.B(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_197),
.C(n_192),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_188),
.Y(n_205)
);


endmodule