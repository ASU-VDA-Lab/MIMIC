module real_aes_10701_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_269;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_0), .Y(n_1222) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1), .Y(n_1348) );
AOI21xp33_ASAP7_75t_L g648 ( .A1(n_2), .A2(n_318), .B(n_506), .Y(n_648) );
INVx1_ASAP7_75t_L g685 ( .A(n_2), .Y(n_685) );
INVx1_ASAP7_75t_L g335 ( .A(n_3), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_3), .A2(n_79), .B1(n_419), .B2(n_425), .C(n_429), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_4), .A2(n_263), .B1(n_318), .B2(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g449 ( .A(n_4), .Y(n_449) );
XOR2xp5_ASAP7_75t_L g1587 ( .A(n_5), .B(n_1588), .Y(n_1587) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_6), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_6), .B(n_200), .Y(n_381) );
AND2x2_ASAP7_75t_L g398 ( .A(n_6), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g462 ( .A(n_6), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_7), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_8), .A2(n_157), .B1(n_349), .B2(n_483), .C(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g527 ( .A(n_8), .Y(n_527) );
INVxp67_ASAP7_75t_L g995 ( .A(n_9), .Y(n_995) );
OAI222xp33_ASAP7_75t_L g1010 ( .A1(n_9), .A2(n_45), .B1(n_255), .B2(n_739), .C1(n_1011), .C2(n_1013), .Y(n_1010) );
OAI211xp5_ASAP7_75t_L g1213 ( .A1(n_10), .A2(n_1214), .B(n_1215), .C(n_1242), .Y(n_1213) );
OAI221xp5_ASAP7_75t_L g846 ( .A1(n_11), .A2(n_847), .B1(n_849), .B2(n_855), .C(n_862), .Y(n_846) );
INVx1_ASAP7_75t_L g889 ( .A(n_11), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_12), .Y(n_1229) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_13), .A2(n_57), .B1(n_402), .B2(n_838), .C(n_839), .Y(n_837) );
INVx1_ASAP7_75t_L g904 ( .A(n_13), .Y(n_904) );
INVx1_ASAP7_75t_L g828 ( .A(n_14), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_14), .A2(n_58), .B1(n_371), .B2(n_629), .Y(n_891) );
AO22x2_ASAP7_75t_L g911 ( .A1(n_15), .A2(n_912), .B1(n_969), .B2(n_970), .Y(n_911) );
CKINVDCx14_ASAP7_75t_R g969 ( .A(n_15), .Y(n_969) );
INVx1_ASAP7_75t_L g1128 ( .A(n_16), .Y(n_1128) );
INVx1_ASAP7_75t_L g1382 ( .A(n_17), .Y(n_1382) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_18), .A2(n_39), .B1(n_347), .B2(n_348), .C(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g455 ( .A(n_18), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_19), .A2(n_253), .B1(n_562), .B2(n_772), .C(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g797 ( .A(n_19), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_20), .Y(n_1174) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_21), .A2(n_559), .B1(n_624), .B2(n_631), .C(n_638), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_21), .A2(n_179), .B1(n_659), .B2(n_671), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g857 ( .A(n_22), .Y(n_857) );
AO221x2_ASAP7_75t_L g1319 ( .A1(n_23), .A2(n_59), .B1(n_1303), .B2(n_1312), .C(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1158 ( .A(n_24), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_24), .A2(n_224), .B1(n_775), .B2(n_1196), .Y(n_1195) );
INVx2_ASAP7_75t_L g326 ( .A(n_25), .Y(n_326) );
OR2x2_ASAP7_75t_L g344 ( .A(n_25), .B(n_331), .Y(n_344) );
AO22x1_ASAP7_75t_L g819 ( .A1(n_26), .A2(n_820), .B1(n_909), .B2(n_910), .Y(n_819) );
INVx1_ASAP7_75t_L g910 ( .A(n_26), .Y(n_910) );
INVx1_ASAP7_75t_L g1336 ( .A(n_27), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_28), .A2(n_234), .B1(n_577), .B2(n_579), .Y(n_576) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_28), .A2(n_234), .B1(n_425), .B2(n_429), .C(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g998 ( .A(n_29), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_30), .A2(n_106), .B1(n_323), .B2(n_1039), .C(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1066 ( .A(n_30), .Y(n_1066) );
BUFx2_ASAP7_75t_L g375 ( .A(n_31), .Y(n_375) );
OR2x2_ASAP7_75t_L g380 ( .A(n_31), .B(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g384 ( .A(n_31), .Y(n_384) );
INVx1_ASAP7_75t_L g397 ( .A(n_31), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_32), .A2(n_210), .B1(n_593), .B2(n_979), .C(n_1072), .Y(n_1223) );
INVx1_ASAP7_75t_L g1257 ( .A(n_32), .Y(n_1257) );
INVx1_ASAP7_75t_L g547 ( .A(n_33), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g1543 ( .A1(n_34), .A2(n_175), .B1(n_1544), .B2(n_1545), .Y(n_1543) );
INVx1_ASAP7_75t_L g1570 ( .A(n_34), .Y(n_1570) );
INVx1_ASAP7_75t_L g915 ( .A(n_35), .Y(n_915) );
AOI21xp33_ASAP7_75t_L g958 ( .A1(n_35), .A2(n_371), .B(n_959), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_36), .A2(n_161), .B1(n_563), .B2(n_1049), .C(n_1051), .Y(n_1048) );
INVx1_ASAP7_75t_L g1077 ( .A(n_36), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_37), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1169 ( .A(n_38), .Y(n_1169) );
INVx1_ASAP7_75t_L g440 ( .A(n_39), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_40), .Y(n_359) );
INVx1_ASAP7_75t_L g1288 ( .A(n_41), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_41), .B(n_1286), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_42), .A2(n_141), .B1(n_371), .B2(n_629), .Y(n_647) );
INVx1_ASAP7_75t_L g686 ( .A(n_42), .Y(n_686) );
INVx1_ASAP7_75t_L g984 ( .A(n_43), .Y(n_984) );
INVx1_ASAP7_75t_L g1129 ( .A(n_44), .Y(n_1129) );
INVxp67_ASAP7_75t_L g993 ( .A(n_45), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_46), .A2(n_204), .B1(n_486), .B2(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g598 ( .A(n_46), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_47), .A2(n_108), .B1(n_721), .B2(n_722), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_47), .A2(n_71), .B1(n_637), .B2(n_750), .C(n_752), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_48), .A2(n_216), .B1(n_961), .B2(n_962), .C(n_964), .Y(n_960) );
INVx1_ASAP7_75t_L g967 ( .A(n_48), .Y(n_967) );
CKINVDCx16_ASAP7_75t_R g1333 ( .A(n_49), .Y(n_1333) );
INVx1_ASAP7_75t_L g854 ( .A(n_50), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_50), .A2(n_149), .B1(n_484), .B2(n_629), .Y(n_885) );
INVx1_ASAP7_75t_L g1377 ( .A(n_51), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_52), .A2(n_162), .B1(n_841), .B2(n_845), .Y(n_840) );
OAI22xp5_ASAP7_75t_SL g873 ( .A1(n_52), .A2(n_162), .B1(n_874), .B2(n_878), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g1044 ( .A(n_53), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_54), .A2(n_1213), .B1(n_1270), .B2(n_1271), .Y(n_1212) );
INVx1_ASAP7_75t_L g1271 ( .A(n_54), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1540 ( .A1(n_55), .A2(n_80), .B1(n_307), .B2(n_1541), .Y(n_1540) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_55), .A2(n_80), .B1(n_1154), .B2(n_1155), .Y(n_1547) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_56), .A2(n_179), .B1(n_361), .B2(n_367), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_56), .A2(n_260), .B1(n_662), .B2(n_667), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_57), .A2(n_115), .B1(n_906), .B2(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g830 ( .A(n_58), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_60), .A2(n_72), .B1(n_347), .B2(n_562), .C(n_563), .Y(n_561) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_60), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_61), .Y(n_501) );
INVx1_ASAP7_75t_L g1108 ( .A(n_62), .Y(n_1108) );
AO22x2_ASAP7_75t_L g1149 ( .A1(n_63), .A2(n_1150), .B1(n_1151), .B2(n_1207), .Y(n_1149) );
INVx1_ASAP7_75t_L g1207 ( .A(n_63), .Y(n_1207) );
CKINVDCx16_ASAP7_75t_R g1295 ( .A(n_64), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_65), .A2(n_150), .B1(n_1531), .B2(n_1532), .Y(n_1530) );
INVxp67_ASAP7_75t_SL g1555 ( .A(n_65), .Y(n_1555) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_66), .A2(n_211), .B1(n_520), .B2(n_979), .C(n_1072), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_66), .A2(n_211), .B1(n_962), .B2(n_1135), .Y(n_1134) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_67), .Y(n_1176) );
INVxp67_ASAP7_75t_L g1121 ( .A(n_68), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_68), .A2(n_126), .B1(n_1054), .B2(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1221 ( .A(n_69), .Y(n_1221) );
AOI221xp5_ASAP7_75t_L g1264 ( .A1(n_69), .A2(n_133), .B1(n_755), .B2(n_1265), .C(n_1267), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_70), .A2(n_185), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
INVx1_ASAP7_75t_L g1064 ( .A(n_70), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_71), .A2(n_130), .B1(n_715), .B2(n_718), .Y(n_714) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_72), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_73), .A2(n_194), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
AOI22xp33_ASAP7_75t_SL g1200 ( .A1(n_73), .A2(n_194), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_74), .Y(n_1167) );
INVx1_ASAP7_75t_L g1237 ( .A(n_75), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_75), .A2(n_237), .B1(n_361), .B2(n_367), .Y(n_1269) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_76), .A2(n_91), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g748 ( .A(n_76), .Y(n_748) );
INVx1_ASAP7_75t_L g1349 ( .A(n_77), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_78), .A2(n_231), .B1(n_569), .B2(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g798 ( .A(n_78), .Y(n_798) );
INVx1_ASAP7_75t_L g339 ( .A(n_79), .Y(n_339) );
INVx1_ASAP7_75t_L g709 ( .A(n_81), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_81), .A2(n_104), .B1(n_738), .B2(n_740), .C(n_741), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_82), .A2(n_152), .B1(n_772), .B2(n_773), .C(n_1025), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_82), .A2(n_169), .B1(n_1028), .B2(n_1029), .C(n_1031), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_83), .Y(n_1178) );
CKINVDCx16_ASAP7_75t_R g1301 ( .A(n_84), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1317 ( .A1(n_85), .A2(n_146), .B1(n_1306), .B2(n_1309), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_86), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_87), .A2(n_208), .B1(n_722), .B2(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g765 ( .A(n_87), .Y(n_765) );
INVx1_ASAP7_75t_L g327 ( .A(n_88), .Y(n_327) );
INVx1_ASAP7_75t_L g331 ( .A(n_88), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_89), .A2(n_247), .B1(n_486), .B2(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g538 ( .A(n_89), .Y(n_538) );
INVx1_ASAP7_75t_L g556 ( .A(n_90), .Y(n_556) );
INVx1_ASAP7_75t_L g764 ( .A(n_91), .Y(n_764) );
INVx1_ASAP7_75t_L g1536 ( .A(n_92), .Y(n_1536) );
OAI221xp5_ASAP7_75t_L g1548 ( .A1(n_92), .A2(n_847), .B1(n_1549), .B2(n_1552), .C(n_1557), .Y(n_1548) );
INVx1_ASAP7_75t_L g632 ( .A(n_93), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_93), .A2(n_159), .B1(n_658), .B2(n_659), .Y(n_657) );
NAND2xp33_ASAP7_75t_SL g312 ( .A(n_94), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g400 ( .A(n_94), .Y(n_400) );
INVx1_ASAP7_75t_L g1561 ( .A(n_95), .Y(n_1561) );
OAI22xp5_ASAP7_75t_L g1572 ( .A1(n_95), .A2(n_121), .B1(n_906), .B2(n_907), .Y(n_1572) );
OAI221xp5_ASAP7_75t_L g1164 ( .A1(n_96), .A2(n_823), .B1(n_1165), .B2(n_1171), .C(n_1175), .Y(n_1164) );
AOI22xp33_ASAP7_75t_SL g1199 ( .A1(n_96), .A2(n_128), .B1(n_755), .B2(n_1039), .Y(n_1199) );
INVx1_ASAP7_75t_L g695 ( .A(n_97), .Y(n_695) );
XNOR2xp5_ASAP7_75t_L g974 ( .A(n_98), .B(n_975), .Y(n_974) );
INVxp67_ASAP7_75t_L g1116 ( .A(n_99), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1141 ( .A1(n_99), .A2(n_120), .B1(n_637), .B2(n_1142), .C(n_1144), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_100), .A2(n_620), .B1(n_690), .B2(n_691), .Y(n_619) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_100), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_101), .Y(n_788) );
INVxp67_ASAP7_75t_L g982 ( .A(n_102), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_102), .A2(n_167), .B1(n_347), .B2(n_348), .C(n_563), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_103), .Y(n_297) );
INVx1_ASAP7_75t_L g705 ( .A(n_104), .Y(n_705) );
INVx1_ASAP7_75t_L g1335 ( .A(n_105), .Y(n_1335) );
INVx1_ASAP7_75t_L g1068 ( .A(n_106), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_107), .A2(n_218), .B1(n_562), .B2(n_637), .C(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g806 ( .A(n_107), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_108), .A2(n_130), .B1(n_755), .B2(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g1235 ( .A(n_109), .Y(n_1235) );
OAI211xp5_ASAP7_75t_L g1254 ( .A1(n_109), .A2(n_1255), .B(n_1256), .C(n_1261), .Y(n_1254) );
INVx1_ASAP7_75t_L g1241 ( .A(n_110), .Y(n_1241) );
OAI211xp5_ASAP7_75t_SL g1243 ( .A1(n_110), .A2(n_1244), .B(n_1245), .C(n_1253), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1562 ( .A1(n_111), .A2(n_121), .B1(n_728), .B2(n_1563), .C(n_1565), .Y(n_1562) );
OAI22xp5_ASAP7_75t_L g1573 ( .A1(n_111), .A2(n_197), .B1(n_1574), .B2(n_1576), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_112), .A2(n_226), .B1(n_573), .B2(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g591 ( .A(n_112), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_113), .Y(n_369) );
AO221x2_ASAP7_75t_L g1346 ( .A1(n_114), .A2(n_187), .B1(n_1297), .B2(n_1303), .C(n_1347), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_115), .A2(n_127), .B1(n_834), .B2(n_835), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_116), .A2(n_209), .B1(n_318), .B2(n_506), .C(n_562), .Y(n_571) );
INVx1_ASAP7_75t_L g590 ( .A(n_116), .Y(n_590) );
INVxp33_ASAP7_75t_L g1104 ( .A(n_117), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_117), .A2(n_148), .B1(n_775), .B2(n_1137), .C(n_1139), .Y(n_1136) );
INVx1_ASAP7_75t_L g1163 ( .A(n_118), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_118), .A2(n_135), .B1(n_1051), .B2(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g272 ( .A(n_119), .Y(n_272) );
INVxp67_ASAP7_75t_L g1118 ( .A(n_120), .Y(n_1118) );
INVx1_ASAP7_75t_L g376 ( .A(n_122), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_123), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_124), .Y(n_923) );
OA22x2_ASAP7_75t_L g766 ( .A1(n_125), .A2(n_767), .B1(n_812), .B2(n_813), .Y(n_766) );
INVx1_ASAP7_75t_L g813 ( .A(n_125), .Y(n_813) );
INVx1_ASAP7_75t_L g1113 ( .A(n_126), .Y(n_1113) );
INVx1_ASAP7_75t_L g902 ( .A(n_127), .Y(n_902) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_128), .A2(n_847), .B1(n_862), .B2(n_1157), .C(n_1161), .Y(n_1156) );
INVx1_ASAP7_75t_L g1106 ( .A(n_129), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_131), .A2(n_178), .B1(n_1303), .B2(n_1312), .Y(n_1318) );
AOI22xp33_ASAP7_75t_SL g302 ( .A1(n_132), .A2(n_214), .B1(n_303), .B2(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g411 ( .A(n_132), .Y(n_411) );
INVx1_ASAP7_75t_L g1219 ( .A(n_133), .Y(n_1219) );
OAI222xp33_ASAP7_75t_L g977 ( .A1(n_134), .A2(n_168), .B1(n_258), .B2(n_379), .C1(n_978), .C2(n_979), .Y(n_977) );
INVx1_ASAP7_75t_L g1004 ( .A(n_134), .Y(n_1004) );
INVx1_ASAP7_75t_L g1162 ( .A(n_135), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_136), .Y(n_508) );
INVx1_ASAP7_75t_L g1321 ( .A(n_137), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_138), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g1518 ( .A(n_139), .Y(n_1518) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_140), .A2(n_264), .B1(n_483), .B2(n_505), .C(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g515 ( .A(n_140), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_141), .A2(n_249), .B1(n_688), .B2(n_689), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_142), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_143), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_144), .Y(n_789) );
INVx1_ASAP7_75t_L g730 ( .A(n_145), .Y(n_730) );
INVx1_ASAP7_75t_L g495 ( .A(n_147), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_147), .A2(n_227), .B1(n_426), .B2(n_520), .C(n_522), .Y(n_519) );
INVxp33_ASAP7_75t_L g1109 ( .A(n_148), .Y(n_1109) );
INVx1_ASAP7_75t_L g852 ( .A(n_149), .Y(n_852) );
INVxp67_ASAP7_75t_SL g1556 ( .A(n_150), .Y(n_1556) );
INVx1_ASAP7_75t_L g1539 ( .A(n_151), .Y(n_1539) );
OAI211xp5_ASAP7_75t_SL g1558 ( .A1(n_151), .A2(n_823), .B(n_1559), .C(n_1566), .Y(n_1558) );
OAI332xp33_ASAP7_75t_L g980 ( .A1(n_152), .A2(n_432), .A3(n_615), .B1(n_936), .B2(n_981), .B3(n_985), .C1(n_988), .C2(n_994), .Y(n_980) );
INVx1_ASAP7_75t_L g916 ( .A(n_153), .Y(n_916) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_153), .A2(n_196), .B1(n_629), .B2(n_957), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_154), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_155), .Y(n_481) );
INVx1_ASAP7_75t_L g560 ( .A(n_156), .Y(n_560) );
INVx1_ASAP7_75t_L g533 ( .A(n_157), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g1324 ( .A1(n_158), .A2(n_173), .B1(n_1306), .B2(n_1309), .Y(n_1324) );
INVx1_ASAP7_75t_L g627 ( .A(n_159), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_160), .Y(n_1181) );
INVx1_ASAP7_75t_L g1079 ( .A(n_161), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g1233 ( .A(n_163), .Y(n_1233) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_163), .A2(n_195), .B1(n_1250), .B2(n_1251), .C(n_1252), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_164), .A2(n_212), .B1(n_379), .B2(n_688), .Y(n_937) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_164), .A2(n_191), .B1(n_371), .B2(n_629), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_165), .A2(n_191), .B1(n_935), .B2(n_936), .Y(n_934) );
INVx1_ASAP7_75t_L g947 ( .A(n_165), .Y(n_947) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_166), .A2(n_484), .B(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_166), .A2(n_248), .B1(n_662), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g986 ( .A(n_167), .Y(n_986) );
INVx1_ASAP7_75t_L g1020 ( .A(n_168), .Y(n_1020) );
INVx1_ASAP7_75t_L g1023 ( .A(n_169), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_170), .Y(n_924) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_171), .B(n_272), .Y(n_1284) );
AND3x2_ASAP7_75t_L g1300 ( .A(n_171), .B(n_272), .C(n_1287), .Y(n_1300) );
OA332x1_ASAP7_75t_L g913 ( .A1(n_172), .A2(n_432), .A3(n_914), .B1(n_919), .B2(n_922), .B3(n_925), .C1(n_930), .C2(n_931), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g952 ( .A1(n_172), .A2(n_506), .B(n_953), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g1325 ( .A1(n_174), .A2(n_206), .B1(n_1297), .B2(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1569 ( .A(n_175), .Y(n_1569) );
INVx2_ASAP7_75t_L g285 ( .A(n_176), .Y(n_285) );
INVx1_ASAP7_75t_L g580 ( .A(n_177), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_180), .A2(n_240), .B1(n_772), .B2(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g803 ( .A(n_180), .Y(n_803) );
INVx1_ASAP7_75t_L g1126 ( .A(n_181), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_182), .Y(n_786) );
OAI211xp5_ASAP7_75t_L g822 ( .A1(n_183), .A2(n_823), .B(n_827), .C(n_832), .Y(n_822) );
INVx1_ASAP7_75t_L g890 ( .A(n_183), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_184), .A2(n_220), .B1(n_942), .B2(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1075 ( .A(n_184), .Y(n_1075) );
INVx1_ASAP7_75t_L g1069 ( .A(n_185), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_186), .A2(n_190), .B1(n_1303), .B2(n_1312), .Y(n_1311) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_188), .Y(n_642) );
INVx1_ASAP7_75t_L g1287 ( .A(n_189), .Y(n_1287) );
CKINVDCx16_ASAP7_75t_R g1332 ( .A(n_192), .Y(n_1332) );
INVx1_ASAP7_75t_L g1379 ( .A(n_193), .Y(n_1379) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_195), .Y(n_1226) );
INVx1_ASAP7_75t_L g920 ( .A(n_196), .Y(n_920) );
INVx1_ASAP7_75t_L g1560 ( .A(n_197), .Y(n_1560) );
OAI22xp33_ASAP7_75t_L g1045 ( .A1(n_198), .A2(n_199), .B1(n_962), .B2(n_1046), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_198), .A2(n_199), .B1(n_520), .B2(n_979), .C(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g287 ( .A(n_200), .Y(n_287) );
INVx2_ASAP7_75t_L g399 ( .A(n_200), .Y(n_399) );
OR2x2_ASAP7_75t_L g621 ( .A(n_201), .B(n_378), .Y(n_621) );
INVx1_ASAP7_75t_L g1124 ( .A(n_202), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_203), .A2(n_238), .B1(n_1306), .B2(n_1309), .Y(n_1305) );
INVx1_ASAP7_75t_L g608 ( .A(n_204), .Y(n_608) );
INVx1_ASAP7_75t_L g866 ( .A(n_205), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_207), .A2(n_551), .B1(n_617), .B2(n_618), .Y(n_550) );
INVx1_ASAP7_75t_L g618 ( .A(n_207), .Y(n_618) );
INVx1_ASAP7_75t_L g733 ( .A(n_208), .Y(n_733) );
INVx1_ASAP7_75t_L g586 ( .A(n_209), .Y(n_586) );
INVx1_ASAP7_75t_L g1260 ( .A(n_210), .Y(n_1260) );
INVx1_ASAP7_75t_L g965 ( .A(n_212), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_213), .Y(n_492) );
INVx1_ASAP7_75t_L g389 ( .A(n_214), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_215), .Y(n_493) );
INVx1_ASAP7_75t_L g968 ( .A(n_216), .Y(n_968) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_217), .Y(n_365) );
INVx1_ASAP7_75t_L g804 ( .A(n_218), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_219), .Y(n_776) );
INVx1_ASAP7_75t_L g1081 ( .A(n_220), .Y(n_1081) );
INVx1_ASAP7_75t_L g1059 ( .A(n_221), .Y(n_1059) );
INVx1_ASAP7_75t_L g1231 ( .A(n_222), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_223), .A2(n_229), .B1(n_579), .B2(n_778), .Y(n_777) );
OAI221xp5_ASAP7_75t_L g800 ( .A1(n_223), .A2(n_229), .B1(n_419), .B2(n_425), .C(n_429), .Y(n_800) );
INVx1_ASAP7_75t_L g1160 ( .A(n_224), .Y(n_1160) );
INVx1_ASAP7_75t_L g1289 ( .A(n_225), .Y(n_1289) );
INVx1_ASAP7_75t_L g584 ( .A(n_226), .Y(n_584) );
INVx1_ASAP7_75t_L g496 ( .A(n_227), .Y(n_496) );
INVx1_ASAP7_75t_L g509 ( .A(n_228), .Y(n_509) );
INVx1_ASAP7_75t_L g570 ( .A(n_230), .Y(n_570) );
INVx1_ASAP7_75t_L g794 ( .A(n_231), .Y(n_794) );
INVx1_ASAP7_75t_L g703 ( .A(n_232), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_232), .A2(n_250), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g987 ( .A(n_233), .Y(n_987) );
INVx1_ASAP7_75t_L g1007 ( .A(n_235), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_236), .Y(n_1131) );
INVx1_ASAP7_75t_L g1239 ( .A(n_237), .Y(n_1239) );
INVx1_ASAP7_75t_L g1515 ( .A(n_238), .Y(n_1515) );
AOI22xp33_ASAP7_75t_L g1581 ( .A1(n_238), .A2(n_1582), .B1(n_1586), .B2(n_1590), .Y(n_1581) );
INVx1_ASAP7_75t_L g1148 ( .A(n_239), .Y(n_1148) );
INVx1_ASAP7_75t_L g807 ( .A(n_240), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_241), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_242), .Y(n_860) );
INVx2_ASAP7_75t_L g284 ( .A(n_243), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_244), .Y(n_503) );
INVx1_ASAP7_75t_L g1091 ( .A(n_245), .Y(n_1091) );
AOI21xp33_ASAP7_75t_L g317 ( .A1(n_246), .A2(n_318), .B(n_323), .Y(n_317) );
INVx1_ASAP7_75t_L g406 ( .A(n_246), .Y(n_406) );
INVx1_ASAP7_75t_L g525 ( .A(n_247), .Y(n_525) );
INVx1_ASAP7_75t_L g630 ( .A(n_248), .Y(n_630) );
INVx1_ASAP7_75t_L g645 ( .A(n_249), .Y(n_645) );
INVx1_ASAP7_75t_L g700 ( .A(n_250), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_251), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g1218 ( .A(n_252), .Y(n_1218) );
INVx1_ASAP7_75t_L g795 ( .A(n_253), .Y(n_795) );
INVx1_ASAP7_75t_L g1525 ( .A(n_254), .Y(n_1525) );
INVxp67_ASAP7_75t_L g989 ( .A(n_255), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_256), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_257), .Y(n_706) );
INVx1_ASAP7_75t_L g1008 ( .A(n_258), .Y(n_1008) );
INVx1_ASAP7_75t_L g1529 ( .A(n_259), .Y(n_1529) );
OAI211xp5_ASAP7_75t_SL g639 ( .A1(n_260), .A2(n_640), .B(n_641), .C(n_644), .Y(n_639) );
BUFx3_ASAP7_75t_L g306 ( .A(n_261), .Y(n_306) );
INVx1_ASAP7_75t_L g311 ( .A(n_261), .Y(n_311) );
INVx1_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
BUFx3_ASAP7_75t_L g310 ( .A(n_262), .Y(n_310) );
INVx1_ASAP7_75t_L g444 ( .A(n_263), .Y(n_444) );
INVx1_ASAP7_75t_L g517 ( .A(n_264), .Y(n_517) );
INVx1_ASAP7_75t_L g555 ( .A(n_265), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_288), .B(n_1274), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x4_ASAP7_75t_L g1580 ( .A(n_270), .B(n_276), .Y(n_1580) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_SL g1585 ( .A(n_271), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_271), .B(n_273), .Y(n_1592) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_273), .B(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g656 ( .A(n_279), .B(n_287), .Y(n_656) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g433 ( .A(n_280), .B(n_434), .Y(n_433) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
OR2x2_ASAP7_75t_L g379 ( .A(n_282), .B(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g448 ( .A(n_282), .Y(n_448) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_282), .Y(n_544) );
INVx2_ASAP7_75t_SL g597 ( .A(n_282), .Y(n_597) );
INVx2_ASAP7_75t_SL g859 ( .A(n_282), .Y(n_859) );
INVx1_ASAP7_75t_L g997 ( .A(n_282), .Y(n_997) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x4_ASAP7_75t_L g394 ( .A(n_284), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g404 ( .A(n_284), .Y(n_404) );
AND2x2_ASAP7_75t_L g410 ( .A(n_284), .B(n_285), .Y(n_410) );
INVx2_ASAP7_75t_L g415 ( .A(n_284), .Y(n_415) );
INVx1_ASAP7_75t_L g454 ( .A(n_284), .Y(n_454) );
INVx2_ASAP7_75t_L g395 ( .A(n_285), .Y(n_395) );
INVx1_ASAP7_75t_L g417 ( .A(n_285), .Y(n_417) );
INVx1_ASAP7_75t_L g423 ( .A(n_285), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_285), .B(n_415), .Y(n_439) );
INVx1_ASAP7_75t_L g453 ( .A(n_285), .Y(n_453) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B1(n_1094), .B2(n_1095), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
XNOR2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_692), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B1(n_548), .B2(n_549), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B1(n_471), .B2(n_472), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_386), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_372), .B1(n_376), .B2(n_377), .Y(n_299) );
NAND4xp25_ASAP7_75t_L g300 ( .A(n_301), .B(n_340), .C(n_358), .D(n_368), .Y(n_300) );
AOI322xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_312), .A3(n_317), .B1(n_328), .B2(n_335), .C1(n_336), .C2(n_339), .Y(n_301) );
BUFx3_ASAP7_75t_L g1541 ( .A(n_303), .Y(n_1541) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_304), .Y(n_371) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_304), .Y(n_484) );
BUFx2_ASAP7_75t_L g500 ( .A(n_304), .Y(n_500) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_304), .Y(n_569) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_304), .Y(n_573) );
BUFx2_ASAP7_75t_L g781 ( .A(n_304), .Y(n_781) );
INVx2_ASAP7_75t_SL g899 ( .A(n_304), .Y(n_899) );
HB1xp67_ASAP7_75t_L g1263 ( .A(n_304), .Y(n_1263) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g364 ( .A(n_305), .Y(n_364) );
AND2x2_ASAP7_75t_L g316 ( .A(n_306), .B(n_310), .Y(n_316) );
INVx2_ASAP7_75t_L g321 ( .A(n_306), .Y(n_321) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x6_ASAP7_75t_L g906 ( .A(n_308), .B(n_901), .Y(n_906) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_309), .Y(n_490) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_309), .Y(n_629) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g322 ( .A(n_310), .Y(n_322) );
INVx1_ASAP7_75t_L g363 ( .A(n_311), .Y(n_363) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g562 ( .A(n_314), .Y(n_562) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_315), .Y(n_483) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_315), .Y(n_762) );
INVx1_ASAP7_75t_L g894 ( .A(n_315), .Y(n_894) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
AND2x2_ASAP7_75t_L g903 ( .A(n_318), .B(n_900), .Y(n_903) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g953 ( .A(n_319), .Y(n_953) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g385 ( .A(n_320), .B(n_329), .Y(n_385) );
INVx6_ASAP7_75t_L g488 ( .A(n_320), .Y(n_488) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g338 ( .A(n_321), .Y(n_338) );
INVx1_ASAP7_75t_L g334 ( .A(n_322), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g506 ( .A(n_324), .Y(n_506) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_324), .Y(n_745) );
INVx1_ASAP7_75t_L g773 ( .A(n_324), .Y(n_773) );
AND2x4_ASAP7_75t_L g887 ( .A(n_324), .B(n_384), .Y(n_887) );
INVx2_ASAP7_75t_L g1268 ( .A(n_324), .Y(n_1268) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AND2x4_ASAP7_75t_L g329 ( .A(n_325), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g352 ( .A(n_326), .B(n_327), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_328), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
INVx2_ASAP7_75t_L g735 ( .A(n_328), .Y(n_735) );
INVx2_ASAP7_75t_SL g961 ( .A(n_328), .Y(n_961) );
INVx1_ASAP7_75t_L g1046 ( .A(n_328), .Y(n_1046) );
INVx1_ASAP7_75t_L g1135 ( .A(n_328), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_328), .A2(n_1257), .B1(n_1258), .B2(n_1260), .Y(n_1256) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AND2x4_ASAP7_75t_L g336 ( .A(n_329), .B(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
AND2x2_ASAP7_75t_L g497 ( .A(n_329), .B(n_337), .Y(n_497) );
AND2x4_ASAP7_75t_L g578 ( .A(n_329), .B(n_332), .Y(n_578) );
INVx1_ASAP7_75t_L g761 ( .A(n_329), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g877 ( .A(n_329), .B(n_459), .Y(n_877) );
AND2x2_ASAP7_75t_L g963 ( .A(n_329), .B(n_337), .Y(n_963) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g875 ( .A(n_333), .Y(n_875) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_SL g579 ( .A(n_336), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_336), .A2(n_578), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI222xp33_ASAP7_75t_SL g1001 ( .A1(n_336), .A2(n_1002), .B1(n_1004), .B2(n_1005), .C1(n_1007), .C2(n_1008), .Y(n_1001) );
INVx2_ASAP7_75t_L g879 ( .A(n_337), .Y(n_879) );
BUFx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B1(n_346), .B2(n_353), .C(n_356), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_341), .A2(n_356), .B1(n_481), .B2(n_482), .C(n_485), .Y(n_480) );
INVx2_ASAP7_75t_SL g559 ( .A(n_341), .Y(n_559) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_341), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_341), .A2(n_356), .B1(n_780), .B2(n_782), .C(n_786), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_341), .A2(n_343), .B1(n_356), .B2(n_998), .C(n_1010), .Y(n_1009) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
BUFx4f_ASAP7_75t_L g348 ( .A(n_342), .Y(n_348) );
AND2x4_ASAP7_75t_L g356 ( .A(n_342), .B(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_342), .Y(n_753) );
INVx1_ASAP7_75t_L g1026 ( .A(n_342), .Y(n_1026) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_342), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1052 ( .A(n_342), .Y(n_1052) );
AND2x4_ASAP7_75t_L g370 ( .A(n_343), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g568 ( .A(n_343), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g361 ( .A(n_344), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g367 ( .A(n_344), .B(n_355), .Y(n_367) );
OR2x2_ASAP7_75t_L g901 ( .A(n_344), .B(n_397), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_344), .A2(n_940), .B(n_943), .C(n_944), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_345), .A2(n_359), .B1(n_464), .B2(n_465), .Y(n_463) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_347), .Y(n_1019) );
INVx2_ASAP7_75t_L g1138 ( .A(n_347), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_348), .A2(n_898), .B1(n_924), .B2(n_926), .Y(n_943) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x6_ASAP7_75t_L g1194 ( .A(n_351), .B(n_374), .Y(n_1194) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g564 ( .A(n_352), .Y(n_564) );
INVx2_ASAP7_75t_SL g637 ( .A(n_352), .Y(n_637) );
INVx1_ASAP7_75t_L g882 ( .A(n_352), .Y(n_882) );
INVx1_ASAP7_75t_L g959 ( .A(n_352), .Y(n_959) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g785 ( .A(n_355), .Y(n_785) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_356), .A2(n_558), .B1(n_560), .B2(n_561), .C(n_565), .Y(n_557) );
INVx1_ASAP7_75t_L g638 ( .A(n_356), .Y(n_638) );
INVx1_ASAP7_75t_L g944 ( .A(n_356), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_356), .A2(n_747), .B1(n_1048), .B2(n_1053), .C(n_1055), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_365), .B2(n_366), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_360), .A2(n_366), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_360), .A2(n_366), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_360), .A2(n_366), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_360), .A2(n_366), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_360), .A2(n_366), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_360), .A2(n_366), .B1(n_1128), .B2(n_1129), .Y(n_1147) );
INVx6_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g626 ( .A(n_362), .Y(n_626) );
INVx1_ASAP7_75t_L g744 ( .A(n_362), .Y(n_744) );
INVx1_ASAP7_75t_L g1012 ( .A(n_362), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1524 ( .A(n_362), .Y(n_1524) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g635 ( .A(n_363), .B(n_364), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_365), .A2(n_369), .B1(n_436), .B2(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_370), .B(n_508), .Y(n_507) );
AOI211xp5_ASAP7_75t_SL g732 ( .A1(n_370), .A2(n_733), .B(n_734), .C(n_737), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_370), .A2(n_1038), .B1(n_1041), .B2(n_1044), .C(n_1045), .Y(n_1037) );
AOI211xp5_ASAP7_75t_L g1133 ( .A1(n_370), .A2(n_1124), .B(n_1134), .C(n_1136), .Y(n_1133) );
INVx1_ASAP7_75t_L g1255 ( .A(n_370), .Y(n_1255) );
INVx2_ASAP7_75t_SL g1143 ( .A(n_371), .Y(n_1143) );
BUFx3_ASAP7_75t_L g1201 ( .A(n_371), .Y(n_1201) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_372), .A2(n_377), .B1(n_553), .B2(n_580), .Y(n_552) );
CKINVDCx8_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
OAI31xp33_ASAP7_75t_L g1152 ( .A1(n_373), .A2(n_1153), .A3(n_1156), .B(n_1164), .Y(n_1152) );
BUFx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g652 ( .A(n_374), .Y(n_652) );
AND2x4_ASAP7_75t_L g655 ( .A(n_374), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g674 ( .A(n_374), .B(n_675), .Y(n_674) );
AND2x4_ASAP7_75t_L g713 ( .A(n_374), .B(n_656), .Y(n_713) );
OR2x2_ASAP7_75t_L g881 ( .A(n_374), .B(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x6_ASAP7_75t_L g432 ( .A(n_375), .B(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g478 ( .A(n_375), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_377), .A2(n_652), .B1(n_769), .B2(n_790), .Y(n_768) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx5_ASAP7_75t_L g510 ( .A(n_378), .Y(n_510) );
INVx1_ASAP7_75t_L g1060 ( .A(n_378), .Y(n_1060) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .Y(n_378) );
INVx3_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
INVx1_ASAP7_75t_L g844 ( .A(n_381), .Y(n_844) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x6_ASAP7_75t_L g867 ( .A(n_383), .B(n_868), .Y(n_867) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_385), .B(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g1003 ( .A(n_385), .Y(n_1003) );
NOR3xp33_ASAP7_75t_SL g386 ( .A(n_387), .B(n_418), .C(n_431), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_405), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_400), .B2(n_401), .Y(n_388) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g514 ( .A(n_391), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_391), .A2(n_401), .B1(n_794), .B2(n_795), .Y(n_793) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_391), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_391), .Y(n_1065) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_391), .Y(n_1105) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
BUFx3_ASAP7_75t_L g470 ( .A(n_392), .Y(n_470) );
INVx2_ASAP7_75t_L g607 ( .A(n_392), .Y(n_607) );
INVx1_ASAP7_75t_L g853 ( .A(n_392), .Y(n_853) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g537 ( .A(n_393), .Y(n_537) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_393), .Y(n_836) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_394), .Y(n_717) );
AND2x4_ASAP7_75t_L g403 ( .A(n_395), .B(n_404), .Y(n_403) );
AND2x6_ASAP7_75t_L g401 ( .A(n_396), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g407 ( .A(n_396), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g412 ( .A(n_396), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g518 ( .A(n_396), .B(n_413), .Y(n_518) );
AND2x2_ASAP7_75t_L g585 ( .A(n_396), .B(n_537), .Y(n_585) );
AND2x2_ASAP7_75t_L g587 ( .A(n_396), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g710 ( .A(n_396), .B(n_413), .Y(n_710) );
AND2x2_ASAP7_75t_L g799 ( .A(n_396), .B(n_413), .Y(n_799) );
AND2x2_ASAP7_75t_L g932 ( .A(n_396), .B(n_871), .Y(n_932) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_396), .B(n_413), .Y(n_1070) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
INVx2_ASAP7_75t_L g826 ( .A(n_398), .Y(n_826) );
AND2x2_ASAP7_75t_L g829 ( .A(n_398), .B(n_414), .Y(n_829) );
AND2x4_ASAP7_75t_L g848 ( .A(n_398), .B(n_673), .Y(n_848) );
INVx1_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
INVx1_ASAP7_75t_L g461 ( .A(n_399), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_401), .A2(n_503), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_401), .A2(n_514), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_401), .A2(n_1064), .B1(n_1065), .B2(n_1066), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_401), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_401), .A2(n_1030), .B1(n_1218), .B2(n_1219), .Y(n_1217) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_402), .B(n_424), .Y(n_430) );
BUFx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_403), .Y(n_588) );
BUFx3_ASAP7_75t_L g660 ( .A(n_403), .Y(n_660) );
BUFx2_ASAP7_75t_L g683 ( .A(n_403), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_411), .B2(n_412), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_407), .A2(n_501), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_407), .A2(n_412), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_407), .A2(n_518), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_407), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_407), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g1028 ( .A(n_407), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_407), .A2(n_1068), .B1(n_1069), .B2(n_1070), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_407), .A2(n_518), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_407), .A2(n_799), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
BUFx2_ASAP7_75t_L g658 ( .A(n_408), .Y(n_658) );
BUFx3_ASAP7_75t_L g727 ( .A(n_408), .Y(n_727) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g871 ( .A(n_409), .Y(n_871) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_410), .Y(n_673) );
INVx1_ASAP7_75t_L g935 ( .A(n_412), .Y(n_935) );
INVx1_ASAP7_75t_L g978 ( .A(n_412), .Y(n_978) );
INVx2_ASAP7_75t_SL g723 ( .A(n_413), .Y(n_723) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g663 ( .A(n_414), .Y(n_663) );
BUFx6f_ASAP7_75t_L g834 ( .A(n_414), .Y(n_834) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g428 ( .A(n_415), .Y(n_428) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g521 ( .A(n_420), .Y(n_521) );
NAND2x1_ASAP7_75t_SL g420 ( .A(n_421), .B(n_424), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g841 ( .A(n_421), .B(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_423), .Y(n_678) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_424), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g677 ( .A(n_424), .B(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g679 ( .A(n_424), .B(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g682 ( .A(n_424), .B(n_683), .Y(n_682) );
BUFx4f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx4f_ASAP7_75t_L g979 ( .A(n_426), .Y(n_979) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x6_ASAP7_75t_L g845 ( .A(n_428), .B(n_843), .Y(n_845) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g522 ( .A(n_430), .Y(n_522) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_430), .Y(n_1072) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .A3(n_445), .B1(n_456), .B2(n_463), .B3(n_468), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g523 ( .A1(n_432), .A2(n_456), .A3(n_524), .B1(n_528), .B2(n_539), .B3(n_541), .Y(n_523) );
OAI33xp33_ASAP7_75t_L g594 ( .A1(n_432), .A2(n_595), .A3(n_603), .B1(n_609), .B2(n_613), .B3(n_615), .Y(n_594) );
OAI33xp33_ASAP7_75t_L g801 ( .A1(n_432), .A2(n_456), .A3(n_802), .B1(n_805), .B2(n_808), .B3(n_811), .Y(n_801) );
OAI33xp33_ASAP7_75t_L g1073 ( .A1(n_432), .A2(n_615), .A3(n_1074), .B1(n_1078), .B2(n_1083), .B3(n_1089), .Y(n_1073) );
OAI33xp33_ASAP7_75t_L g1111 ( .A1(n_432), .A2(n_456), .A3(n_1112), .B1(n_1117), .B2(n_1122), .B3(n_1127), .Y(n_1111) );
OAI33xp33_ASAP7_75t_L g1224 ( .A1(n_432), .A2(n_456), .A3(n_1225), .B1(n_1230), .B2(n_1234), .B3(n_1238), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_440), .B1(n_441), .B2(n_444), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_436), .A2(n_536), .B1(n_806), .B2(n_807), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_436), .A2(n_776), .B1(n_789), .B2(n_809), .Y(n_808) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g927 ( .A(n_437), .Y(n_927) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_438), .Y(n_611) );
INVx1_ASAP7_75t_L g1086 ( .A(n_438), .Y(n_1086) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g532 ( .A(n_439), .Y(n_532) );
BUFx2_ASAP7_75t_L g851 ( .A(n_439), .Y(n_851) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g612 ( .A(n_442), .Y(n_612) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g669 ( .A(n_443), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B1(n_450), .B2(n_455), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g464 ( .A(n_447), .Y(n_464) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_450), .A2(n_464), .B1(n_803), .B2(n_804), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_450), .A2(n_858), .B1(n_920), .B2(n_921), .Y(n_919) );
BUFx3_ASAP7_75t_L g1232 ( .A(n_450), .Y(n_1232) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g546 ( .A(n_451), .Y(n_546) );
BUFx3_ASAP7_75t_L g614 ( .A(n_451), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g922 ( .A1(n_451), .A2(n_544), .B1(n_923), .B2(n_924), .Y(n_922) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x2_ASAP7_75t_L g467 ( .A(n_453), .B(n_454), .Y(n_467) );
INVx1_ASAP7_75t_L g681 ( .A(n_454), .Y(n_681) );
CKINVDCx8_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
INVx5_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx6_ASAP7_75t_L g616 ( .A(n_458), .Y(n_616) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx2_ASAP7_75t_L g675 ( .A(n_460), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_464), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g811 ( .A1(n_464), .A2(n_599), .B1(n_786), .B2(n_788), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_465), .A2(n_858), .B1(n_861), .B2(n_1162), .C(n_1163), .Y(n_1161) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g526 ( .A(n_466), .Y(n_526) );
INVx2_ASAP7_75t_L g1166 ( .A(n_466), .Y(n_1166) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g601 ( .A(n_467), .Y(n_601) );
INVx3_ASAP7_75t_L g856 ( .A(n_467), .Y(n_856) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
XNOR2x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_547), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_511), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_479), .B1(n_509), .B2(n_510), .Y(n_474) );
AOI21xp5_ASAP7_75t_SL g999 ( .A1(n_475), .A2(n_1000), .B(n_1027), .Y(n_999) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AOI31xp33_ASAP7_75t_L g731 ( .A1(n_476), .A2(n_732), .A3(n_746), .B(n_763), .Y(n_731) );
AOI31xp33_ASAP7_75t_L g1132 ( .A1(n_476), .A2(n_1133), .A3(n_1140), .B(n_1147), .Y(n_1132) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI31xp33_ASAP7_75t_L g938 ( .A1(n_477), .A2(n_939), .A3(n_945), .B(n_960), .Y(n_938) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g864 ( .A(n_478), .Y(n_864) );
NAND5xp2_ASAP7_75t_L g479 ( .A(n_480), .B(n_491), .C(n_494), .D(n_498), .E(n_507), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_481), .A2(n_492), .B1(n_542), .B2(n_545), .Y(n_541) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_483), .Y(n_1144) );
BUFx3_ASAP7_75t_L g1042 ( .A(n_484), .Y(n_1042) );
INVx2_ASAP7_75t_L g1050 ( .A(n_484), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_484), .Y(n_1196) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g505 ( .A(n_487), .Y(n_505) );
INVx4_ASAP7_75t_L g1040 ( .A(n_487), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g757 ( .A(n_488), .Y(n_757) );
INVx1_ASAP7_75t_L g772 ( .A(n_488), .Y(n_772) );
INVx2_ASAP7_75t_L g941 ( .A(n_488), .Y(n_941) );
INVx1_ASAP7_75t_L g957 ( .A(n_488), .Y(n_957) );
INVx1_ASAP7_75t_L g502 ( .A(n_489), .Y(n_502) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_489), .Y(n_758) );
INVx1_ASAP7_75t_L g1533 ( .A(n_489), .Y(n_1533) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_490), .Y(n_566) );
INVx1_ASAP7_75t_L g575 ( .A(n_490), .Y(n_575) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_490), .Y(n_942) );
INVx2_ASAP7_75t_L g1013 ( .A(n_490), .Y(n_1013) );
INVx1_ASAP7_75t_L g1015 ( .A(n_490), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_493), .A2(n_508), .B1(n_536), .B2(n_540), .Y(n_539) );
INVx2_ASAP7_75t_SL g736 ( .A(n_497), .Y(n_736) );
OAI221xp5_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_501), .B1(n_502), .B2(n_503), .C(n_504), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_510), .A2(n_730), .B(n_731), .Y(n_729) );
AOI21xp33_ASAP7_75t_SL g1130 ( .A1(n_510), .A2(n_1131), .B(n_1132), .Y(n_1130) );
INVx1_ASAP7_75t_L g1214 ( .A(n_510), .Y(n_1214) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_519), .C(n_523), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_533), .B1(n_534), .B2(n_538), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g540 ( .A(n_530), .Y(n_540) );
INVx2_ASAP7_75t_L g1080 ( .A(n_530), .Y(n_1080) );
INVx2_ASAP7_75t_L g1123 ( .A(n_530), .Y(n_1123) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g605 ( .A(n_532), .Y(n_605) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_537), .Y(n_918) );
INVx1_ASAP7_75t_L g992 ( .A(n_537), .Y(n_992) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_544), .A2(n_555), .B1(n_560), .B2(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_544), .Y(n_1090) );
OAI22xp33_ASAP7_75t_L g1230 ( .A1(n_544), .A2(n_1231), .B1(n_1232), .B2(n_1233), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g1238 ( .A1(n_544), .A2(n_1239), .B1(n_1240), .B2(n_1241), .Y(n_1238) );
OAI22xp5_ASAP7_75t_SL g994 ( .A1(n_545), .A2(n_995), .B1(n_996), .B2(n_998), .Y(n_994) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_547), .A2(n_1381), .B1(n_1382), .B2(n_1383), .Y(n_1380) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
XOR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_619), .Y(n_549) );
INVx1_ASAP7_75t_L g617 ( .A(n_551), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_581), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .C(n_567), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_556), .A2(n_570), .B1(n_610), .B2(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B1(n_571), .B2(n_572), .C(n_576), .Y(n_567) );
INVx1_ASAP7_75t_L g640 ( .A(n_568), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_568), .A2(n_771), .B1(n_774), .B2(n_776), .C(n_777), .Y(n_770) );
INVx1_ASAP7_75t_L g739 ( .A(n_569), .Y(n_739) );
INVx1_ASAP7_75t_L g751 ( .A(n_569), .Y(n_751) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g778 ( .A(n_578), .Y(n_778) );
INVx4_ASAP7_75t_L g1006 ( .A(n_578), .Y(n_1006) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_592), .C(n_594), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_589), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_586), .B2(n_587), .Y(n_583) );
INVx2_ASAP7_75t_L g688 ( .A(n_585), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_587), .Y(n_689) );
INVxp67_ASAP7_75t_L g936 ( .A(n_587), .Y(n_936) );
INVx2_ASAP7_75t_SL g719 ( .A(n_588), .Y(n_719) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x6_ASAP7_75t_L g862 ( .A(n_601), .B(n_843), .Y(n_862) );
OAI22xp33_ASAP7_75t_L g985 ( .A1(n_601), .A2(n_858), .B1(n_986), .B2(n_987), .Y(n_985) );
OR2x2_ASAP7_75t_L g1557 ( .A(n_601), .B(n_843), .Y(n_1557) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_607), .B2(n_608), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g983 ( .A(n_605), .Y(n_983) );
INVx2_ASAP7_75t_SL g1554 ( .A(n_605), .Y(n_1554) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g1074 ( .A1(n_614), .A2(n_1075), .B1(n_1076), .B2(n_1077), .Y(n_1074) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_614), .A2(n_1055), .B1(n_1057), .B2(n_1090), .Y(n_1089) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI33xp33_ASAP7_75t_L g711 ( .A1(n_616), .A2(n_712), .A3(n_714), .B1(n_720), .B2(n_724), .B3(n_726), .Y(n_711) );
INVx1_ASAP7_75t_L g930 ( .A(n_616), .Y(n_930) );
INVx1_ASAP7_75t_L g691 ( .A(n_620), .Y(n_691) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .C(n_653), .D(n_684), .Y(n_620) );
OAI31xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_639), .A3(n_649), .B(n_650), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_628), .B2(n_630), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g884 ( .A(n_626), .Y(n_884) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_626), .Y(n_1247) );
INVx2_ASAP7_75t_L g1535 ( .A(n_626), .Y(n_1535) );
INVx1_ASAP7_75t_L g1575 ( .A(n_626), .Y(n_1575) );
INVx1_ASAP7_75t_L g1202 ( .A(n_628), .Y(n_1202) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx3_ASAP7_75t_L g740 ( .A(n_629), .Y(n_740) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_629), .Y(n_775) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_636), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_633), .A2(n_857), .B1(n_860), .B2(n_884), .C(n_885), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_633), .A2(n_743), .B1(n_889), .B2(n_890), .C(n_891), .Y(n_888) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g646 ( .A(n_634), .Y(n_646) );
INVx1_ASAP7_75t_L g955 ( .A(n_634), .Y(n_955) );
BUFx4f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g742 ( .A(n_635), .Y(n_742) );
INVx2_ASAP7_75t_L g908 ( .A(n_635), .Y(n_908) );
INVx1_ASAP7_75t_L g950 ( .A(n_635), .Y(n_950) );
INVx1_ASAP7_75t_L g1528 ( .A(n_635), .Y(n_1528) );
BUFx2_ASAP7_75t_L g1252 ( .A(n_637), .Y(n_1252) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_642), .A2(n_643), .B1(n_677), .B2(n_679), .C(n_682), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_647), .C(n_648), .Y(n_644) );
OAI31xp33_ASAP7_75t_L g1242 ( .A1(n_650), .A2(n_1243), .A3(n_1254), .B(n_1269), .Y(n_1242) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI31xp33_ASAP7_75t_SL g1546 ( .A1(n_651), .A2(n_1547), .A3(n_1548), .B(n_1558), .Y(n_1546) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp67_ASAP7_75t_L g868 ( .A(n_652), .B(n_869), .Y(n_868) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_654), .B(n_676), .Y(n_653) );
AOI33xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .A3(n_661), .B1(n_666), .B2(n_670), .B3(n_674), .Y(n_654) );
BUFx2_ASAP7_75t_SL g861 ( .A(n_656), .Y(n_861) );
INVx1_ASAP7_75t_L g1551 ( .A(n_656), .Y(n_1551) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g824 ( .A(n_660), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g810 ( .A(n_665), .Y(n_810) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g831 ( .A(n_669), .B(n_825), .Y(n_831) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g721 ( .A(n_672), .Y(n_721) );
INVx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx6f_ASAP7_75t_L g838 ( .A(n_673), .Y(n_838) );
INVx2_ASAP7_75t_SL g839 ( .A(n_675), .Y(n_839) );
INVx1_ASAP7_75t_L g1565 ( .A(n_675), .Y(n_1565) );
INVx1_ASAP7_75t_L g702 ( .A(n_677), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_677), .A2(n_679), .B1(n_682), .B2(n_967), .C(n_968), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g1031 ( .A1(n_677), .A2(n_682), .B(n_1007), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_678), .B(n_870), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_678), .B(n_870), .Y(n_1568) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_679), .Y(n_699) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_682), .A2(n_699), .B1(n_700), .B2(n_701), .C(n_703), .Y(n_698) );
XNOR2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_816), .Y(n_692) );
AO22x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_766), .B1(n_814), .B2(n_815), .Y(n_693) );
INVx1_ASAP7_75t_L g815 ( .A(n_694), .Y(n_815) );
XNOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
AND2x4_ASAP7_75t_L g696 ( .A(n_697), .B(n_729), .Y(n_696) );
AND4x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_704), .C(n_707), .D(n_711), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_706), .A2(n_708), .B1(n_742), .B2(n_743), .C(n_745), .Y(n_741) );
BUFx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_716), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_716), .A2(n_996), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
INVx4_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx3_ASAP7_75t_L g725 ( .A(n_717), .Y(n_725) );
INVx2_ASAP7_75t_SL g929 ( .A(n_717), .Y(n_929) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_717), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1173 ( .A(n_717), .Y(n_1173) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g728 ( .A(n_719), .Y(n_728) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1082 ( .A(n_725), .Y(n_1082) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g1576 ( .A(n_739), .B(n_901), .Y(n_1576) );
OAI221xp5_ASAP7_75t_L g1139 ( .A1(n_742), .A2(n_745), .B1(n_884), .B2(n_1106), .C(n_1108), .Y(n_1139) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_749), .B2(n_754), .C(n_759), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_747), .A2(n_759), .B1(n_1126), .B2(n_1141), .C(n_1145), .Y(n_1140) );
INVx1_ASAP7_75t_L g1244 ( .A(n_747), .Y(n_1244) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_753), .B(n_895), .Y(n_1206) );
INVx1_ASAP7_75t_L g1266 ( .A(n_753), .Y(n_1266) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g1253 ( .A(n_759), .Y(n_1253) );
AND2x4_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_761), .B(n_879), .Y(n_1259) );
INVx3_ASAP7_75t_L g814 ( .A(n_766), .Y(n_814) );
INVx1_ASAP7_75t_L g812 ( .A(n_767), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_791), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_779), .C(n_787), .Y(n_769) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g1022 ( .A(n_784), .Y(n_1022) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_785), .Y(n_1146) );
NOR3xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_800), .C(n_801), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_796), .Y(n_792) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_971), .B1(n_972), .B2(n_1092), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g1093 ( .A(n_818), .Y(n_1093) );
XNOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_911), .Y(n_818) );
INVx1_ASAP7_75t_L g909 ( .A(n_820), .Y(n_909) );
NAND4xp25_ASAP7_75t_L g820 ( .A(n_821), .B(n_865), .C(n_872), .D(n_896), .Y(n_820) );
OAI21xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_846), .B(n_863), .Y(n_821) );
INVx8_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_827) );
INVx3_ASAP7_75t_L g1154 ( .A(n_829), .Y(n_1154) );
INVx3_ASAP7_75t_L g1155 ( .A(n_831), .Y(n_1155) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_837), .B(n_840), .Y(n_832) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_835), .Y(n_1120) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx3_ASAP7_75t_L g1088 ( .A(n_836), .Y(n_1088) );
INVx1_ASAP7_75t_L g1564 ( .A(n_838), .Y(n_1564) );
INVx1_ASAP7_75t_L g1170 ( .A(n_839), .Y(n_1170) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g870 ( .A(n_843), .Y(n_870) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
CKINVDCx11_ASAP7_75t_R g1179 ( .A(n_845), .Y(n_1179) );
CKINVDCx6p67_ASAP7_75t_R g847 ( .A(n_848), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_852), .B1(n_853), .B2(n_854), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_850), .A2(n_915), .B1(n_916), .B2(n_917), .Y(n_914) );
BUFx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g991 ( .A(n_851), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_858), .B2(n_860), .C(n_861), .Y(n_855) );
INVx1_ASAP7_75t_L g1115 ( .A(n_856), .Y(n_1115) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_856), .Y(n_1125) );
OAI221xp5_ASAP7_75t_L g1549 ( .A1(n_858), .A2(n_1125), .B1(n_1525), .B2(n_1529), .C(n_1550), .Y(n_1549) );
INVx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
BUFx8_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g1035 ( .A(n_864), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_867), .B(n_1181), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_867), .B(n_1518), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
NOR3xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_880), .C(n_892), .Y(n_872) );
INVx2_ASAP7_75t_L g1190 ( .A(n_874), .Y(n_1190) );
NAND2x1p5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
OR2x6_ASAP7_75t_L g878 ( .A(n_877), .B(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g895 ( .A(n_877), .Y(n_895) );
OR2x2_ASAP7_75t_L g1545 ( .A(n_877), .B(n_879), .Y(n_1545) );
INVx2_ASAP7_75t_L g1191 ( .A(n_878), .Y(n_1191) );
OAI22xp5_ASAP7_75t_SL g880 ( .A1(n_881), .A2(n_883), .B1(n_886), .B2(n_888), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g1520 ( .A1(n_886), .A2(n_1521), .B1(n_1523), .B2(n_1534), .Y(n_1520) );
INVx4_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
BUFx4f_ASAP7_75t_L g1203 ( .A(n_887), .Y(n_1203) );
BUFx2_ASAP7_75t_L g1542 ( .A(n_892), .Y(n_1542) );
AND2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_895), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_902), .B1(n_903), .B2(n_904), .C(n_905), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_897), .A2(n_903), .B1(n_1169), .B2(n_1172), .Y(n_1187) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_900), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g1250 ( .A(n_899), .Y(n_1250) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OR2x6_ASAP7_75t_L g907 ( .A(n_901), .B(n_908), .Y(n_907) );
OR2x2_ASAP7_75t_L g1574 ( .A(n_901), .B(n_1575), .Y(n_1574) );
CKINVDCx6p67_ASAP7_75t_R g1185 ( .A(n_906), .Y(n_1185) );
CKINVDCx6p67_ASAP7_75t_R g1186 ( .A(n_907), .Y(n_1186) );
INVx1_ASAP7_75t_L g1538 ( .A(n_908), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_910), .A2(n_1283), .B1(n_1292), .B2(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_SL g970 ( .A(n_912), .Y(n_970) );
NAND4xp75_ASAP7_75t_L g912 ( .A(n_913), .B(n_933), .C(n_938), .D(n_966), .Y(n_912) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
OAI211xp5_ASAP7_75t_L g954 ( .A1(n_921), .A2(n_955), .B(n_956), .C(n_958), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_923), .A2(n_928), .B1(n_941), .B2(n_942), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_928), .B2(n_929), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g1559 ( .A1(n_929), .A2(n_1080), .B1(n_1560), .B2(n_1561), .C(n_1562), .Y(n_1559) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
NOR2x1_ASAP7_75t_L g933 ( .A(n_934), .B(n_937), .Y(n_933) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_941), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_941), .Y(n_1198) );
INVx2_ASAP7_75t_SL g1248 ( .A(n_942), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_954), .Y(n_945) );
OAI211xp5_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_948), .B(n_951), .C(n_952), .Y(n_946) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx3_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
XNOR2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_1032), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
AND2x2_ASAP7_75t_L g975 ( .A(n_976), .B(n_999), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_980), .Y(n_976) );
OAI221xp5_ASAP7_75t_SL g1014 ( .A1(n_984), .A2(n_987), .B1(n_1011), .B2(n_1015), .C(n_1016), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_990), .B1(n_992), .B2(n_993), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_990), .A2(n_1226), .B1(n_1227), .B2(n_1229), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_990), .A2(n_1235), .B1(n_1236), .B2(n_1237), .Y(n_1234) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g1228 ( .A(n_992), .Y(n_1228) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1076 ( .A(n_997), .Y(n_1076) );
INVx1_ASAP7_75t_L g1168 ( .A(n_997), .Y(n_1168) );
NAND4xp25_ASAP7_75t_SL g1000 ( .A(n_1001), .B(n_1009), .C(n_1014), .D(n_1017), .Y(n_1000) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1013), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1020), .B1(n_1021), .B2(n_1023), .C(n_1024), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1026), .Y(n_1251) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
XNOR2x1_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1091), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1061), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B1(n_1059), .B2(n_1060), .Y(n_1034) );
NAND3xp33_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1047), .C(n_1056), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_1044), .A2(n_1058), .B1(n_1084), .B2(n_1087), .Y(n_1083) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
NOR3xp33_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1071), .C(n_1073), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1067), .Y(n_1062) );
OAI22xp5_ASAP7_75t_SL g1078 ( .A1(n_1079), .A2(n_1080), .B1(n_1081), .B2(n_1082), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_1080), .A2(n_1118), .B1(n_1119), .B2(n_1121), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_1080), .A2(n_1158), .B1(n_1159), .B2(n_1160), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_1084), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1171) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1088), .Y(n_1236) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_1090), .A2(n_1113), .B1(n_1114), .B2(n_1116), .Y(n_1112) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_1096), .A2(n_1097), .B1(n_1209), .B2(n_1272), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1099), .B1(n_1149), .B2(n_1208), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
XNOR2x1_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1148), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1130), .Y(n_1100) );
NOR3xp33_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1110), .C(n_1111), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1107), .Y(n_1102) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1115), .Y(n_1240) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1122) );
INVx2_ASAP7_75t_SL g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1143), .Y(n_1531) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1149), .Y(n_1208) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
NAND3xp33_ASAP7_75t_SL g1151 ( .A(n_1152), .B(n_1180), .C(n_1182), .Y(n_1151) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1167), .B1(n_1168), .B2(n_1169), .C(n_1170), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_1167), .A2(n_1174), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1177), .B1(n_1178), .B2(n_1179), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_1176), .A2(n_1178), .B1(n_1190), .B2(n_1191), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_1179), .A2(n_1567), .B1(n_1569), .B2(n_1570), .Y(n_1566) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1188), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1187), .Y(n_1183) );
NAND3xp33_ASAP7_75t_SL g1188 ( .A(n_1189), .B(n_1192), .C(n_1204), .Y(n_1188) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1190), .Y(n_1544) );
AOI33xp33_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1195), .A3(n_1197), .B1(n_1199), .B2(n_1200), .B3(n_1203), .Y(n_1192) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1194), .Y(n_1522) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1281 ( .A1(n_1207), .A2(n_1282), .B1(n_1289), .B2(n_1290), .Y(n_1281) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1210), .Y(n_1273) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1213), .Y(n_1270) );
NOR3xp33_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1223), .C(n_1224), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1220), .Y(n_1216) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_1218), .A2(n_1222), .B1(n_1248), .B2(n_1262), .C(n_1264), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_1227), .A2(n_1553), .B1(n_1555), .B2(n_1556), .Y(n_1552) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_1228), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1245 ( .A1(n_1229), .A2(n_1231), .B1(n_1246), .B2(n_1248), .C(n_1249), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
OAI221xp5_ASAP7_75t_SL g1274 ( .A1(n_1275), .A2(n_1381), .B1(n_1513), .B2(n_1577), .C(n_1581), .Y(n_1274) );
AND5x1_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1423), .C(n_1461), .D(n_1473), .E(n_1496), .Y(n_1275) );
A2O1A1Ixp33_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1279), .B(n_1366), .C(n_1399), .Y(n_1276) );
OAI211xp5_ASAP7_75t_L g1277 ( .A1(n_1278), .A2(n_1313), .B(n_1353), .C(n_1355), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1304), .Y(n_1278) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1279), .Y(n_1364) );
INVx3_ASAP7_75t_L g1385 ( .A(n_1279), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1279), .B(n_1345), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1279), .B(n_1398), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1279), .B(n_1409), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1279), .B(n_1304), .Y(n_1455) );
INVx3_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1280), .B(n_1304), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1280), .B(n_1388), .Y(n_1387) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1294), .Y(n_1280) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_1282), .A2(n_1292), .B1(n_1335), .B2(n_1336), .Y(n_1334) );
OAI22xp33_ASAP7_75t_L g1347 ( .A1(n_1282), .A2(n_1292), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
BUFx3_ASAP7_75t_L g1381 ( .A(n_1282), .Y(n_1381) );
BUFx6f_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1285), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1284), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1284), .Y(n_1308) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1285), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1288), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1288), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g1383 ( .A(n_1290), .Y(n_1383) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1293), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_1295), .A2(n_1296), .B1(n_1301), .B2(n_1302), .Y(n_1294) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1297), .Y(n_1378) );
AND2x4_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1300), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1298), .B(n_1300), .Y(n_1312) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1299), .B(n_1300), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_1302), .A2(n_1331), .B1(n_1332), .B2(n_1333), .Y(n_1330) );
INVx1_ASAP7_75t_SL g1302 ( .A(n_1303), .Y(n_1302) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1303), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1304), .B(n_1345), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1304), .B(n_1345), .Y(n_1372) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1304), .B(n_1346), .Y(n_1388) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1304), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1304), .B(n_1346), .Y(n_1409) );
OAI211xp5_ASAP7_75t_L g1437 ( .A1(n_1304), .A2(n_1438), .B(n_1440), .C(n_1443), .Y(n_1437) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_1304), .A2(n_1353), .B1(n_1464), .B2(n_1466), .C(n_1467), .Y(n_1463) );
OAI211xp5_ASAP7_75t_L g1475 ( .A1(n_1304), .A2(n_1476), .B(n_1478), .C(n_1484), .Y(n_1475) );
AND2x4_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1311), .Y(n_1304) );
AND2x4_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
OAI21xp33_ASAP7_75t_SL g1591 ( .A1(n_1307), .A2(n_1585), .B(n_1592), .Y(n_1591) );
AND2x4_ASAP7_75t_L g1309 ( .A(n_1308), .B(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1312), .Y(n_1331) );
AOI211xp5_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1322), .B(n_1337), .C(n_1340), .Y(n_1313) );
AOI21xp33_ASAP7_75t_L g1417 ( .A1(n_1314), .A2(n_1418), .B(n_1420), .Y(n_1417) );
AOI21xp5_ASAP7_75t_L g1471 ( .A1(n_1314), .A2(n_1420), .B(n_1457), .Y(n_1471) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1315), .B(n_1338), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1315), .B(n_1328), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1315), .B(n_1322), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1315), .B(n_1323), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1319), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1316), .B(n_1319), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1316), .B(n_1352), .Y(n_1351) );
NOR2xp33_ASAP7_75t_L g1359 ( .A(n_1316), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1316), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1316), .B(n_1329), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1318), .Y(n_1316) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1319), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1319), .B(n_1393), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1319), .B(n_1328), .Y(n_1408) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_1319), .B(n_1328), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1319), .B(n_1322), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1322), .B(n_1392), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1322), .B(n_1430), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1328), .Y(n_1322) );
INVx4_ASAP7_75t_L g1338 ( .A(n_1323), .Y(n_1338) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1323), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1323), .B(n_1354), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1406 ( .A(n_1323), .B(n_1339), .Y(n_1406) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1323), .B(n_1343), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1323), .B(n_1477), .Y(n_1476) );
NOR2xp33_ASAP7_75t_L g1487 ( .A(n_1323), .B(n_1328), .Y(n_1487) );
AND2x6_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1325), .Y(n_1323) );
INVx2_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_1327), .A2(n_1377), .B1(n_1378), .B2(n_1379), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1328), .B(n_1352), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1328), .B(n_1352), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1434 ( .A(n_1328), .B(n_1435), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1328), .B(n_1392), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1328), .B(n_1370), .Y(n_1465) );
CKINVDCx6p67_ASAP7_75t_R g1328 ( .A(n_1329), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1329), .B(n_1339), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1329), .B(n_1370), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1329), .B(n_1393), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1329), .B(n_1392), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1329), .B(n_1430), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1329), .B(n_1351), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1329), .B(n_1393), .Y(n_1495) );
OR2x6_ASAP7_75t_SL g1329 ( .A(n_1330), .B(n_1334), .Y(n_1329) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1338), .B(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1338), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1338), .B(n_1445), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1338), .B(n_1495), .Y(n_1501) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1339), .Y(n_1430) );
NOR2xp33_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1350), .Y(n_1340) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1341), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1342), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1342), .B(n_1408), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1342), .B(n_1415), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1342), .B(n_1439), .Y(n_1438) );
OAI21xp33_ASAP7_75t_L g1456 ( .A1(n_1342), .A2(n_1418), .B(n_1457), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1342), .B(n_1470), .Y(n_1469) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_1342), .B(n_1398), .Y(n_1481) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1344), .Y(n_1363) );
O2A1O1Ixp33_ASAP7_75t_L g1412 ( .A1(n_1344), .A2(n_1413), .B(n_1414), .C(n_1417), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1493 ( .A(n_1344), .B(n_1494), .Y(n_1493) );
INVx2_ASAP7_75t_SL g1344 ( .A(n_1345), .Y(n_1344) );
INVx2_ASAP7_75t_SL g1345 ( .A(n_1346), .Y(n_1345) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_1346), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1350), .B(n_1452), .Y(n_1451) );
NOR3xp33_ASAP7_75t_L g1459 ( .A(n_1350), .B(n_1385), .C(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
OAI222xp33_ASAP7_75t_L g1386 ( .A1(n_1354), .A2(n_1387), .B1(n_1389), .B2(n_1391), .C1(n_1394), .C2(n_1396), .Y(n_1386) );
NOR2xp33_ASAP7_75t_L g1472 ( .A(n_1354), .B(n_1387), .Y(n_1472) );
OAI22xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1359), .B1(n_1362), .B2(n_1365), .Y(n_1355) );
NOR2x1_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1494 ( .A(n_1357), .B(n_1495), .Y(n_1494) );
NOR2x1_ASAP7_75t_R g1507 ( .A(n_1357), .B(n_1508), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_1357), .B(n_1372), .Y(n_1512) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_1361), .A2(n_1405), .B1(n_1407), .B2(n_1409), .C(n_1410), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1361), .B(n_1411), .Y(n_1410) );
A2O1A1Ixp33_ASAP7_75t_L g1467 ( .A1(n_1361), .A2(n_1375), .B(n_1468), .C(n_1471), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1364), .Y(n_1362) );
O2A1O1Ixp33_ASAP7_75t_SL g1423 ( .A1(n_1364), .A2(n_1424), .B(n_1437), .C(n_1446), .Y(n_1423) );
INVxp67_ASAP7_75t_SL g1366 ( .A(n_1367), .Y(n_1366) );
OAI211xp5_ASAP7_75t_L g1399 ( .A1(n_1367), .A2(n_1400), .B(n_1404), .C(n_1412), .Y(n_1399) );
AOI21xp5_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1384), .B(n_1386), .Y(n_1367) );
OAI21xp5_ASAP7_75t_SL g1368 ( .A1(n_1369), .A2(n_1371), .B(n_1373), .Y(n_1368) );
OAI21xp5_ASAP7_75t_SL g1431 ( .A1(n_1371), .A2(n_1432), .B(n_1436), .Y(n_1431) );
OAI21xp33_ASAP7_75t_SL g1447 ( .A1(n_1371), .A2(n_1448), .B(n_1449), .Y(n_1447) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1372), .B(n_1483), .Y(n_1482) );
CKINVDCx14_ASAP7_75t_R g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1375), .B(n_1385), .Y(n_1384) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_1375), .Y(n_1402) );
AOI31xp33_ASAP7_75t_L g1446 ( .A1(n_1375), .A2(n_1447), .A3(n_1450), .B(n_1454), .Y(n_1446) );
OR2x6_ASAP7_75t_SL g1375 ( .A(n_1376), .B(n_1380), .Y(n_1375) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1384), .Y(n_1474) );
INVx1_ASAP7_75t_SL g1403 ( .A(n_1385), .Y(n_1403) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1387), .Y(n_1462) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1388), .Y(n_1445) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1390), .B(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1391), .Y(n_1411) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1392), .Y(n_1508) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1454 ( .A1(n_1395), .A2(n_1414), .B1(n_1455), .B2(n_1456), .C(n_1459), .Y(n_1454) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
AOI21xp5_ASAP7_75t_L g1450 ( .A1(n_1397), .A2(n_1413), .B(n_1451), .Y(n_1450) );
NOR2xp33_ASAP7_75t_L g1466 ( .A(n_1397), .B(n_1428), .Y(n_1466) );
A2O1A1Ixp33_ASAP7_75t_L g1424 ( .A1(n_1398), .A2(n_1425), .B(n_1426), .C(n_1431), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1398), .B(n_1402), .Y(n_1492) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1403), .Y(n_1401) );
OAI21xp33_ASAP7_75t_L g1499 ( .A1(n_1402), .A2(n_1428), .B(n_1500), .Y(n_1499) );
AOI21xp5_ASAP7_75t_L g1506 ( .A1(n_1402), .A2(n_1445), .B(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1407), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1409), .B(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1409), .Y(n_1505) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1414), .Y(n_1504) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_1415), .B(n_1439), .Y(n_1480) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1425), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1426), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1429), .Y(n_1426) );
OAI21xp33_ASAP7_75t_L g1484 ( .A1(n_1427), .A2(n_1485), .B(n_1488), .Y(n_1484) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1428), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1430), .B(n_1487), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1430), .B(n_1511), .Y(n_1510) );
AOI211xp5_ASAP7_75t_L g1461 ( .A1(n_1432), .A2(n_1462), .B(n_1463), .C(n_1472), .Y(n_1461) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1438), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1439), .B(n_1442), .Y(n_1441) );
INVxp67_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1475), .B1(n_1491), .B2(n_1493), .Y(n_1473) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1476), .Y(n_1498) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1477), .Y(n_1483) );
AOI21xp5_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1481), .B(n_1482), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVxp67_ASAP7_75t_SL g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
OAI321xp33_ASAP7_75t_L g1496 ( .A1(n_1492), .A2(n_1497), .A3(n_1498), .B1(n_1499), .B2(n_1502), .C(n_1509), .Y(n_1496) );
INVxp33_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
A2O1A1Ixp33_ASAP7_75t_L g1502 ( .A1(n_1503), .A2(n_1504), .B(n_1505), .C(n_1506), .Y(n_1502) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
XNOR2xp5_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1516), .Y(n_1514) );
HB1xp67_ASAP7_75t_L g1589 ( .A(n_1516), .Y(n_1589) );
AND4x1_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1519), .C(n_1546), .D(n_1571), .Y(n_1516) );
NOR3xp33_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1542), .C(n_1543), .Y(n_1519) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
OAI221xp5_ASAP7_75t_L g1523 ( .A1(n_1524), .A2(n_1525), .B1(n_1526), .B2(n_1529), .C(n_1530), .Y(n_1523) );
INVx2_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
OAI221xp5_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1536), .B1(n_1537), .B2(n_1539), .C(n_1540), .Y(n_1534) );
INVx2_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx2_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
BUFx2_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
HB1xp67_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
INVx4_ASAP7_75t_SL g1577 ( .A(n_1578), .Y(n_1577) );
BUFx3_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
BUFx2_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_1584), .Y(n_1583) );
INVxp33_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
HB1xp67_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
endmodule