module fake_jpeg_13384_n_402 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_402);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_402;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_28),
.A2(n_14),
.B(n_1),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_82),
.B(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_63),
.B(n_66),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_64),
.Y(n_103)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g106 ( 
.A(n_65),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_1),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_81),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_54),
.B1(n_53),
.B2(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_36),
.B(n_1),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_37),
.B1(n_33),
.B2(n_41),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_5),
.B(n_7),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_37),
.B1(n_32),
.B2(n_17),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_92),
.A2(n_94),
.B1(n_114),
.B2(n_130),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_40),
.B1(n_32),
.B2(n_35),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_40),
.B1(n_25),
.B2(n_26),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_70),
.A2(n_35),
.B1(n_38),
.B2(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_42),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_42),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_8),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_19),
.B1(n_38),
.B2(n_22),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_122),
.B1(n_3),
.B2(n_4),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_67),
.A2(n_68),
.B1(n_74),
.B2(n_49),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_59),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_60),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_80),
.B1(n_72),
.B2(n_45),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_147),
.B1(n_174),
.B2(n_176),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_115),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_137),
.B(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_65),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_141),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_64),
.B1(n_69),
.B2(n_75),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_140),
.A2(n_154),
.B1(n_157),
.B2(n_109),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_64),
.C(n_58),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_146),
.C(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_148),
.Y(n_183)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_87),
.C(n_124),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_83),
.B1(n_64),
.B2(n_5),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_3),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_3),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_153),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_104),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_4),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_5),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_164),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_102),
.B(n_7),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_104),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_7),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_9),
.Y(n_194)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_108),
.B(n_8),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_178),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_120),
.A2(n_8),
.B1(n_9),
.B2(n_98),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_97),
.B(n_8),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_111),
.C(n_112),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_95),
.A2(n_9),
.B1(n_99),
.B2(n_101),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_88),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_194),
.B(n_210),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_150),
.A2(n_125),
.B1(n_86),
.B2(n_88),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_134),
.B1(n_158),
.B2(n_160),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_125),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_142),
.B(n_102),
.CI(n_103),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_156),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_131),
.B(n_103),
.C(n_106),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_169),
.B(n_155),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_137),
.B(n_89),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_216),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_89),
.C(n_111),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_138),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_137),
.B(n_86),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_145),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_150),
.B1(n_154),
.B2(n_135),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_177),
.B1(n_149),
.B2(n_151),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_172),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_222),
.B(n_198),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_226),
.A2(n_201),
.B(n_210),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_146),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_249),
.C(n_213),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_199),
.B1(n_206),
.B2(n_208),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_159),
.B1(n_178),
.B2(n_171),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_234),
.B1(n_252),
.B2(n_190),
.Y(n_263)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_236),
.B(n_239),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_241),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_192),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_246),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_248),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_187),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_136),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_181),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_256),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_205),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_251),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_207),
.B1(n_191),
.B2(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_206),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_181),
.B(n_194),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_195),
.B(n_203),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_259),
.A2(n_262),
.B(n_268),
.C(n_270),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_246),
.B(n_241),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_263),
.A2(n_259),
.B1(n_268),
.B2(n_260),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_280),
.B1(n_235),
.B2(n_230),
.Y(n_296)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_219),
.A3(n_185),
.B1(n_197),
.B2(n_218),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_275),
.Y(n_313)
);

NOR2x1_ASAP7_75t_R g268 ( 
.A(n_223),
.B(n_202),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_276),
.C(n_227),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_198),
.B(n_204),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_217),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_198),
.C(n_199),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_255),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_203),
.B1(n_190),
.B2(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_297),
.C(n_300),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_290),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_224),
.B1(n_248),
.B2(n_223),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_291),
.A2(n_306),
.B1(n_310),
.B2(n_266),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_225),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_312),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_203),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_222),
.C(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_231),
.C(n_225),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_307),
.C(n_314),
.Y(n_325)
);

NAND5xp2_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_231),
.C(n_236),
.D(n_256),
.E(n_247),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_243),
.Y(n_307)
);

AO221x1_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_254),
.B1(n_208),
.B2(n_220),
.C(n_209),
.Y(n_308)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_258),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_260),
.A2(n_259),
.B1(n_262),
.B2(n_270),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_282),
.A2(n_244),
.B1(n_228),
.B2(n_235),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_311),
.A2(n_257),
.B1(n_282),
.B2(n_283),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_271),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_229),
.Y(n_314)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_320),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_322),
.A2(n_333),
.B1(n_294),
.B2(n_302),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_272),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_329),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_301),
.Y(n_326)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_293),
.Y(n_328)
);

INVx13_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_330),
.A2(n_305),
.B(n_313),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_332),
.A2(n_296),
.B(n_305),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_291),
.A2(n_261),
.B1(n_287),
.B2(n_274),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_273),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_304),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_273),
.C(n_284),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_324),
.C(n_289),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_333),
.C(n_334),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g365 ( 
.A1(n_339),
.A2(n_332),
.B(n_316),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_340),
.A2(n_330),
.B(n_326),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_315),
.Y(n_355)
);

BUFx12_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_349),
.Y(n_361)
);

BUFx12f_ASAP7_75t_SL g346 ( 
.A(n_329),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_315),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_300),
.C(n_305),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_348),
.C(n_351),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_305),
.C(n_301),
.Y(n_348)
);

AOI321xp33_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_306),
.A3(n_279),
.B1(n_278),
.B2(n_298),
.C(n_294),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_303),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_298),
.C(n_293),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_353),
.C(n_327),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_286),
.C(n_274),
.Y(n_353)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_364),
.C(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_331),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_360),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_340),
.B(n_332),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_278),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_363),
.Y(n_373)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_365),
.A2(n_341),
.B1(n_345),
.B2(n_346),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_316),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_339),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_368),
.B(n_369),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_338),
.C(n_347),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_376),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_318),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_374),
.B(n_257),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_348),
.C(n_337),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_SL g384 ( 
.A(n_375),
.B(n_350),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_378),
.A2(n_359),
.B1(n_365),
.B2(n_336),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_383),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_377),
.A2(n_355),
.B1(n_350),
.B2(n_354),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_381),
.A2(n_368),
.B1(n_369),
.B2(n_344),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_336),
.B1(n_366),
.B2(n_328),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_386),
.B(n_342),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_372),
.A2(n_321),
.B1(n_342),
.B2(n_272),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_387),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_281),
.Y(n_387)
);

NOR2x1p5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_393),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_392),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_344),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_388),
.B(n_382),
.CI(n_379),
.CON(n_395),
.SN(n_395)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_395),
.A2(n_396),
.B(n_221),
.Y(n_399)
);

AOI322xp5_ASAP7_75t_L g396 ( 
.A1(n_389),
.A2(n_382),
.A3(n_281),
.B1(n_209),
.B2(n_220),
.C1(n_242),
.C2(n_221),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_397),
.A2(n_221),
.B(n_211),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_399),
.C(n_395),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_394),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_401),
.B(n_394),
.Y(n_402)
);


endmodule