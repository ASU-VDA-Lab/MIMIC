module fake_ariane_1764_n_1857 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1857);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1857;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_14),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_38),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_74),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_73),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_109),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_18),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_41),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_100),
.Y(n_199)
);

BUFx8_ASAP7_75t_SL g200 ( 
.A(n_75),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_3),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_45),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_96),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_58),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_26),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_136),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_69),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_144),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_139),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_18),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_157),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_133),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_128),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_37),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

INVx4_ASAP7_75t_R g225 ( 
.A(n_146),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_95),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_69),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_31),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_107),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_81),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_91),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_103),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_98),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_68),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_46),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_105),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_101),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_51),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_138),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_132),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_64),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_79),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_24),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_102),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_65),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_141),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_42),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_110),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_13),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_83),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_145),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_44),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_14),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_127),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_2),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_38),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_28),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_6),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_129),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_43),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_60),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_183),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_7),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_137),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_168),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_71),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_3),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_2),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_55),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_1),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_153),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_150),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_67),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_89),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_43),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_25),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_78),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_169),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_62),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_5),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_90),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_122),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_56),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_99),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_34),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_11),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_29),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_39),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_123),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_176),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_33),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_165),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_23),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_155),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_70),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_97),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_130),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_143),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_167),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_20),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_63),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_154),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_156),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_10),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_118),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_62),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_106),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_42),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_25),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_4),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_104),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_50),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_117),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_44),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_9),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_60),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_39),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_17),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_61),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_86),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_0),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_119),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_131),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_108),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_87),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_50),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_52),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_152),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_30),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_175),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_49),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_29),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_57),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_59),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_48),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_173),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_57),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_177),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_67),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_49),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_82),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_48),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_134),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_68),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_200),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_268),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_194),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_244),
.B(n_4),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_187),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_237),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g381 ( 
.A(n_184),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_294),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_187),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_187),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_341),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_250),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_5),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_187),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_270),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_295),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_213),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_187),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_198),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_198),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_340),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_214),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_214),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_214),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_205),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_244),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_296),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_214),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_254),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_254),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_354),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_254),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_254),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_262),
.B(n_6),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_205),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_230),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_231),
.Y(n_413)
);

INVxp33_ASAP7_75t_SL g414 ( 
.A(n_184),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_254),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_246),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_211),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_233),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_246),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_240),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_243),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_302),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_192),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_7),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_255),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_302),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_276),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_310),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_206),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_186),
.B(n_8),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_257),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_289),
.B(n_9),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_310),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_261),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_269),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_271),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_353),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_282),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_272),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_358),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_190),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_213),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_289),
.B(n_291),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_210),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_273),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_324),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_324),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_216),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_274),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_222),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_242),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_259),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_275),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_189),
.B(n_11),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_264),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_280),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_267),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_281),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_290),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_293),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_291),
.B(n_12),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_330),
.B(n_12),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_297),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_299),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_304),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_276),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_306),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_330),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_195),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_393),
.B(n_346),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_384),
.A2(n_392),
.B(n_388),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_378),
.B(n_363),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_209),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_410),
.B(n_199),
.Y(n_483)
);

BUFx8_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_394),
.B(n_346),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_388),
.A2(n_218),
.B(n_215),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_379),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_430),
.A2(n_232),
.B(n_224),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_391),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_403),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_391),
.B(n_348),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_376),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_394),
.B(n_348),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_406),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_422),
.B(n_199),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_363),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_455),
.A2(n_428),
.B(n_426),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_408),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_424),
.B(n_185),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_426),
.B(n_329),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_428),
.B(n_287),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

AND3x1_ASAP7_75t_L g518 ( 
.A(n_387),
.B(n_343),
.C(n_333),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_415),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_417),
.B(n_241),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_433),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_400),
.B(n_344),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_433),
.A2(n_236),
.B(n_234),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

XNOR2x2_ASAP7_75t_L g526 ( 
.A(n_444),
.B(n_251),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_411),
.B(n_239),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_427),
.B(n_345),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_438),
.B(n_245),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

CKINVDCx6p67_ASAP7_75t_R g533 ( 
.A(n_417),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_416),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_385),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_445),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_467),
.B(n_449),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_449),
.B(n_360),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_381),
.B(n_248),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_451),
.B(n_249),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_451),
.B(n_361),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_386),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_463),
.C(n_462),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_476),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_545),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_SL g555 ( 
.A1(n_483),
.A2(n_432),
.B(n_378),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_526),
.A2(n_432),
.B1(n_414),
.B2(n_423),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_540),
.B(n_439),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_395),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_515),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_478),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_494),
.B(n_412),
.Y(n_561)
);

BUFx8_ASAP7_75t_SL g562 ( 
.A(n_482),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_477),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_418),
.C(n_413),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_494),
.B(n_420),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_484),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_494),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_539),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_529),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_541),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_496),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_529),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_512),
.B(n_421),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_542),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_526),
.A2(n_443),
.B1(n_447),
.B2(n_364),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_540),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_518),
.A2(n_436),
.B1(n_457),
.B2(n_454),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_529),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_470),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_477),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_496),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_512),
.B(n_425),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_496),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_431),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_482),
.B(n_452),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_484),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_478),
.B(n_434),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_486),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_478),
.B(n_437),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_540),
.B(n_446),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_540),
.B(n_450),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

AND3x2_ASAP7_75t_L g597 ( 
.A(n_520),
.B(n_469),
.C(n_401),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_541),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_541),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_538),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_538),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_508),
.B(n_287),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_544),
.B(n_452),
.Y(n_604)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_491),
.A2(n_288),
.B(n_279),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_540),
.A2(n_201),
.B1(n_197),
.B2(n_192),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_544),
.B(n_453),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_522),
.B(n_453),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_506),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_520),
.A2(n_533),
.B1(n_540),
.B2(n_316),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_540),
.B(n_389),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_500),
.B(n_456),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_522),
.B(n_456),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_540),
.B(n_301),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_540),
.B(n_390),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_522),
.B(n_458),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_477),
.A2(n_370),
.B1(n_347),
.B2(n_337),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_SL g620 ( 
.A1(n_491),
.A2(n_468),
.B(n_459),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_508),
.B(n_287),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_525),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_543),
.B(n_458),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_500),
.B(n_459),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_529),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_525),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_531),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_506),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_531),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_543),
.B(n_460),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_527),
.B(n_508),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_527),
.B(n_508),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_482),
.B(n_468),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_534),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_504),
.B(n_402),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_510),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_508),
.B(n_287),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_501),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_484),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_515),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_506),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_529),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_544),
.B(n_460),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_508),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_SL g648 ( 
.A1(n_526),
.A2(n_405),
.B1(n_313),
.B2(n_338),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_504),
.B(n_461),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_514),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_509),
.A2(n_241),
.B1(n_278),
.B2(n_464),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_514),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_500),
.B(n_461),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_482),
.B(n_464),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_470),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_470),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_500),
.B(n_466),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_510),
.B(n_319),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_484),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_510),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_514),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_548),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_529),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_536),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_529),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_536),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_500),
.B(n_465),
.Y(n_667)
);

AND3x1_ASAP7_75t_L g668 ( 
.A(n_501),
.B(n_466),
.C(n_465),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_504),
.B(n_474),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_514),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_498),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_471),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_509),
.B(n_287),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_471),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_509),
.A2(n_513),
.B1(n_547),
.B2(n_544),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_473),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_515),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_486),
.Y(n_679)
);

INVxp33_ASAP7_75t_SL g680 ( 
.A(n_548),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_473),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_471),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_486),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_488),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_544),
.B(n_327),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_544),
.B(n_349),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_475),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_488),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_500),
.B(n_208),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_523),
.A2(n_320),
.B1(n_318),
.B2(n_283),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_547),
.B(n_351),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_488),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_546),
.A2(n_227),
.B1(n_203),
.B2(n_202),
.Y(n_693)
);

INVx4_ASAP7_75t_SL g694 ( 
.A(n_515),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_515),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_583),
.Y(n_696)
);

BUFx8_ASAP7_75t_L g697 ( 
.A(n_674),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_550),
.A2(n_484),
.B1(n_486),
.B2(n_513),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_582),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_649),
.B(n_523),
.Y(n_700)
);

NAND3xp33_ASAP7_75t_SL g701 ( 
.A(n_580),
.B(n_380),
.C(n_377),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_582),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_575),
.A2(n_350),
.B1(n_227),
.B2(n_322),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_674),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_566),
.B(n_185),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_669),
.B(n_523),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_585),
.B(n_528),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_554),
.B(n_484),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_631),
.B(n_632),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_623),
.B(n_528),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_572),
.B(n_528),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_639),
.B(n_188),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_630),
.B(n_474),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_572),
.B(n_547),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_662),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_672),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_604),
.B(n_474),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_638),
.B(n_533),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_604),
.B(n_485),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_672),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_607),
.B(n_485),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_563),
.B(n_533),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_675),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_607),
.B(n_485),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_645),
.B(n_613),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_645),
.B(n_547),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_639),
.B(n_188),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_657),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_613),
.B(n_624),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_613),
.B(n_547),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_549),
.B(n_513),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_655),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_560),
.A2(n_595),
.B(n_572),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_635),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_682),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_595),
.A2(n_546),
.B(n_475),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_624),
.B(n_547),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_597),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_646),
.B(n_524),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_624),
.B(n_509),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_561),
.B(n_509),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_659),
.B(n_646),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_590),
.B(n_524),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_655),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_668),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_587),
.B(n_509),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_682),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_684),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_592),
.B(n_513),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_549),
.Y(n_750)
);

INVxp33_ASAP7_75t_L g751 ( 
.A(n_638),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_591),
.B(n_513),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_676),
.B(n_472),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_656),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_591),
.B(n_191),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_554),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_656),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_677),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_569),
.B(n_480),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_571),
.B(n_480),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_636),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_576),
.B(n_530),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_659),
.B(n_191),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_554),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_662),
.B(n_407),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_688),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_662),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_681),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_687),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_680),
.B(n_429),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_606),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_608),
.B(n_614),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_617),
.B(n_530),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_588),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_622),
.B(n_532),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_578),
.B(n_440),
.Y(n_777)
);

AND2x6_ASAP7_75t_SL g778 ( 
.A(n_588),
.B(n_633),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_688),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_692),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_594),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_555),
.B(n_284),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_591),
.B(n_193),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_692),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_564),
.B(n_532),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_562),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_611),
.B(n_292),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_588),
.B(n_441),
.Y(n_788)
);

BUFx5_ASAP7_75t_L g789 ( 
.A(n_636),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_549),
.B(n_193),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_598),
.B(n_196),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_562),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_599),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_619),
.B(n_322),
.C(n_203),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_556),
.B(n_486),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_657),
.A2(n_339),
.B1(n_365),
.B2(n_356),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_551),
.B(n_552),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_633),
.B(n_241),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_693),
.A2(n_339),
.B1(n_365),
.B2(n_362),
.C(n_356),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_679),
.A2(n_486),
.B1(n_532),
.B2(n_535),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_626),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_627),
.B(n_532),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_SL g803 ( 
.A(n_680),
.B(n_567),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_629),
.B(n_535),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_R g805 ( 
.A(n_567),
.B(n_335),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_689),
.B(n_300),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_634),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_647),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_657),
.B(n_690),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_664),
.B(n_535),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_551),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_666),
.B(n_535),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_612),
.B(n_479),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_657),
.A2(n_633),
.B1(n_654),
.B2(n_653),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_616),
.B(n_479),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_557),
.A2(n_219),
.B1(n_221),
.B2(n_373),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_593),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_551),
.B(n_196),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_685),
.B(n_686),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_551),
.B(n_204),
.Y(n_820)
);

INVx8_ASAP7_75t_L g821 ( 
.A(n_633),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_685),
.B(n_497),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_686),
.B(n_497),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_551),
.B(n_204),
.Y(n_824)
);

INVx8_ASAP7_75t_L g825 ( 
.A(n_654),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_557),
.B(n_303),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_573),
.B(n_577),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_573),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_552),
.B(n_207),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_691),
.B(n_305),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_691),
.B(n_505),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_577),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_584),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_620),
.A2(n_492),
.B(n_489),
.C(n_517),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_584),
.Y(n_835)
);

OAI221xp5_ASAP7_75t_L g836 ( 
.A1(n_651),
.A2(n_347),
.B1(n_369),
.B2(n_370),
.C(n_372),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_654),
.B(n_350),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_558),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_552),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_679),
.B(n_309),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_586),
.B(n_505),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_552),
.B(n_207),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_602),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_586),
.B(n_511),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_552),
.B(n_212),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_603),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_602),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_602),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_660),
.A2(n_601),
.B(n_609),
.C(n_600),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_610),
.B(n_516),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_610),
.B(n_516),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_589),
.B(n_355),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_660),
.B(n_679),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_817),
.A2(n_658),
.B(n_568),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_696),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_775),
.B(n_728),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_707),
.B(n_618),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_704),
.B(n_589),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_699),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_848),
.Y(n_860)
);

AOI21xp33_ASAP7_75t_L g861 ( 
.A1(n_787),
.A2(n_648),
.B(n_683),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_700),
.B(n_628),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_734),
.B(n_683),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_709),
.A2(n_568),
.B(n_565),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_809),
.A2(n_640),
.B(n_642),
.C(n_670),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_786),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_733),
.A2(n_568),
.B(n_579),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_702),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_750),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_697),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_703),
.A2(n_640),
.B(n_642),
.C(n_644),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_710),
.B(n_644),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_751),
.B(n_278),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_706),
.B(n_713),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_795),
.A2(n_683),
.B1(n_621),
.B2(n_637),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_771),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_772),
.B(n_745),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_729),
.A2(n_652),
.B1(n_650),
.B2(n_661),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_839),
.B(n_650),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_750),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_732),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_697),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_774),
.B(n_652),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_725),
.B(n_670),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_809),
.A2(n_673),
.B1(n_602),
.B2(n_637),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_355),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_806),
.B(n_553),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_806),
.B(n_711),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_853),
.A2(n_615),
.B(n_574),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_805),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_723),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_711),
.B(n_553),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_739),
.A2(n_615),
.B(n_492),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_763),
.B(n_602),
.Y(n_894)
);

O2A1O1Ixp5_ASAP7_75t_L g895 ( 
.A1(n_790),
.A2(n_663),
.B(n_665),
.C(n_574),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_739),
.A2(n_783),
.B(n_755),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_797),
.A2(n_581),
.B(n_570),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_730),
.A2(n_570),
.B1(n_581),
.B2(n_665),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_787),
.B(n_369),
.C(n_362),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_717),
.B(n_602),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_719),
.B(n_621),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_839),
.B(n_596),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_755),
.A2(n_368),
.B(n_359),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_838),
.B(n_756),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_736),
.A2(n_643),
.B(n_625),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_786),
.B(n_625),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_708),
.A2(n_673),
.B1(n_637),
.B2(n_621),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_839),
.B(n_643),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_750),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_813),
.A2(n_663),
.B(n_643),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_721),
.B(n_621),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_744),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_805),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_724),
.B(n_621),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_815),
.A2(n_671),
.B(n_605),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_754),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_849),
.A2(n_671),
.B(n_637),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_765),
.B(n_671),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_757),
.Y(n_919)
);

AOI21xp33_ASAP7_75t_L g920 ( 
.A1(n_826),
.A2(n_605),
.B(n_372),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_827),
.A2(n_605),
.B(n_489),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_773),
.B(n_621),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_801),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_783),
.A2(n_492),
.B(n_489),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_741),
.A2(n_366),
.B(n_321),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_753),
.B(n_637),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_751),
.B(n_722),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_752),
.A2(n_321),
.B(n_228),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_768),
.B(n_517),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_752),
.A2(n_228),
.B(n_217),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_737),
.A2(n_314),
.B1(n_311),
.B2(n_312),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_807),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_834),
.A2(n_673),
.B(n_519),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_714),
.A2(n_749),
.B(n_760),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_852),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_SL g936 ( 
.A1(n_834),
.A2(n_521),
.B(n_519),
.C(n_493),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_708),
.A2(n_521),
.B(n_490),
.C(n_493),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_714),
.A2(n_223),
.B(n_217),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_728),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_740),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_761),
.A2(n_223),
.B(n_220),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_808),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_726),
.B(n_673),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_766),
.B(n_278),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_814),
.A2(n_673),
.B1(n_226),
.B2(n_326),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_746),
.B(n_673),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_759),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_716),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_738),
.B(n_374),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_790),
.A2(n_212),
.B(n_226),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_775),
.B(n_694),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_830),
.B(n_325),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_715),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_830),
.B(n_328),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_750),
.B(n_328),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_837),
.B(n_323),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_811),
.B(n_331),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_811),
.B(n_331),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_836),
.A2(n_493),
.B(n_503),
.C(n_502),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_698),
.A2(n_336),
.B1(n_342),
.B2(n_352),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_792),
.B(n_336),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_848),
.Y(n_962)
);

INVx11_ASAP7_75t_L g963 ( 
.A(n_731),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_818),
.A2(n_352),
.B(n_342),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_818),
.A2(n_357),
.B(n_366),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_769),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_770),
.B(n_826),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_800),
.A2(n_503),
.B(n_490),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_819),
.B(n_357),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_800),
.A2(n_840),
.B(n_832),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_821),
.Y(n_971)
);

OR2x2_ASAP7_75t_SL g972 ( 
.A(n_701),
.B(n_803),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_820),
.A2(n_373),
.B(n_235),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_782),
.B(n_488),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_782),
.B(n_490),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_840),
.B(n_490),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_820),
.A2(n_308),
.B(n_238),
.Y(n_977)
);

AND2x2_ASAP7_75t_SL g978 ( 
.A(n_795),
.B(n_225),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_824),
.A2(n_315),
.B(n_247),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_852),
.B(n_495),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_811),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_828),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_731),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_824),
.A2(n_317),
.B(n_252),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_698),
.A2(n_495),
.B1(n_502),
.B2(n_503),
.Y(n_985)
);

OAI321xp33_ASAP7_75t_L g986 ( 
.A1(n_814),
.A2(n_495),
.A3(n_503),
.B1(n_502),
.B2(n_487),
.C(n_481),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_798),
.B(n_720),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_835),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_796),
.A2(n_502),
.B(n_481),
.C(n_487),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_735),
.B(n_481),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_788),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_829),
.A2(n_298),
.B(n_253),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_821),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_715),
.B(n_16),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_778),
.B(n_16),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_747),
.Y(n_996)
);

CKINVDCx10_ASAP7_75t_R g997 ( 
.A(n_799),
.Y(n_997)
);

AO22x1_ASAP7_75t_L g998 ( 
.A1(n_777),
.A2(n_695),
.B1(n_559),
.B2(n_678),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_781),
.B(n_481),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_731),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_793),
.B(n_487),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_821),
.B(n_17),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_825),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_794),
.A2(n_487),
.B(n_498),
.C(n_499),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_825),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_742),
.A2(n_498),
.B1(n_499),
.B2(n_507),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_825),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_748),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_731),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_833),
.A2(n_515),
.B(n_695),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_731),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_847),
.B(n_694),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_776),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_762),
.B(n_498),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_742),
.Y(n_1015)
);

NOR2x1p5_ASAP7_75t_L g1016 ( 
.A(n_822),
.B(n_256),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_843),
.B(n_694),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_816),
.B(n_258),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_842),
.A2(n_307),
.B(n_260),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_762),
.B(n_498),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_846),
.B(n_263),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_845),
.B(n_19),
.Y(n_1022)
);

NOR2xp67_ASAP7_75t_L g1023 ( 
.A(n_876),
.B(n_785),
.Y(n_1023)
);

OAI22x1_ASAP7_75t_L g1024 ( 
.A1(n_995),
.A2(n_956),
.B1(n_945),
.B2(n_935),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_877),
.B(n_791),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_864),
.A2(n_705),
.B(n_727),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_854),
.A2(n_712),
.B(n_764),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_874),
.B(n_802),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_1022),
.A2(n_812),
.B(n_804),
.C(n_810),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_855),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_993),
.B(n_758),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_858),
.B(n_767),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_952),
.A2(n_851),
.B(n_850),
.C(n_844),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_R g1034 ( 
.A(n_913),
.B(n_823),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_991),
.B(n_877),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_887),
.A2(n_841),
.B(n_789),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_1000),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_940),
.B(n_831),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_956),
.B(n_779),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_923),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_1022),
.A2(n_784),
.B(n_780),
.C(n_499),
.Y(n_1041)
);

OAI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_954),
.A2(n_265),
.B(n_266),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_960),
.A2(n_277),
.B(n_285),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_932),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_934),
.A2(n_789),
.B(n_762),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_967),
.A2(n_789),
.B1(n_762),
.B2(n_286),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_921),
.A2(n_789),
.B(n_762),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_888),
.A2(n_863),
.B1(n_983),
.B2(n_963),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_1000),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_994),
.A2(n_789),
.B(n_20),
.C(n_22),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_1000),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_865),
.A2(n_515),
.B(n_789),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_1000),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_859),
.A2(n_498),
.B1(n_499),
.B2(n_507),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_863),
.A2(n_507),
.B1(n_499),
.B2(n_641),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_983),
.A2(n_507),
.B1(n_499),
.B2(n_641),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_927),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_994),
.A2(n_931),
.B(n_1004),
.C(n_857),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_873),
.B(n_944),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_890),
.A2(n_953),
.B1(n_949),
.B2(n_1002),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_883),
.A2(n_695),
.B(n_678),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_983),
.B(n_695),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_983),
.A2(n_507),
.B1(n_499),
.B2(n_641),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1009),
.B(n_695),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_939),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_866),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_949),
.A2(n_515),
.B1(n_641),
.B2(n_559),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_1009),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_1009),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_1004),
.A2(n_19),
.B(n_22),
.C(n_28),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_861),
.A2(n_515),
.B1(n_641),
.B2(n_559),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_920),
.A2(n_507),
.B(n_499),
.C(n_678),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_942),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1014),
.A2(n_678),
.B(n_559),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1009),
.B(n_507),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_980),
.B(n_32),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_904),
.B(n_229),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_SL g1078 ( 
.A(n_993),
.B(n_515),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_939),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_951),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_904),
.B(n_1013),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_966),
.B(n_32),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_868),
.B(n_33),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_865),
.A2(n_515),
.B(n_334),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_881),
.B(n_34),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_856),
.B(n_334),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_912),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_916),
.B(n_36),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_886),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_899),
.B(n_47),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_866),
.Y(n_1092)
);

INVx8_ASAP7_75t_L g1093 ( 
.A(n_951),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_987),
.B(n_51),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_970),
.A2(n_334),
.B(n_229),
.C(n_54),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_995),
.B(n_52),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1011),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1011),
.A2(n_919),
.B1(n_884),
.B2(n_872),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_1012),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_922),
.A2(n_334),
.B(n_229),
.C(n_63),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_856),
.B(n_53),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_862),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_1102)
);

OAI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1002),
.A2(n_66),
.B1(n_334),
.B2(n_229),
.C(n_77),
.Y(n_1103)
);

OAI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_961),
.A2(n_882),
.B1(n_1018),
.B2(n_969),
.C(n_997),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_982),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_937),
.A2(n_334),
.B(n_229),
.C(n_84),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1005),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1015),
.B(n_929),
.Y(n_1108)
);

OA22x2_ASAP7_75t_L g1109 ( 
.A1(n_870),
.A2(n_885),
.B1(n_988),
.B2(n_971),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_972),
.B(n_72),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1016),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_948),
.Y(n_1112)
);

NAND2x1_ASAP7_75t_L g1113 ( 
.A(n_869),
.B(n_76),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1003),
.B(n_334),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_L g1115 ( 
.A1(n_924),
.A2(n_229),
.B(n_92),
.C(n_93),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_971),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1007),
.B(n_88),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_894),
.A2(n_229),
.B(n_115),
.C(n_116),
.Y(n_1118)
);

AND2x6_ASAP7_75t_L g1119 ( 
.A(n_869),
.B(n_112),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_943),
.A2(n_120),
.B1(n_124),
.B2(n_140),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1015),
.B(n_149),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_996),
.B(n_181),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_937),
.A2(n_163),
.B(n_164),
.C(n_166),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_869),
.Y(n_1124)
);

XNOR2xp5_ASAP7_75t_L g1125 ( 
.A(n_906),
.B(n_170),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_978),
.B(n_892),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1008),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_891),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_941),
.B(n_938),
.C(n_925),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_880),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_981),
.A2(n_918),
.B1(n_901),
.B2(n_914),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_900),
.A2(n_911),
.B1(n_875),
.B2(n_933),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_955),
.A2(n_958),
.B(n_957),
.C(n_936),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1020),
.A2(n_915),
.B(n_867),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_875),
.A2(n_946),
.B1(n_974),
.B2(n_975),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_981),
.A2(n_918),
.B1(n_909),
.B2(n_957),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_909),
.Y(n_1137)
);

INVx3_ASAP7_75t_SL g1138 ( 
.A(n_955),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_958),
.A2(n_936),
.B(n_871),
.C(n_878),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_L g1140 ( 
.A(n_950),
.B(n_964),
.C(n_965),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1020),
.A2(n_910),
.B(n_897),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_909),
.B(n_928),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_930),
.B(n_926),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_898),
.A2(n_905),
.B(n_895),
.C(n_973),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_999),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1017),
.Y(n_1146)
);

BUFx4f_ASAP7_75t_L g1147 ( 
.A(n_1017),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_986),
.B(n_907),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1012),
.B(n_860),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_998),
.B(n_902),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1021),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_860),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_908),
.B(n_879),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_903),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_959),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_917),
.A2(n_989),
.B(n_889),
.C(n_968),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_962),
.Y(n_1157)
);

OAI21xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1001),
.A2(n_1010),
.B(n_1019),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_962),
.Y(n_1159)
);

AOI221xp5_ASAP7_75t_L g1160 ( 
.A1(n_977),
.A2(n_992),
.B1(n_979),
.B2(n_984),
.C(n_985),
.Y(n_1160)
);

NOR3xp33_ASAP7_75t_SL g1161 ( 
.A(n_1006),
.B(n_990),
.C(n_896),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_893),
.B(n_639),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_864),
.A2(n_817),
.B(n_854),
.Y(n_1163)
);

NOR4xp25_ASAP7_75t_L g1164 ( 
.A(n_1088),
.B(n_1090),
.C(n_1103),
.D(n_1050),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1156),
.A2(n_1135),
.B(n_1095),
.Y(n_1165)
);

AOI221x1_ASAP7_75t_L g1166 ( 
.A1(n_1024),
.A2(n_1102),
.B1(n_1097),
.B2(n_1100),
.C(n_1088),
.Y(n_1166)
);

AO32x2_ASAP7_75t_L g1167 ( 
.A1(n_1098),
.A2(n_1135),
.A3(n_1132),
.B1(n_1131),
.B2(n_1136),
.Y(n_1167)
);

BUFx2_ASAP7_75t_R g1168 ( 
.A(n_1066),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1093),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1025),
.B(n_1053),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1035),
.A2(n_1091),
.B1(n_1059),
.B2(n_1096),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1028),
.A2(n_1082),
.B1(n_1058),
.B2(n_1101),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1132),
.A2(n_1072),
.A3(n_1041),
.B(n_1154),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_1093),
.B(n_1101),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1109),
.A2(n_1127),
.B1(n_1057),
.B2(n_1039),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1104),
.A2(n_1094),
.B1(n_1043),
.B2(n_1070),
.C(n_1079),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_1046),
.C(n_1077),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1052),
.A2(n_1144),
.B(n_1139),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1080),
.B(n_1057),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1040),
.Y(n_1180)
);

NAND2x2_ASAP7_75t_L g1181 ( 
.A(n_1111),
.B(n_1092),
.Y(n_1181)
);

CKINVDCx16_ASAP7_75t_R g1182 ( 
.A(n_1034),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1080),
.B(n_1065),
.Y(n_1183)
);

AOI221x1_ASAP7_75t_L g1184 ( 
.A1(n_1140),
.A2(n_1110),
.B1(n_1118),
.B2(n_1085),
.C(n_1048),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1030),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1038),
.B(n_1032),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1085),
.A2(n_1143),
.B(n_1142),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1060),
.B(n_1116),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1161),
.A2(n_1115),
.B(n_1126),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1133),
.A2(n_1106),
.B(n_1042),
.C(n_1033),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_1117),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1138),
.B(n_1151),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1029),
.A2(n_1148),
.B(n_1158),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1044),
.B(n_1073),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1105),
.B(n_1081),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1123),
.A2(n_1023),
.B(n_1083),
.C(n_1160),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1155),
.A2(n_1086),
.B1(n_1089),
.B2(n_1084),
.Y(n_1197)
);

BUFx10_ASAP7_75t_L g1198 ( 
.A(n_1124),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_1053),
.Y(n_1199)
);

CKINVDCx11_ASAP7_75t_R g1200 ( 
.A(n_1107),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1055),
.A2(n_1145),
.B(n_1150),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1112),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1150),
.A2(n_1162),
.B(n_1054),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1076),
.A2(n_1147),
.B1(n_1159),
.B2(n_1107),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1128),
.Y(n_1205)
);

INVx8_ASAP7_75t_L g1206 ( 
.A(n_1093),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1162),
.A2(n_1054),
.B(n_1075),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_SL g1208 ( 
.A(n_1053),
.B(n_1153),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1129),
.A2(n_1067),
.B(n_1061),
.Y(n_1209)
);

AO21x1_ASAP7_75t_L g1210 ( 
.A1(n_1121),
.A2(n_1120),
.B(n_1114),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1074),
.A2(n_1071),
.B(n_1153),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1125),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1122),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_L g1214 ( 
.A(n_1037),
.B(n_1049),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1153),
.A2(n_1157),
.B1(n_1146),
.B2(n_1152),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1108),
.B(n_1099),
.Y(n_1216)
);

OAI22x1_ASAP7_75t_L g1217 ( 
.A1(n_1087),
.A2(n_1031),
.B1(n_1099),
.B2(n_1149),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1157),
.B(n_1051),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1152),
.A2(n_1064),
.B(n_1130),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1049),
.B(n_1068),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1124),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1068),
.A2(n_1069),
.B1(n_1130),
.B2(n_1137),
.Y(n_1222)
);

INVx5_ASAP7_75t_L g1223 ( 
.A(n_1119),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1062),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1119),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1113),
.A2(n_1056),
.B(n_1063),
.C(n_1078),
.Y(n_1226)
);

NOR4xp25_ASAP7_75t_L g1227 ( 
.A(n_1119),
.B(n_1088),
.C(n_1090),
.D(n_1103),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1047),
.A2(n_1134),
.B(n_1045),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1095),
.A2(n_888),
.B(n_863),
.C(n_874),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1095),
.A2(n_888),
.B(n_863),
.C(n_874),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1134),
.A2(n_920),
.B(n_970),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1134),
.A2(n_1163),
.B(n_1141),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1047),
.A2(n_1134),
.B(n_1045),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1135),
.A2(n_924),
.A3(n_1132),
.B(n_1072),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1025),
.A2(n_575),
.B(n_585),
.C(n_1022),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1040),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1066),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1025),
.A2(n_734),
.B(n_575),
.C(n_585),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1025),
.A2(n_734),
.B(n_575),
.C(n_585),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1092),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1035),
.B(n_858),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_L g1252 ( 
.A1(n_1025),
.A2(n_708),
.B(n_1022),
.C(n_1027),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1146),
.B(n_993),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1035),
.B(n_734),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1095),
.A2(n_920),
.B1(n_1024),
.B2(n_1022),
.C(n_550),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1025),
.A2(n_877),
.B1(n_787),
.B2(n_803),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1025),
.A2(n_575),
.B(n_585),
.C(n_1022),
.Y(n_1258)
);

AOI21xp33_ASAP7_75t_L g1259 ( 
.A1(n_1025),
.A2(n_787),
.B(n_956),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1040),
.Y(n_1260)
);

OAI22x1_ASAP7_75t_L g1261 ( 
.A1(n_1060),
.A2(n_995),
.B1(n_1138),
.B2(n_1096),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1080),
.B(n_1057),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_SL g1263 ( 
.A1(n_1095),
.A2(n_888),
.B(n_863),
.C(n_874),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1035),
.B(n_734),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1025),
.A2(n_575),
.B(n_585),
.C(n_1022),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1266)
);

AO32x2_ASAP7_75t_L g1267 ( 
.A1(n_1098),
.A2(n_1135),
.A3(n_1132),
.B1(n_1088),
.B2(n_1131),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1025),
.A2(n_877),
.B1(n_787),
.B2(n_803),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1035),
.B(n_858),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1035),
.B(n_734),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1092),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1025),
.A2(n_575),
.B(n_585),
.C(n_1022),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1080),
.B(n_1057),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1035),
.B(n_858),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1279)
);

NOR4xp25_ASAP7_75t_L g1280 ( 
.A(n_1088),
.B(n_1090),
.C(n_1103),
.D(n_1050),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1047),
.A2(n_1134),
.B(n_1045),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1040),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1093),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1025),
.B(n_680),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1066),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1066),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1047),
.A2(n_1134),
.B(n_1045),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1066),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1040),
.Y(n_1292)
);

BUFx2_ASAP7_75t_R g1293 ( 
.A(n_1066),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1163),
.A2(n_1028),
.B(n_1036),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1156),
.A2(n_970),
.B(n_865),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1040),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1035),
.B(n_734),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_SL g1299 ( 
.A1(n_1095),
.A2(n_888),
.B(n_863),
.C(n_874),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1065),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1065),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1146),
.B(n_993),
.Y(n_1302)
);

NOR4xp25_ASAP7_75t_L g1303 ( 
.A(n_1088),
.B(n_1090),
.C(n_1103),
.D(n_1050),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1040),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1025),
.B(n_550),
.C(n_1091),
.Y(n_1305)
);

AOI31xp67_ASAP7_75t_L g1306 ( 
.A1(n_1103),
.A2(n_743),
.A3(n_976),
.B(n_1014),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1194),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1243),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1288),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1249),
.Y(n_1310)
);

OAI21xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1257),
.A2(n_1268),
.B(n_1165),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1180),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1257),
.A2(n_1268),
.B1(n_1259),
.B2(n_1286),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1242),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1305),
.A2(n_1258),
.B1(n_1272),
.B2(n_1240),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1200),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1171),
.A2(n_1261),
.B1(n_1176),
.B2(n_1175),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1172),
.B(n_1265),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1305),
.B1(n_1182),
.B2(n_1197),
.Y(n_1319)
);

BUFx5_ASAP7_75t_L g1320 ( 
.A(n_1198),
.Y(n_1320)
);

CKINVDCx16_ASAP7_75t_R g1321 ( 
.A(n_1287),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1186),
.B(n_1260),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1174),
.A2(n_1165),
.B1(n_1245),
.B2(n_1246),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1282),
.B(n_1292),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1212),
.A2(n_1188),
.B1(n_1192),
.B2(n_1269),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1291),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1174),
.A2(n_1223),
.B1(n_1284),
.B2(n_1241),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1251),
.A2(n_1278),
.B1(n_1213),
.B2(n_1255),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1297),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1304),
.Y(n_1330)
);

INVx3_ASAP7_75t_SL g1331 ( 
.A(n_1185),
.Y(n_1331)
);

CKINVDCx6p67_ASAP7_75t_R g1332 ( 
.A(n_1271),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1187),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1174),
.A2(n_1227),
.B1(n_1303),
.B2(n_1164),
.Y(n_1334)
);

CKINVDCx6p67_ASAP7_75t_R g1335 ( 
.A(n_1287),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1206),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1202),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1223),
.A2(n_1203),
.B1(n_1295),
.B2(n_1284),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1264),
.A2(n_1270),
.B1(n_1298),
.B2(n_1275),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1241),
.A2(n_1244),
.B1(n_1254),
.B2(n_1295),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1179),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1262),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1195),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1183),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1168),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1199),
.B(n_1225),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1191),
.A2(n_1296),
.B1(n_1248),
.B2(n_1244),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1193),
.B(n_1170),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1191),
.A2(n_1296),
.B1(n_1248),
.B2(n_1254),
.Y(n_1350)
);

INVx3_ASAP7_75t_SL g1351 ( 
.A(n_1221),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1181),
.Y(n_1352)
);

CKINVDCx11_ASAP7_75t_R g1353 ( 
.A(n_1198),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1293),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1300),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1301),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1234),
.A2(n_1210),
.B1(n_1204),
.B2(n_1201),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1234),
.A2(n_1217),
.B1(n_1189),
.B2(n_1178),
.Y(n_1358)
);

OAI21xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1227),
.A2(n_1164),
.B(n_1280),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1189),
.A2(n_1211),
.B1(n_1216),
.B2(n_1280),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1211),
.A2(n_1303),
.B1(n_1256),
.B2(n_1166),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1190),
.A2(n_1196),
.B1(n_1215),
.B2(n_1267),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1169),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1199),
.B(n_1224),
.Y(n_1364)
);

BUFx8_ASAP7_75t_SL g1365 ( 
.A(n_1169),
.Y(n_1365)
);

BUFx12f_ASAP7_75t_L g1366 ( 
.A(n_1285),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1285),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1285),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1253),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1220),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1208),
.B(n_1239),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1184),
.A2(n_1302),
.B(n_1253),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1224),
.Y(n_1373)
);

CKINVDCx10_ASAP7_75t_R g1374 ( 
.A(n_1218),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1267),
.A2(n_1167),
.B1(n_1207),
.B2(n_1214),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1236),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1222),
.Y(n_1377)
);

BUFx5_ASAP7_75t_L g1378 ( 
.A(n_1177),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1173),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1219),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1252),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1267),
.A2(n_1167),
.B1(n_1209),
.B2(n_1263),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1173),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1239),
.B(n_1247),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1229),
.A2(n_1250),
.B1(n_1276),
.B2(n_1274),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1236),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1230),
.B(n_1266),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1167),
.A2(n_1273),
.B1(n_1238),
.B2(n_1294),
.Y(n_1388)
);

BUFx4_ASAP7_75t_R g1389 ( 
.A(n_1231),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1232),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1233),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1306),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1299),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1235),
.Y(n_1394)
);

CKINVDCx6p67_ASAP7_75t_R g1395 ( 
.A(n_1226),
.Y(n_1395)
);

CKINVDCx14_ASAP7_75t_R g1396 ( 
.A(n_1277),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1279),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1283),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1289),
.A2(n_1228),
.B1(n_1237),
.B2(n_1281),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1290),
.A2(n_1259),
.B1(n_526),
.B2(n_578),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1259),
.A2(n_526),
.B1(n_578),
.B2(n_1305),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1182),
.A2(n_648),
.B1(n_526),
.B2(n_380),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1259),
.A2(n_526),
.B1(n_578),
.B2(n_1305),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1249),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1200),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1287),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1194),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1200),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1182),
.A2(n_648),
.B1(n_526),
.B2(n_380),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1206),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1257),
.A2(n_1268),
.B1(n_771),
.B2(n_803),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1172),
.B(n_1240),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1194),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1259),
.A2(n_526),
.B1(n_578),
.B2(n_1305),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1251),
.B(n_1269),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1305),
.A2(n_1257),
.B1(n_1268),
.B2(n_1258),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1182),
.A2(n_648),
.B1(n_526),
.B2(n_380),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1257),
.A2(n_1268),
.B1(n_771),
.B2(n_803),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1257),
.A2(n_1268),
.B1(n_771),
.B2(n_803),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1243),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1259),
.A2(n_526),
.B1(n_578),
.B2(n_1305),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1185),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1194),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1185),
.Y(n_1424)
);

BUFx2_ASAP7_75t_R g1425 ( 
.A(n_1212),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1249),
.Y(n_1426)
);

BUFx10_ASAP7_75t_L g1427 ( 
.A(n_1243),
.Y(n_1427)
);

NAND2x1p5_ASAP7_75t_L g1428 ( 
.A(n_1223),
.B(n_1053),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1399),
.A2(n_1385),
.B(n_1388),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1333),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1345),
.B(n_1307),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1333),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1312),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1348),
.B(n_1355),
.Y(n_1434)
);

INVx5_ASAP7_75t_SL g1435 ( 
.A(n_1395),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1356),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1386),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1398),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1348),
.B(n_1416),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1384),
.A2(n_1358),
.B(n_1357),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1416),
.B(n_1350),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1331),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1399),
.A2(n_1388),
.B(n_1387),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1329),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1330),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1376),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1337),
.Y(n_1450)
);

INVxp33_ASAP7_75t_L g1451 ( 
.A(n_1325),
.Y(n_1451)
);

OAI21xp33_ASAP7_75t_L g1452 ( 
.A1(n_1359),
.A2(n_1311),
.B(n_1361),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1370),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1339),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1376),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1371),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1371),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1324),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1394),
.B(n_1382),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1384),
.A2(n_1375),
.B(n_1392),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1349),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1341),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1341),
.B(n_1396),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1344),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1338),
.B(n_1415),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1338),
.B(n_1361),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1360),
.B(n_1362),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1375),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1318),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1358),
.A2(n_1357),
.B(n_1327),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1362),
.A2(n_1315),
.A3(n_1412),
.B(n_1318),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1412),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1360),
.B(n_1327),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1381),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1313),
.A2(n_1315),
.B(n_1323),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1323),
.A2(n_1428),
.B(n_1347),
.Y(n_1477)
);

INVxp33_ASAP7_75t_SL g1478 ( 
.A(n_1354),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1328),
.B(n_1407),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1402),
.A2(n_1409),
.B1(n_1417),
.B2(n_1401),
.Y(n_1480)
);

INVx3_ASAP7_75t_SL g1481 ( 
.A(n_1351),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1391),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1413),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1423),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1322),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1397),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1328),
.B(n_1319),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1342),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1428),
.A2(n_1347),
.B(n_1364),
.Y(n_1489)
);

OAI211xp5_ASAP7_75t_L g1490 ( 
.A1(n_1411),
.A2(n_1419),
.B(n_1418),
.C(n_1414),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1343),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1322),
.B(n_1378),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1378),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1378),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1378),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1364),
.A2(n_1372),
.B(n_1378),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1334),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1390),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1390),
.Y(n_1499)
);

OAI31xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1389),
.A2(n_1417),
.A3(n_1409),
.B(n_1402),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1380),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1393),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1377),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1393),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1369),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1373),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1320),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1400),
.A2(n_1317),
.B(n_1401),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1403),
.A2(n_1414),
.B1(n_1421),
.B2(n_1400),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1403),
.A2(n_1421),
.B1(n_1340),
.B2(n_1351),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1321),
.B(n_1404),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1352),
.A2(n_1346),
.B1(n_1310),
.B2(n_1426),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1437),
.B(n_1406),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1437),
.B(n_1331),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1470),
.B(n_1332),
.Y(n_1515)
);

NOR2x1_ASAP7_75t_SL g1516 ( 
.A(n_1498),
.B(n_1410),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_SL g1517 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1481),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1478),
.B(n_1425),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1444),
.B(n_1425),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1481),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1485),
.B(n_1335),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1464),
.B(n_1427),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1436),
.B(n_1308),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1509),
.A2(n_1368),
.B1(n_1366),
.B2(n_1363),
.Y(n_1525)
);

AND2x4_ASAP7_75t_SL g1526 ( 
.A(n_1439),
.B(n_1420),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1500),
.A2(n_1336),
.B(n_1316),
.C(n_1405),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1501),
.B(n_1353),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1440),
.A2(n_1408),
.B(n_1326),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1309),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1434),
.B(n_1365),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1475),
.B(n_1374),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1480),
.A2(n_1508),
.B1(n_1459),
.B2(n_1510),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1481),
.Y(n_1534)
);

AO32x2_ASAP7_75t_L g1535 ( 
.A1(n_1453),
.A2(n_1367),
.A3(n_1434),
.B1(n_1472),
.B2(n_1479),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1452),
.A2(n_1440),
.B(n_1443),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1490),
.A2(n_1452),
.B1(n_1467),
.B2(n_1497),
.Y(n_1537)
);

NOR3xp33_ASAP7_75t_SL g1538 ( 
.A(n_1499),
.B(n_1504),
.C(n_1502),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1459),
.A2(n_1467),
.B(n_1443),
.C(n_1468),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1466),
.B(n_1459),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_SL g1541 ( 
.A1(n_1502),
.A2(n_1504),
.B(n_1497),
.C(n_1511),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1441),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1459),
.A2(n_1468),
.B(n_1474),
.C(n_1463),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1463),
.A2(n_1474),
.B(n_1473),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1446),
.A2(n_1429),
.B(n_1471),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1487),
.A2(n_1435),
.B1(n_1469),
.B2(n_1476),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1477),
.A2(n_1446),
.B(n_1496),
.Y(n_1548)
);

AO32x2_ASAP7_75t_L g1549 ( 
.A1(n_1472),
.A2(n_1479),
.A3(n_1492),
.B1(n_1469),
.B2(n_1488),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1506),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1439),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1433),
.Y(n_1552)
);

INVxp33_ASAP7_75t_L g1553 ( 
.A(n_1451),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1487),
.A2(n_1471),
.B(n_1477),
.C(n_1476),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1458),
.B(n_1506),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1482),
.A2(n_1461),
.B(n_1462),
.C(n_1486),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1431),
.Y(n_1557)
);

NAND2x1_ASAP7_75t_L g1558 ( 
.A(n_1461),
.B(n_1462),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1445),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1472),
.B(n_1456),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1483),
.A2(n_1484),
.B1(n_1465),
.B2(n_1435),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1442),
.A2(n_1486),
.B(n_1489),
.Y(n_1562)
);

OAI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1512),
.A2(n_1472),
.B(n_1442),
.C(n_1430),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1472),
.B(n_1456),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1442),
.A2(n_1489),
.B(n_1457),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1438),
.B(n_1507),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1536),
.A2(n_1442),
.B1(n_1460),
.B2(n_1488),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1560),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1560),
.B(n_1472),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1564),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1493),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1564),
.B(n_1447),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1559),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1549),
.B(n_1494),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1546),
.B(n_1545),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1546),
.B(n_1495),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1536),
.A2(n_1491),
.B1(n_1435),
.B2(n_1483),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1537),
.A2(n_1450),
.B1(n_1447),
.B2(n_1454),
.C(n_1448),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1535),
.B(n_1555),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1535),
.B(n_1455),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1535),
.B(n_1455),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1563),
.B(n_1448),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1540),
.B(n_1449),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1533),
.A2(n_1491),
.B1(n_1435),
.B2(n_1484),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1556),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1566),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1565),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1562),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1550),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1565),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1566),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1537),
.A2(n_1435),
.B1(n_1465),
.B2(n_1450),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1430),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1569),
.B(n_1544),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1577),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1593),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1588),
.A2(n_1539),
.B1(n_1543),
.B2(n_1538),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1584),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1576),
.B(n_1514),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1584),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1573),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1513),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1573),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1588),
.B(n_1518),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1569),
.B(n_1557),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1573),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1593),
.B(n_1515),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1569),
.B(n_1554),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1572),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1576),
.B(n_1513),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1576),
.B(n_1580),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1523),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1569),
.B(n_1432),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1572),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1529),
.C(n_1541),
.Y(n_1623)
);

INVxp67_ASAP7_75t_SL g1624 ( 
.A(n_1592),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1574),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1517),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1580),
.B(n_1522),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1579),
.A2(n_1516),
.B(n_1547),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_R g1629 ( 
.A(n_1597),
.B(n_1521),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1583),
.Y(n_1630)
);

INVx5_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1594),
.A2(n_1547),
.B1(n_1527),
.B2(n_1529),
.C(n_1525),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1583),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1581),
.B(n_1534),
.Y(n_1634)
);

AND2x4_ASAP7_75t_SL g1635 ( 
.A(n_1596),
.B(n_1534),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1595),
.B(n_1586),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1596),
.B(n_1551),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1618),
.B(n_1636),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1601),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1621),
.B(n_1570),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1615),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1623),
.B(n_1596),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1570),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1618),
.B(n_1581),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1600),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1600),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1636),
.B(n_1581),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1602),
.A2(n_1579),
.B1(n_1567),
.B2(n_1587),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1620),
.B(n_1568),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1605),
.B(n_1619),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1631),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1620),
.B(n_1594),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1607),
.B(n_1571),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1610),
.B(n_1531),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1615),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1605),
.B(n_1581),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1616),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1622),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1619),
.B(n_1582),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1622),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1530),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1614),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1625),
.Y(n_1667)
);

NOR2xp67_ASAP7_75t_L g1668 ( 
.A(n_1631),
.B(n_1592),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1629),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1582),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1628),
.A2(n_1578),
.B1(n_1587),
.B2(n_1579),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1608),
.B(n_1617),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1617),
.B(n_1582),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1582),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1607),
.B(n_1571),
.Y(n_1675)
);

INVx3_ASAP7_75t_SL g1676 ( 
.A(n_1669),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1667),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1645),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1639),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1665),
.B(n_1599),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1665),
.B(n_1599),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1651),
.B(n_1672),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1648),
.B(n_1614),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1648),
.B(n_1611),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1651),
.B(n_1634),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_SL g1686 ( 
.A(n_1642),
.B(n_1528),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1669),
.B(n_1519),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1667),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1611),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1641),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1642),
.B(n_1571),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1651),
.B(n_1634),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1571),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1641),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1645),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1657),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1657),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1658),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1640),
.B(n_1609),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1664),
.B(n_1628),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1640),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1645),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1658),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1646),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1638),
.B(n_1662),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1660),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1643),
.B(n_1654),
.Y(n_1709)
);

OAI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1671),
.A2(n_1585),
.B1(n_1637),
.B2(n_1598),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1711)
);

AND3x2_ASAP7_75t_L g1712 ( 
.A(n_1656),
.B(n_1520),
.C(n_1532),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1660),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1643),
.B(n_1575),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1654),
.B(n_1575),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1653),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1654),
.B(n_1609),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1650),
.B(n_1612),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1656),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1676),
.B(n_1719),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1676),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1682),
.B(n_1662),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1662),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1612),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1676),
.Y(n_1726)
);

AOI33xp33_ASAP7_75t_L g1727 ( 
.A1(n_1710),
.A2(n_1644),
.A3(n_1597),
.B1(n_1674),
.B2(n_1567),
.B3(n_1659),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1690),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1701),
.A2(n_1671),
.B(n_1598),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1681),
.B(n_1650),
.Y(n_1730)
);

INVxp67_ASAP7_75t_SL g1731 ( 
.A(n_1701),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1686),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1695),
.B(n_1644),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1690),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1695),
.B(n_1644),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1705),
.B(n_1707),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1702),
.B(n_1647),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1681),
.B(n_1650),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1683),
.B(n_1653),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1686),
.B(n_1680),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1687),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1684),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1679),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1686),
.B(n_1691),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1716),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1694),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1716),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1705),
.B(n_1659),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1716),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1709),
.B(n_1647),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1694),
.Y(n_1751)
);

AND2x4_ASAP7_75t_SL g1752 ( 
.A(n_1685),
.B(n_1532),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1707),
.B(n_1659),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1677),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1697),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1709),
.B(n_1689),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1685),
.B(n_1670),
.Y(n_1757)
);

OAI32xp33_ASAP7_75t_L g1758 ( 
.A1(n_1740),
.A2(n_1693),
.A3(n_1714),
.B1(n_1715),
.B2(n_1688),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1729),
.B(n_1653),
.Y(n_1759)
);

O2A1O1Ixp33_ASAP7_75t_SL g1760 ( 
.A1(n_1726),
.A2(n_1677),
.B(n_1688),
.C(n_1524),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1746),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1731),
.A2(n_1668),
.B(n_1632),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1746),
.Y(n_1763)
);

AOI33xp33_ASAP7_75t_L g1764 ( 
.A1(n_1726),
.A2(n_1698),
.A3(n_1713),
.B1(n_1697),
.B2(n_1708),
.B3(n_1699),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1752),
.Y(n_1765)
);

XNOR2x1_ASAP7_75t_L g1766 ( 
.A(n_1740),
.B(n_1530),
.Y(n_1766)
);

OR4x1_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1704),
.C(n_1698),
.D(n_1699),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1751),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1741),
.A2(n_1668),
.B(n_1598),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1732),
.A2(n_1635),
.B(n_1674),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1722),
.B(n_1633),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1732),
.A2(n_1585),
.B(n_1711),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1744),
.A2(n_1692),
.B1(n_1711),
.B2(n_1720),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1721),
.B(n_1647),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1742),
.A2(n_1727),
.B(n_1737),
.C(n_1730),
.Y(n_1775)
);

O2A1O1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1739),
.A2(n_1704),
.B(n_1713),
.C(n_1708),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1752),
.B(n_1692),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1751),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1743),
.B(n_1700),
.Y(n_1779)
);

OAI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1739),
.A2(n_1585),
.B1(n_1637),
.B2(n_1591),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1733),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1739),
.A2(n_1591),
.B1(n_1594),
.B2(n_1585),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1756),
.B(n_1700),
.Y(n_1783)
);

AOI21xp33_ASAP7_75t_SL g1784 ( 
.A1(n_1759),
.A2(n_1739),
.B(n_1749),
.Y(n_1784)
);

OAI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1759),
.A2(n_1747),
.B(n_1745),
.C(n_1734),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1761),
.Y(n_1786)
);

O2A1O1Ixp5_ASAP7_75t_L g1787 ( 
.A1(n_1762),
.A2(n_1745),
.B(n_1734),
.C(n_1728),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1763),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1776),
.A2(n_1739),
.B(n_1754),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1768),
.Y(n_1790)
);

OAI32xp33_ASAP7_75t_L g1791 ( 
.A1(n_1782),
.A2(n_1730),
.A3(n_1738),
.B1(n_1745),
.B2(n_1754),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1778),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1764),
.B(n_1747),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1779),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1782),
.A2(n_1738),
.B1(n_1725),
.B2(n_1750),
.C(n_1678),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1775),
.A2(n_1755),
.B(n_1736),
.Y(n_1796)
);

NAND2x1_ASAP7_75t_SL g1797 ( 
.A(n_1771),
.B(n_1755),
.Y(n_1797)
);

AO22x1_ASAP7_75t_L g1798 ( 
.A1(n_1771),
.A2(n_1736),
.B1(n_1723),
.B2(n_1724),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1775),
.A2(n_1703),
.B1(n_1696),
.B2(n_1706),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1774),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1777),
.B(n_1781),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1772),
.A2(n_1724),
.B(n_1723),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1767),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1797),
.B(n_1765),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1799),
.A2(n_1780),
.B1(n_1766),
.B2(n_1760),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1786),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1787),
.A2(n_1760),
.B(n_1780),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1801),
.B(n_1783),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1800),
.B(n_1748),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1800),
.B(n_1801),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1788),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1798),
.B(n_1748),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1797),
.Y(n_1813)
);

AOI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1791),
.A2(n_1758),
.B(n_1769),
.C(n_1770),
.Y(n_1814)
);

AOI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1807),
.A2(n_1789),
.B(n_1784),
.C(n_1796),
.Y(n_1815)
);

OAI211xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1814),
.A2(n_1785),
.B(n_1793),
.C(n_1803),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1813),
.A2(n_1803),
.B1(n_1795),
.B2(n_1794),
.C(n_1792),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_SL g1818 ( 
.A(n_1805),
.B(n_1790),
.C(n_1773),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1808),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1810),
.B(n_1802),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1809),
.B(n_1733),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1804),
.A2(n_1678),
.B1(n_1706),
.B2(n_1703),
.Y(n_1822)
);

NAND4xp25_ASAP7_75t_L g1823 ( 
.A(n_1804),
.B(n_1753),
.C(n_1757),
.D(n_1735),
.Y(n_1823)
);

NAND3xp33_ASAP7_75t_L g1824 ( 
.A(n_1806),
.B(n_1753),
.C(n_1757),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1811),
.A2(n_1696),
.B(n_1678),
.Y(n_1825)
);

NAND3x1_ASAP7_75t_L g1826 ( 
.A(n_1819),
.B(n_1817),
.C(n_1821),
.Y(n_1826)
);

O2A1O1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1816),
.A2(n_1815),
.B(n_1820),
.C(n_1818),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1824),
.Y(n_1828)
);

AOI21xp33_ASAP7_75t_L g1829 ( 
.A1(n_1822),
.A2(n_1812),
.B(n_1703),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1823),
.A2(n_1825),
.B1(n_1706),
.B2(n_1696),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1819),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_SL g1832 ( 
.A(n_1827),
.B(n_1735),
.C(n_1720),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1831),
.B(n_1630),
.Y(n_1833)
);

NOR4xp25_ASAP7_75t_L g1834 ( 
.A(n_1826),
.B(n_1718),
.C(n_1717),
.D(n_1542),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_L g1835 ( 
.A1(n_1829),
.A2(n_1674),
.B(n_1718),
.C(n_1717),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1828),
.A2(n_1553),
.B1(n_1674),
.B2(n_1591),
.C(n_1655),
.Y(n_1836)
);

AOI311xp33_ASAP7_75t_L g1837 ( 
.A1(n_1830),
.A2(n_1661),
.A3(n_1663),
.B(n_1666),
.C(n_1613),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1832),
.B(n_1674),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_L g1839 ( 
.A(n_1833),
.B(n_1633),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1834),
.B(n_1633),
.Y(n_1840)
);

XOR2x2_ASAP7_75t_L g1841 ( 
.A(n_1835),
.B(n_1637),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1836),
.Y(n_1842)
);

AOI322xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1838),
.A3(n_1839),
.B1(n_1840),
.B2(n_1837),
.C1(n_1841),
.C2(n_1591),
.Y(n_1843)
);

AOI211x1_ASAP7_75t_L g1844 ( 
.A1(n_1842),
.A2(n_1649),
.B(n_1652),
.C(n_1655),
.Y(n_1844)
);

AND4x1_ASAP7_75t_L g1845 ( 
.A(n_1839),
.B(n_1578),
.C(n_1673),
.D(n_1670),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1845),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1846),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1847),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1847),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1848),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1846),
.B1(n_1844),
.B2(n_1843),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1851),
.A2(n_1630),
.B1(n_1631),
.B2(n_1627),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1852),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1853),
.B(n_1850),
.Y(n_1854)
);

XNOR2xp5_ASAP7_75t_L g1855 ( 
.A(n_1854),
.B(n_1526),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_R g1856 ( 
.A1(n_1855),
.A2(n_1603),
.B1(n_1631),
.B2(n_1675),
.C(n_1606),
.Y(n_1856)
);

AOI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1551),
.B(n_1649),
.C(n_1652),
.Y(n_1857)
);


endmodule