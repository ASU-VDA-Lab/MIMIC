module real_jpeg_30155_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_42),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_42),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_4),
.A2(n_9),
.B1(n_42),
.B2(n_65),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_39),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_44),
.B1(n_67),
.B2(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_8),
.A2(n_9),
.B1(n_44),
.B2(n_65),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_9),
.B(n_64),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_8),
.A2(n_10),
.B(n_37),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_8),
.B(n_62),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_8),
.A2(n_22),
.B(n_38),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_76),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_9),
.A2(n_10),
.B1(n_65),
.B2(n_77),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_9),
.A2(n_44),
.B(n_123),
.C(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_113),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_112),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_98),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_16),
.B(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_83),
.B2(n_97),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_21),
.A2(n_29),
.B1(n_53),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_21),
.B(n_24),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_27),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_29),
.A2(n_50),
.B(n_91),
.Y(n_136)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_29),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_32),
.A2(n_33),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_32),
.A2(n_33),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_33),
.B(n_90),
.C(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_33),
.B(n_130),
.C(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_34),
.B(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_37),
.A2(n_39),
.B(n_44),
.C(n_147),
.Y(n_146)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_40),
.B(n_44),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_63),
.B(n_68),
.C(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_44),
.B(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_59),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_54),
.B1(n_55),
.B2(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_55),
.B1(n_146),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_54),
.A2(n_55),
.B1(n_106),
.B2(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_120),
.C(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_55),
.B(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B(n_58),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_73),
.B1(n_74),
.B2(n_82),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_106),
.C(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_60),
.A2(n_82),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_69),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_70),
.B1(n_71),
.B2(n_85),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_72)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.C(n_92),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_92),
.B1(n_93),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_90),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_90),
.B(n_165),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_93),
.B1(n_132),
.B2(n_137),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_93),
.B(n_133),
.C(n_136),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_96),
.B(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.C(n_104),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_99),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_190),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_185),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_175),
.B(n_184),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_142),
.B(n_174),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_119),
.B(n_129),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_132),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_169),
.B(n_173),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_154),
.B(n_168),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B(n_167),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_166),
.Y(n_158)
);

INVx5_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_177),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);


endmodule