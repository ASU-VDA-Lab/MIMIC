module fake_jpeg_31467_n_111 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_4),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_23),
.B(n_16),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_20),
.B1(n_19),
.B2(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_29),
.B1(n_0),
.B2(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_17),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_20),
.B1(n_13),
.B2(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_51),
.B1(n_27),
.B2(n_29),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_20),
.B1(n_19),
.B2(n_12),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_36),
.B1(n_32),
.B2(n_37),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_68),
.B1(n_44),
.B2(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_11),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_66),
.B1(n_49),
.B2(n_63),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_9),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_43),
.B(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_47),
.B1(n_49),
.B2(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_44),
.B1(n_55),
.B2(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_82),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_89),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_63),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_71),
.C(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_77),
.C(n_82),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_60),
.B(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_76),
.B1(n_80),
.B2(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_88),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_92),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_93),
.C(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_94),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_105),
.Y(n_106)
);

AOI211xp5_ASAP7_75t_SL g108 ( 
.A1(n_106),
.A2(n_107),
.B(n_104),
.C(n_103),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_104),
.B(n_106),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_60),
.A3(n_79),
.B1(n_105),
.B2(n_108),
.C(n_107),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_110),
.Y(n_111)
);


endmodule