module real_aes_7423_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_884;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_767;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp5_ASAP7_75t_SL g443 ( .A1(n_0), .A2(n_244), .B1(n_360), .B2(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_1), .A2(n_274), .B1(n_342), .B2(n_350), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_2), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_3), .A2(n_253), .B1(n_707), .B2(n_795), .Y(n_794) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_4), .A2(n_90), .B1(n_264), .B2(n_320), .C1(n_326), .C2(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_5), .A2(n_121), .B1(n_405), .B2(n_481), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_6), .A2(n_24), .B1(n_410), .B2(n_455), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_7), .A2(n_64), .B1(n_332), .B2(n_540), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_8), .B(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_9), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_10), .A2(n_132), .B1(n_683), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_11), .A2(n_76), .B1(n_772), .B2(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g522 ( .A(n_12), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_13), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_14), .A2(n_133), .B1(n_591), .B2(n_654), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_15), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_16), .A2(n_270), .B1(n_477), .B2(n_790), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_17), .A2(n_151), .B1(n_548), .B2(n_657), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_18), .A2(n_127), .B1(n_426), .B2(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_19), .A2(n_57), .B1(n_423), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_20), .A2(n_119), .B1(n_335), .B2(n_479), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_21), .A2(n_161), .B1(n_331), .B2(n_335), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_22), .A2(n_176), .B1(n_382), .B2(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g393 ( .A(n_23), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_25), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_26), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_27), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_28), .A2(n_172), .B1(n_470), .B2(n_585), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_29), .A2(n_278), .B1(n_655), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_30), .A2(n_245), .B1(n_405), .B2(n_406), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_31), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_32), .A2(n_128), .B1(n_365), .B2(n_371), .Y(n_621) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_33), .A2(n_92), .B1(n_307), .B2(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g836 ( .A(n_33), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_34), .B(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_35), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_36), .A2(n_219), .B1(n_320), .B2(n_455), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_37), .A2(n_162), .B1(n_426), .B2(n_429), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_38), .A2(n_165), .B1(n_441), .B2(n_446), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_39), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_40), .A2(n_263), .B1(n_378), .B2(n_424), .Y(n_680) );
INVx1_ASAP7_75t_L g693 ( .A(n_41), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_42), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_43), .A2(n_130), .B1(n_423), .B2(n_428), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_44), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_45), .A2(n_254), .B1(n_418), .B2(n_428), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_46), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_47), .Y(n_541) );
INVx1_ASAP7_75t_L g677 ( .A(n_48), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_49), .Y(n_630) );
AO22x2_ASAP7_75t_L g310 ( .A1(n_50), .A2(n_95), .B1(n_307), .B2(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g837 ( .A(n_50), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_51), .A2(n_138), .B1(n_327), .B2(n_338), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_52), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_53), .A2(n_149), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_54), .A2(n_178), .B1(n_332), .B2(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_55), .A2(n_275), .B1(n_343), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_56), .A2(n_164), .B1(n_446), .B2(n_447), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_58), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_59), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_60), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_61), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_62), .A2(n_260), .B1(n_319), .B2(n_326), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g819 ( .A1(n_63), .A2(n_195), .B1(n_269), .B2(n_320), .C1(n_483), .C2(n_543), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_65), .Y(n_770) );
AOI22xp5_ASAP7_75t_SL g439 ( .A1(n_66), .A2(n_158), .B1(n_440), .B2(n_441), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_67), .A2(n_261), .B1(n_423), .B2(n_424), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_68), .A2(n_272), .B1(n_697), .B2(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_69), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_70), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_71), .A2(n_233), .B1(n_463), .B2(n_465), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_72), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_73), .A2(n_281), .B1(n_587), .B2(n_588), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_74), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_75), .A2(n_199), .B1(n_371), .B2(n_470), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_77), .A2(n_188), .B1(n_447), .B2(n_657), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_78), .A2(n_204), .B1(n_588), .B2(n_657), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_79), .A2(n_197), .B1(n_335), .B2(n_479), .Y(n_628) );
AOI22xp5_ASAP7_75t_SL g438 ( .A1(n_80), .A2(n_146), .B1(n_420), .B2(n_424), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_81), .A2(n_232), .B1(n_343), .B2(n_352), .Y(n_456) );
XNOR2x2_ASAP7_75t_L g459 ( .A(n_82), .B(n_460), .Y(n_459) );
AO22x2_ASAP7_75t_L g560 ( .A1(n_83), .A2(n_561), .B1(n_592), .B2(n_593), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_83), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_84), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_85), .A2(n_242), .B1(n_584), .B2(n_585), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_86), .Y(n_532) );
AOI211xp5_ASAP7_75t_L g529 ( .A1(n_87), .A2(n_530), .B(n_531), .C(n_537), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_88), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_89), .A2(n_152), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g686 ( .A(n_91), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_93), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_94), .A2(n_144), .B1(n_410), .B2(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_96), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_97), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_98), .A2(n_210), .B1(n_358), .B2(n_429), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_99), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_100), .Y(n_820) );
AND2x2_ASAP7_75t_L g293 ( .A(n_101), .B(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_SL g688 ( .A1(n_102), .A2(n_689), .B1(n_716), .B2(n_717), .Y(n_688) );
INVx1_ASAP7_75t_L g717 ( .A(n_102), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_103), .A2(n_782), .B1(n_802), .B2(n_803), .Y(n_781) );
INVx1_ASAP7_75t_L g803 ( .A(n_103), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_104), .A2(n_134), .B1(n_383), .B2(n_385), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_105), .A2(n_208), .B1(n_657), .B2(n_658), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_106), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_107), .A2(n_213), .B1(n_405), .B2(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_108), .A2(n_212), .B1(n_426), .B2(n_548), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_109), .A2(n_840), .B1(n_865), .B2(n_866), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_109), .Y(n_865) );
INVx1_ASAP7_75t_L g290 ( .A(n_110), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_111), .A2(n_171), .B1(n_661), .B2(n_662), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_112), .A2(n_150), .B1(n_320), .B2(n_327), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_113), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g374 ( .A1(n_114), .A2(n_249), .B1(n_375), .B2(n_378), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_115), .A2(n_192), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_116), .A2(n_248), .B1(n_424), .B2(n_901), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_117), .B(n_650), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_118), .A2(n_236), .B1(n_612), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g497 ( .A(n_120), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_122), .A2(n_166), .B1(n_735), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_123), .A2(n_229), .B1(n_420), .B2(n_423), .Y(n_897) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_124), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_125), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_126), .A2(n_155), .B1(n_371), .B2(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_129), .A2(n_247), .B1(n_428), .B2(n_440), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_131), .A2(n_231), .B1(n_356), .B2(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g523 ( .A(n_135), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_136), .A2(n_211), .B1(n_712), .B2(n_861), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_137), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_139), .A2(n_186), .B1(n_338), .B2(n_405), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_140), .A2(n_222), .B1(n_331), .B2(n_335), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_141), .A2(n_279), .B1(n_365), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_142), .A2(n_167), .B1(n_385), .B2(n_418), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_143), .Y(n_847) );
AOI22xp5_ASAP7_75t_SL g743 ( .A1(n_145), .A2(n_744), .B1(n_774), .B2(n_775), .Y(n_743) );
INVx1_ASAP7_75t_L g775 ( .A(n_145), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_147), .B(n_477), .Y(n_535) );
INVx2_ASAP7_75t_L g294 ( .A(n_148), .Y(n_294) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_153), .A2(n_183), .B1(n_365), .B2(n_371), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_154), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_156), .A2(n_217), .B1(n_479), .B2(n_481), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_157), .Y(n_747) );
AND2x6_ASAP7_75t_L g289 ( .A(n_159), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_159), .Y(n_830) );
AO22x2_ASAP7_75t_L g314 ( .A1(n_160), .A2(n_240), .B1(n_307), .B2(n_311), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_163), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_168), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_169), .A2(n_209), .B1(n_378), .B2(n_420), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_170), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_173), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_174), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_175), .A2(n_268), .B1(n_446), .B2(n_658), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_177), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_179), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_180), .A2(n_191), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_181), .A2(n_287), .B(n_295), .C(n_838), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_182), .A2(n_604), .B1(n_635), .B2(n_636), .Y(n_603) );
INVx1_ASAP7_75t_L g635 ( .A(n_182), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_184), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_185), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_187), .A2(n_225), .B1(n_356), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_189), .A2(n_266), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_190), .A2(n_257), .B1(n_654), .B2(n_655), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_193), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_194), .Y(n_742) );
AO22x2_ASAP7_75t_L g316 ( .A1(n_196), .A2(n_255), .B1(n_307), .B2(n_308), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_198), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_200), .A2(n_228), .B1(n_385), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_201), .A2(n_258), .B1(n_543), .B2(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_202), .Y(n_886) );
INVx1_ASAP7_75t_L g557 ( .A(n_203), .Y(n_557) );
INVx1_ASAP7_75t_L g494 ( .A(n_205), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g876 ( .A(n_206), .Y(n_876) );
AOI22xp5_ASAP7_75t_SL g880 ( .A1(n_206), .A2(n_876), .B1(n_881), .B2(n_902), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_207), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_214), .A2(n_282), .B1(n_406), .B2(n_633), .Y(n_678) );
INVx1_ASAP7_75t_L g692 ( .A(n_215), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_216), .Y(n_893) );
INVx1_ASAP7_75t_L g519 ( .A(n_218), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_220), .B(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_221), .A2(n_259), .B1(n_420), .B2(n_441), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_223), .B(n_444), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_224), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_226), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_227), .A2(n_256), .B1(n_429), .B2(n_584), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_230), .A2(n_276), .B1(n_385), .B2(n_418), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_234), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_235), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_237), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_238), .A2(n_246), .B1(n_682), .B2(n_683), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_239), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_240), .B(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_241), .B(n_650), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_243), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_250), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_251), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_252), .A2(n_262), .B1(n_477), .B2(n_650), .Y(n_813) );
INVx1_ASAP7_75t_L g833 ( .A(n_255), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_265), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_267), .A2(n_285), .B1(n_382), .B2(n_385), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_271), .Y(n_848) );
INVx1_ASAP7_75t_L g307 ( .A(n_273), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_273), .Y(n_309) );
INVx1_ASAP7_75t_L g398 ( .A(n_277), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_280), .A2(n_284), .B1(n_801), .B2(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_283), .Y(n_644) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_290), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g874 ( .A1(n_291), .A2(n_828), .B(n_875), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_600), .B1(n_823), .B2(n_824), .C(n_825), .Y(n_295) );
INVx1_ASAP7_75t_L g823 ( .A(n_296), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_388), .B1(n_598), .B2(n_599), .Y(n_296) );
INVx1_ASAP7_75t_L g598 ( .A(n_297), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_354), .C(n_373), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_329), .Y(n_300) );
OAI21xp5_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_317), .B(n_318), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_SL g403 ( .A(n_303), .Y(n_403) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g451 ( .A(n_304), .Y(n_451) );
INVx4_ASAP7_75t_L g484 ( .A(n_304), .Y(n_484) );
INVx2_ASAP7_75t_SL g501 ( .A(n_304), .Y(n_501) );
BUFx3_ASAP7_75t_L g530 ( .A(n_304), .Y(n_530) );
INVx2_ASAP7_75t_L g645 ( .A(n_304), .Y(n_645) );
AND2x6_ASAP7_75t_L g304 ( .A(n_305), .B(n_312), .Y(n_304) );
AND2x4_ASAP7_75t_L g338 ( .A(n_305), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g579 ( .A(n_305), .Y(n_579) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_310), .Y(n_305) );
AND2x2_ASAP7_75t_L g325 ( .A(n_306), .B(n_314), .Y(n_325) );
INVx2_ASAP7_75t_L g349 ( .A(n_306), .Y(n_349) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_309), .Y(n_311) );
INVx2_ASAP7_75t_L g324 ( .A(n_310), .Y(n_324) );
INVx1_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
OR2x2_ASAP7_75t_L g348 ( .A(n_310), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g353 ( .A(n_310), .B(n_349), .Y(n_353) );
AND2x6_ASAP7_75t_L g377 ( .A(n_312), .B(n_347), .Y(n_377) );
AND2x4_ASAP7_75t_L g380 ( .A(n_312), .B(n_353), .Y(n_380) );
AND2x2_ASAP7_75t_L g384 ( .A(n_312), .B(n_359), .Y(n_384) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
AND2x2_ASAP7_75t_L g346 ( .A(n_313), .B(n_316), .Y(n_346) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_314), .B(n_316), .Y(n_363) );
AND2x2_ASAP7_75t_L g370 ( .A(n_314), .B(n_340), .Y(n_370) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g323 ( .A(n_316), .Y(n_323) );
INVx1_ASAP7_75t_L g340 ( .A(n_316), .Y(n_340) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g503 ( .A(n_320), .Y(n_503) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx4f_ASAP7_75t_SL g410 ( .A(n_321), .Y(n_410) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_321), .Y(n_540) );
BUFx2_ASAP7_75t_L g572 ( .A(n_321), .Y(n_572) );
BUFx6f_ASAP7_75t_L g890 ( .A(n_321), .Y(n_890) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g328 ( .A(n_323), .Y(n_328) );
AND2x2_ASAP7_75t_L g359 ( .A(n_324), .B(n_349), .Y(n_359) );
INVx1_ASAP7_75t_L g414 ( .A(n_324), .Y(n_414) );
AND2x4_ASAP7_75t_L g327 ( .A(n_325), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g332 ( .A(n_325), .B(n_333), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_325), .B(n_414), .Y(n_413) );
BUFx4f_ASAP7_75t_L g752 ( .A(n_326), .Y(n_752) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx12f_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_327), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_341), .Y(n_329) );
BUFx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g455 ( .A(n_332), .Y(n_455) );
INVx1_ASAP7_75t_L g480 ( .A(n_332), .Y(n_480) );
BUFx2_ASAP7_75t_L g815 ( .A(n_332), .Y(n_815) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x6_ASAP7_75t_L g372 ( .A(n_334), .B(n_363), .Y(n_372) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_SL g406 ( .A(n_338), .Y(n_406) );
BUFx2_ASAP7_75t_SL g481 ( .A(n_338), .Y(n_481) );
BUFx3_ASAP7_75t_L g735 ( .A(n_338), .Y(n_735) );
INVx1_ASAP7_75t_L g580 ( .A(n_339), .Y(n_580) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx5_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g477 ( .A(n_344), .Y(n_477) );
INVx2_ASAP7_75t_L g673 ( .A(n_344), .Y(n_673) );
INVx2_ASAP7_75t_L g733 ( .A(n_344), .Y(n_733) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AND2x6_ASAP7_75t_L g352 ( .A(n_346), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g358 ( .A(n_346), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g400 ( .A(n_346), .B(n_353), .Y(n_400) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g396 ( .A(n_348), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
BUFx4f_ASAP7_75t_L g650 ( .A(n_352), .Y(n_650) );
BUFx2_ASAP7_75t_L g790 ( .A(n_352), .Y(n_790) );
AND2x2_ASAP7_75t_L g369 ( .A(n_353), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_353), .B(n_370), .Y(n_517) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_364), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_357), .A2(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g856 ( .A(n_357), .Y(n_856) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
BUFx3_ASAP7_75t_L g447 ( .A(n_358), .Y(n_447) );
BUFx3_ASAP7_75t_L g588 ( .A(n_358), .Y(n_588) );
BUFx3_ASAP7_75t_L g682 ( .A(n_358), .Y(n_682) );
AND2x4_ASAP7_75t_L g361 ( .A(n_359), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_370), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_359), .B(n_370), .Y(n_520) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_SL g418 ( .A(n_361), .Y(n_418) );
INVx1_ASAP7_75t_L g515 ( .A(n_361), .Y(n_515) );
BUFx2_ASAP7_75t_L g548 ( .A(n_361), .Y(n_548) );
BUFx3_ASAP7_75t_L g591 ( .A(n_361), .Y(n_591) );
BUFx3_ASAP7_75t_L g655 ( .A(n_361), .Y(n_655) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_361), .Y(n_707) );
BUFx3_ASAP7_75t_L g761 ( .A(n_361), .Y(n_761) );
AND2x2_ASAP7_75t_L g444 ( .A(n_362), .B(n_414), .Y(n_444) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx4_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
INVx1_ASAP7_75t_L g470 ( .A(n_368), .Y(n_470) );
INVx2_ASAP7_75t_L g584 ( .A(n_368), .Y(n_584) );
INVx5_ASAP7_75t_L g662 ( .A(n_368), .Y(n_662) );
BUFx3_ASAP7_75t_L g710 ( .A(n_368), .Y(n_710) );
INVx8_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx6_ASAP7_75t_SL g429 ( .A(n_372), .Y(n_429) );
INVx1_ASAP7_75t_L g471 ( .A(n_372), .Y(n_471) );
INVx1_ASAP7_75t_SL g683 ( .A(n_372), .Y(n_683) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_381), .Y(n_373) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx3_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
INVx2_ASAP7_75t_SL g712 ( .A(n_376), .Y(n_712) );
INVx11_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx11_ASAP7_75t_L g464 ( .A(n_377), .Y(n_464) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g423 ( .A(n_379), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g508 ( .A1(n_379), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_379), .A2(n_551), .B1(n_552), .B2(n_553), .Y(n_550) );
INVx3_ASAP7_75t_L g661 ( .A(n_379), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_379), .A2(n_765), .B1(n_766), .B2(n_768), .Y(n_764) );
INVx2_ASAP7_75t_L g861 ( .A(n_379), .Y(n_861) );
INVx6_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g441 ( .A(n_380), .Y(n_441) );
BUFx3_ASAP7_75t_L g465 ( .A(n_380), .Y(n_465) );
INVx1_ASAP7_75t_SL g556 ( .A(n_382), .Y(n_556) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g612 ( .A(n_383), .Y(n_612) );
INVx3_ASAP7_75t_L g715 ( .A(n_383), .Y(n_715) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_SL g440 ( .A(n_384), .Y(n_440) );
INVx2_ASAP7_75t_L g509 ( .A(n_384), .Y(n_509) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_384), .Y(n_772) );
BUFx4f_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g614 ( .A(n_386), .Y(n_614) );
BUFx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g446 ( .A(n_387), .Y(n_446) );
BUFx3_ASAP7_75t_L g654 ( .A(n_387), .Y(n_654) );
BUFx3_ASAP7_75t_L g797 ( .A(n_387), .Y(n_797) );
INVx1_ASAP7_75t_L g599 ( .A(n_388), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_431), .B1(n_596), .B2(n_597), .Y(n_388) );
INVx1_ASAP7_75t_SL g596 ( .A(n_389), .Y(n_596) );
XNOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_430), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_415), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_401), .C(n_407), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_398), .B2(n_399), .Y(n_392) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g565 ( .A(n_395), .Y(n_565) );
INVx2_ASAP7_75t_L g624 ( .A(n_395), .Y(n_624) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_396), .A2(n_494), .B(n_495), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_396), .A2(n_399), .B1(n_747), .B2(n_748), .Y(n_746) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_396), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_399), .A2(n_413), .B1(n_497), .B2(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g534 ( .A(n_399), .Y(n_534) );
BUFx3_ASAP7_75t_L g626 ( .A(n_399), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_399), .A2(n_624), .B1(n_692), .B2(n_693), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_399), .A2(n_565), .B1(n_843), .B2(n_844), .Y(n_842) );
BUFx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g475 ( .A(n_400), .Y(n_475) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_404), .Y(n_401) );
OAI222xp33_ASAP7_75t_L g845 ( .A1(n_403), .A2(n_503), .B1(n_632), .B2(n_846), .C1(n_847), .C2(n_848), .Y(n_845) );
INVx2_ASAP7_75t_L g544 ( .A(n_405), .Y(n_544) );
BUFx4f_ASAP7_75t_SL g787 ( .A(n_405), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_411), .B2(n_412), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g629 ( .A1(n_409), .A2(n_501), .B1(n_630), .B2(n_631), .C1(n_632), .C2(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_412), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_849) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx4_ASAP7_75t_L g576 ( .A(n_413), .Y(n_576) );
BUFx3_ASAP7_75t_L g701 ( .A(n_413), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_421), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g619 ( .A(n_418), .Y(n_619) );
INVx1_ASAP7_75t_L g552 ( .A(n_420), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g585 ( .A(n_429), .Y(n_585) );
BUFx2_ASAP7_75t_L g763 ( .A(n_429), .Y(n_763) );
BUFx4f_ASAP7_75t_SL g858 ( .A(n_429), .Y(n_858) );
BUFx2_ASAP7_75t_L g901 ( .A(n_429), .Y(n_901) );
INVx1_ASAP7_75t_L g597 ( .A(n_431), .Y(n_597) );
XOR2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_485), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_458), .B2(n_459), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_435), .A2(n_436), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
XOR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_457), .Y(n_436) );
NAND4xp75_ASAP7_75t_SL g437 ( .A(n_438), .B(n_439), .C(n_442), .D(n_448), .Y(n_437) );
INVx1_ASAP7_75t_L g609 ( .A(n_441), .Y(n_609) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_453), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_452), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND4xp75_ASAP7_75t_L g460 ( .A(n_461), .B(n_467), .C(n_472), .D(n_482), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
INVx2_ASAP7_75t_L g607 ( .A(n_463), .Y(n_607) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_464), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_SL g590 ( .A(n_464), .Y(n_590) );
INVx5_ASAP7_75t_SL g658 ( .A(n_464), .Y(n_658) );
INVx4_ASAP7_75t_L g767 ( .A(n_464), .Y(n_767) );
INVx2_ASAP7_75t_L g795 ( .A(n_464), .Y(n_795) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
OA211x2_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_476), .C(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g567 ( .A(n_475), .Y(n_567) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI21xp5_ASAP7_75t_SL g749 ( .A1(n_484), .A2(n_750), .B(n_751), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_524), .B2(n_525), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
XNOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_523), .Y(n_490) );
AND3x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_504), .C(n_512), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .C(n_499), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_499) );
OAI21xp5_ASAP7_75t_SL g887 ( .A1(n_501), .A2(n_888), .B(n_889), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
INVx3_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
INVx3_ASAP7_75t_L g657 ( .A(n_509), .Y(n_657) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .C(n_521), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_560), .B1(n_594), .B2(n_595), .Y(n_525) );
INVx2_ASAP7_75t_L g594 ( .A(n_526), .Y(n_594) );
XNOR2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_545), .Y(n_528) );
INVx3_ASAP7_75t_L g570 ( .A(n_530), .Y(n_570) );
OAI211xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_535), .C(n_536), .Y(n_531) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_541), .B2(n_542), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_540), .Y(n_697) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .C(n_554), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_558), .A2(n_770), .B1(n_771), .B2(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g595 ( .A(n_560), .Y(n_595) );
INVx1_ASAP7_75t_SL g592 ( .A(n_561), .Y(n_592) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_581), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_568), .C(n_573), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_567), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_883) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_571), .Y(n_568) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_570), .A2(n_695), .B(n_696), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_577), .B2(n_578), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx3_ASAP7_75t_SL g754 ( .A(n_576), .Y(n_754) );
CKINVDCx16_ASAP7_75t_R g704 ( .A(n_578), .Y(n_704) );
BUFx2_ASAP7_75t_L g756 ( .A(n_578), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_578), .A2(n_754), .B1(n_892), .B2(n_893), .Y(n_891) );
OR2x6_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND4x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .C(n_586), .D(n_589), .Y(n_581) );
BUFx2_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
INVx1_ASAP7_75t_L g824 ( .A(n_600), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_721), .B2(n_822), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_637), .B1(n_719), .B2(n_720), .Y(n_602) );
INVx1_ASAP7_75t_L g719 ( .A(n_603), .Y(n_719) );
INVx1_ASAP7_75t_L g636 ( .A(n_604), .Y(n_636) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_622), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_615), .Y(n_605) );
OAI221xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B1(n_609), .B2(n_610), .C(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_618), .B1(n_619), .B2(n_620), .C(n_621), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_629), .Y(n_622) );
OAI221xp5_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_625), .B1(n_626), .B2(n_627), .C(n_628), .Y(n_623) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx3_ASAP7_75t_L g698 ( .A(n_633), .Y(n_698) );
INVx1_ASAP7_75t_L g720 ( .A(n_637), .Y(n_720) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_665), .B2(n_718), .Y(n_638) );
INVx3_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
XOR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_664), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_642), .B(n_651), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_646), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_645), .A2(n_677), .B(n_678), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g727 ( .A1(n_645), .A2(n_728), .B(n_729), .Y(n_727) );
OAI21xp5_ASAP7_75t_SL g784 ( .A1(n_645), .A2(n_785), .B(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_659), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_662), .Y(n_801) );
INVx1_ASAP7_75t_L g718 ( .A(n_665), .Y(n_718) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B1(n_687), .B2(n_688), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
XOR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_686), .Y(n_668) );
NAND4xp75_ASAP7_75t_SL g669 ( .A(n_670), .B(n_679), .C(n_684), .D(n_685), .Y(n_669) );
NOR2xp67_ASAP7_75t_SL g670 ( .A(n_671), .B(n_676), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .C(n_675), .Y(n_671) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_SL g716 ( .A(n_689), .Y(n_716) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_690), .B(n_705), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .C(n_699), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_699) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g852 ( .A(n_704), .Y(n_852) );
AND4x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .C(n_711), .D(n_713), .Y(n_705) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g822 ( .A(n_721), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_778), .B2(n_821), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AO22x2_ASAP7_75t_SL g723 ( .A1(n_724), .A2(n_743), .B1(n_776), .B2(n_777), .Y(n_723) );
INVx4_ASAP7_75t_SL g776 ( .A(n_724), .Y(n_776) );
AO22x2_ASAP7_75t_L g805 ( .A1(n_724), .A2(n_776), .B1(n_806), .B2(n_807), .Y(n_805) );
XOR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_742), .Y(n_724) );
NAND3x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_736), .C(n_739), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .C(n_734), .Y(n_730) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g777 ( .A(n_743), .Y(n_777) );
INVx1_ASAP7_75t_L g774 ( .A(n_744), .Y(n_774) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_758), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .C(n_753), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_754), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_764), .C(n_769), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g821 ( .A(n_778), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B1(n_804), .B2(n_805), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_SL g802 ( .A(n_782), .Y(n_802) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_792), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_788), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_789), .B(n_791), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_798), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g864 ( .A(n_797), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
XOR2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_820), .Y(n_807) );
NAND4xp75_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .C(n_816), .D(n_819), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
AND2x2_ASAP7_75t_SL g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx1_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_831), .Y(n_826) );
OR2x2_ASAP7_75t_SL g905 ( .A(n_827), .B(n_832), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_828), .Y(n_868) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_829), .B(n_872), .Y(n_875) );
CKINVDCx16_ASAP7_75t_R g872 ( .A(n_830), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
OAI322xp33_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_867), .A3(n_869), .B1(n_873), .B2(n_876), .C1(n_877), .C2(n_903), .Y(n_838) );
INVx1_ASAP7_75t_L g866 ( .A(n_840), .Y(n_866) );
AND2x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_853), .Y(n_840) );
NOR3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_845), .C(n_849), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_859), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_857), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g859 ( .A(n_860), .B(n_862), .Y(n_859) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g902 ( .A(n_881), .Y(n_902) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_894), .Y(n_881) );
NOR3xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_887), .C(n_891), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_898), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_904), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_905), .Y(n_904) );
endmodule