module fake_jpeg_9815_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_48),
.B1(n_26),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_34),
.B1(n_25),
.B2(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_25),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_60),
.Y(n_73)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_57),
.Y(n_76)
);

CKINVDCx12_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_21),
.B(n_17),
.C(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_32),
.B1(n_36),
.B2(n_24),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_69),
.B1(n_72),
.B2(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_26),
.B1(n_25),
.B2(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_34),
.B1(n_62),
.B2(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_68),
.B1(n_70),
.B2(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_89),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_51),
.C(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_47),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_37),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_99),
.B(n_19),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_39),
.B1(n_61),
.B2(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_40),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_102),
.C(n_27),
.D(n_20),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_38),
.B(n_20),
.C(n_50),
.D(n_31),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_80),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_116),
.C(n_93),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_95),
.B1(n_90),
.B2(n_85),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_107),
.B1(n_119),
.B2(n_120),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_54),
.B1(n_61),
.B2(n_40),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_117),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_22),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_39),
.C(n_80),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_92),
.B(n_83),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_15),
.B1(n_33),
.B2(n_38),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_15),
.B1(n_33),
.B2(n_38),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_131),
.B(n_110),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_92),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_125),
.C(n_22),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_135),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_99),
.B(n_101),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_134),
.B(n_65),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_91),
.C(n_102),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_27),
.C(n_65),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_33),
.B1(n_31),
.B2(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_100),
.B1(n_84),
.B2(n_21),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_110),
.B1(n_103),
.B2(n_16),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_141),
.C(n_146),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_153),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_109),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_154),
.C(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_84),
.B1(n_17),
.B2(n_19),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_151),
.B1(n_139),
.B2(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_27),
.B1(n_20),
.B2(n_65),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_122),
.C(n_132),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_156),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_165),
.B(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_151),
.B1(n_160),
.B2(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_142),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_134),
.B(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_1),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_156),
.C(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_126),
.C(n_7),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_7),
.C(n_12),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_8),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_0),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_172),
.B(n_173),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_183),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_170),
.B(n_177),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_180),
.B(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_190),
.B(n_8),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_195),
.B(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_177),
.B(n_11),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_13),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_200),
.B1(n_197),
.B2(n_1),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_3),
.Y(n_202)
);


endmodule