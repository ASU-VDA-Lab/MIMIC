module fake_jpeg_23694_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_27),
.B(n_28),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_47),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_16),
.B1(n_26),
.B2(n_25),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_56),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_36),
.B1(n_22),
.B2(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_58),
.B1(n_61),
.B2(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_33),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_35),
.B1(n_47),
.B2(n_45),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_13),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_52),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_39),
.C(n_38),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_83),
.C(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_31),
.B(n_16),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_25),
.B(n_23),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_39),
.C(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_39),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_61),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_93),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_99),
.C(n_86),
.Y(n_110)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_56),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_66),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_24),
.B(n_23),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_66),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_19),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_60),
.C(n_58),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_73),
.B1(n_70),
.B2(n_78),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_103),
.B1(n_98),
.B2(n_24),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_82),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_108),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_112),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_107),
.C(n_90),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_81),
.B1(n_76),
.B2(n_24),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_93),
.B1(n_97),
.B2(n_87),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_88),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.C(n_23),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_95),
.C(n_89),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_102),
.B1(n_104),
.B2(n_96),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_128),
.B1(n_125),
.B2(n_121),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_125),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_107),
.B(n_117),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_19),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_137),
.B1(n_135),
.B2(n_132),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_141),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_21),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_17),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

OAI322xp33_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_131),
.A3(n_127),
.B1(n_119),
.B2(n_123),
.C1(n_21),
.C2(n_20),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_20),
.B1(n_17),
.B2(n_13),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_20),
.B1(n_17),
.B2(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_1),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_139),
.C(n_142),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_2),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_155),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_146),
.B(n_151),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_150),
.B(n_1),
.Y(n_159)
);

AOI31xp67_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_148),
.A3(n_147),
.B(n_4),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_7),
.B(n_9),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_5),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_152),
.B(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_10),
.C(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_164),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_163),
.B(n_11),
.Y(n_172)
);

NOR4xp25_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_172),
.C(n_167),
.D(n_11),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.C(n_168),
.Y(n_174)
);

OAI311xp33_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_175),
.A3(n_10),
.B1(n_12),
.C1(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_12),
.Y(n_177)
);


endmodule