module real_aes_6642_n_5 (n_4, n_0, n_3, n_2, n_1, n_5);
input n_4;
input n_0;
input n_3;
input n_2;
input n_1;
output n_5;
wire n_16;
wire n_13;
wire n_15;
wire n_7;
wire n_9;
wire n_6;
wire n_12;
wire n_8;
wire n_14;
wire n_10;
wire n_11;
AOI22xp5_ASAP7_75t_SL g5 ( .A1(n_0), .A2(n_6), .B1(n_14), .B2(n_16), .Y(n_5) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
CKINVDCx14_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_1), .B(n_9), .Y(n_13) );
OAI21xp5_ASAP7_75t_L g6 ( .A1(n_2), .A2(n_3), .B(n_7), .Y(n_6) );
NAND3xp33_ASAP7_75t_SL g15 ( .A(n_2), .B(n_4), .C(n_12), .Y(n_15) );
INVx1_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
AOI21xp5_ASAP7_75t_L g10 ( .A1(n_3), .A2(n_11), .B(n_12), .Y(n_10) );
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
AOI21xp5_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_9), .B(n_10), .Y(n_7) );
INVx1_ASAP7_75t_SL g12 ( .A(n_13), .Y(n_12) );
INVx1_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
endmodule