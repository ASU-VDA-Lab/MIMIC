module fake_jpeg_17896_n_235 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_47),
.Y(n_71)
);

NOR2x1_ASAP7_75t_R g47 ( 
.A(n_35),
.B(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_29),
.B1(n_18),
.B2(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_24),
.B1(n_14),
.B2(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_31),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_37),
.B(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_68),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_32),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_57),
.B1(n_55),
.B2(n_34),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_32),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_58),
.B(n_22),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_76),
.Y(n_84)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22x1_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_58),
.B1(n_30),
.B2(n_17),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_98),
.B(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_44),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_69),
.B(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_49),
.B1(n_42),
.B2(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_97),
.B1(n_48),
.B2(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_42),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_0),
.Y(n_98)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_73),
.B(n_71),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_105),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_117),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_75),
.B1(n_60),
.B2(n_61),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_93),
.B1(n_87),
.B2(n_91),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_71),
.C(n_52),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_112),
.C(n_115),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_52),
.C(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_36),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_120),
.B1(n_34),
.B2(n_40),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_52),
.C(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_69),
.B1(n_66),
.B2(n_48),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_66),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_111),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_86),
.B1(n_97),
.B2(n_92),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_92),
.B1(n_98),
.B2(n_95),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_98),
.B1(n_80),
.B2(n_81),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_129),
.B(n_140),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_121),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_80),
.B1(n_55),
.B2(n_69),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_129),
.B1(n_103),
.B2(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_99),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_132),
.B1(n_140),
.B2(n_131),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_76),
.B(n_1),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_112),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_147),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_125),
.B1(n_126),
.B2(n_141),
.C(n_122),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_104),
.B(n_117),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_0),
.B(n_1),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_153),
.B(n_157),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_106),
.C(n_105),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_152),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_105),
.B(n_107),
.C(n_106),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_28),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_109),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_101),
.B2(n_40),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_103),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_99),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_175),
.B1(n_150),
.B2(n_147),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_139),
.B1(n_133),
.B2(n_116),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_170),
.B1(n_157),
.B2(n_153),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_76),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_100),
.B1(n_99),
.B2(n_63),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_156),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_177),
.C(n_160),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_100),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_149),
.B1(n_155),
.B2(n_158),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_192),
.B1(n_170),
.B2(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_186),
.C(n_190),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_188),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_171),
.B1(n_176),
.B2(n_174),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_150),
.C(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_151),
.B(n_11),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_11),
.B(n_12),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_63),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_28),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_21),
.C(n_33),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_165),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_21),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_173),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_10),
.B(n_13),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_16),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_197),
.C(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_8),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_185),
.B(n_183),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_197),
.B1(n_195),
.B2(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_183),
.C(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_213),
.B1(n_7),
.B2(n_13),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_36),
.C(n_7),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_21),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_202),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_221),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_3),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_0),
.C(n_1),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_211),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_226),
.B(n_225),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_214),
.B(n_5),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

AOI31xp33_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_220),
.A3(n_221),
.B(n_216),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_4),
.B(n_6),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_230),
.B1(n_9),
.B2(n_10),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_231),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_12),
.Y(n_235)
);


endmodule