module fake_jpeg_881_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_80),
.Y(n_90)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_0),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

OR2x6_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_1),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_64),
.B1(n_70),
.B2(n_57),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_59),
.B1(n_56),
.B2(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_92),
.B1(n_64),
.B2(n_67),
.Y(n_102)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_59),
.B1(n_71),
.B2(n_65),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_57),
.B(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_99),
.C(n_54),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_88),
.B1(n_51),
.B2(n_61),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_50),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_68),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_70),
.B1(n_58),
.B2(n_69),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_72),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_69),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_68),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_55),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_127),
.Y(n_148)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_94),
.B1(n_51),
.B2(n_60),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_135),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_5),
.Y(n_152)
);

NAND2x1_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_130),
.B(n_8),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_72),
.B(n_4),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_61),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_108),
.B1(n_98),
.B2(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_2),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_2),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_103),
.C(n_27),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_145),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_4),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_130),
.B(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_160),
.B(n_159),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_28),
.C(n_47),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_26),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_38),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_48),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_161),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_16),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_8),
.B(n_9),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_30),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_163),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_169),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_172),
.B1(n_178),
.B2(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_15),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_180),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_138),
.B(n_149),
.C(n_160),
.D(n_147),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_191),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_139),
.C(n_158),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_173),
.C(n_166),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_174),
.B(n_168),
.C(n_170),
.D(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_199),
.C(n_157),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_197),
.A2(n_192),
.B1(n_185),
.B2(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_179),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_164),
.C(n_166),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_191),
.B(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_190),
.B1(n_144),
.B2(n_20),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_196),
.B1(n_199),
.B2(n_194),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_207),
.A2(n_208),
.B1(n_202),
.B2(n_31),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_210),
.B(n_36),
.C(n_40),
.D(n_41),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_206),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_207),
.B(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);


endmodule