module fake_jpeg_8948_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_45),
.B(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_32),
.B1(n_18),
.B2(n_17),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_64),
.B1(n_38),
.B2(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_54),
.Y(n_78)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_55),
.B1(n_19),
.B2(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_32),
.B1(n_18),
.B2(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_26),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_69),
.Y(n_83)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_26),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_25),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_38),
.B1(n_22),
.B2(n_20),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_87),
.B1(n_88),
.B2(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_89),
.B1(n_61),
.B2(n_27),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_39),
.B(n_26),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_20),
.B1(n_22),
.B2(n_34),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_20),
.B1(n_22),
.B2(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_78),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_36),
.B1(n_23),
.B2(n_27),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_27),
.B1(n_25),
.B2(n_28),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_53),
.B(n_47),
.C(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_104),
.B1(n_113),
.B2(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_107),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_39),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_115),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_111),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_61),
.B1(n_59),
.B2(n_50),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_68),
.B1(n_63),
.B2(n_48),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_86),
.B1(n_57),
.B2(n_62),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_97),
.B1(n_118),
.B2(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_36),
.B1(n_60),
.B2(n_63),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_60),
.A3(n_42),
.B1(n_44),
.B2(n_36),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_106),
.B(n_102),
.C(n_107),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_0),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_76),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_52),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_119),
.B1(n_98),
.B2(n_97),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_76),
.B1(n_92),
.B2(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_137),
.B1(n_152),
.B2(n_125),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_104),
.B(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_137),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_90),
.B1(n_86),
.B2(n_73),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_142),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_73),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_30),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_75),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_147),
.B(n_150),
.C(n_33),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_90),
.B1(n_51),
.B2(n_92),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_44),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_44),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_33),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_30),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_30),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_157),
.B(n_171),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_99),
.B(n_100),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_124),
.B1(n_131),
.B2(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_178),
.B1(n_133),
.B2(n_136),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_163),
.B(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_170),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_33),
.B1(n_31),
.B2(n_24),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_174),
.B(n_147),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_163),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_131),
.B1(n_130),
.B2(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_140),
.C(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_193),
.C(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_199),
.B1(n_207),
.B2(n_156),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_145),
.C(n_127),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_133),
.B1(n_142),
.B2(n_143),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_136),
.C(n_143),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_31),
.B1(n_147),
.B2(n_77),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_205),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_77),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_204),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_72),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_9),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_168),
.B(n_154),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_173),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_180),
.B1(n_179),
.B2(n_175),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_95),
.B(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

BUFx12_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_225),
.Y(n_246)
);

XNOR2x2_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_164),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_218),
.B(n_189),
.Y(n_240)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_223),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_153),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_175),
.B1(n_177),
.B2(n_176),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_229),
.B1(n_196),
.B2(n_197),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_230),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_190),
.A2(n_156),
.B1(n_162),
.B2(n_157),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_1),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_186),
.C(n_203),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_235),
.C(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_193),
.C(n_204),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_190),
.B(n_192),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_244),
.B(n_229),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_226),
.B1(n_232),
.B2(n_218),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_202),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_95),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_253),
.C(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_220),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_95),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_240),
.B1(n_251),
.B2(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_219),
.B(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_259),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_221),
.B1(n_214),
.B2(n_10),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_236),
.B(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_8),
.B(n_15),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_239),
.C(n_249),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_10),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_246),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.C(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_235),
.C(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_2),
.C(n_3),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_244),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_262),
.C(n_254),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_273),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_277),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_247),
.C(n_252),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_251),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_265),
.C(n_268),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_265),
.C(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_290),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_270),
.A3(n_287),
.B1(n_277),
.B2(n_283),
.C1(n_272),
.C2(n_291),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_234),
.C(n_269),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_261),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_250),
.C(n_5),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_270),
.B(n_275),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_14),
.B(n_15),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_11),
.A3(n_6),
.B1(n_7),
.B2(n_10),
.C1(n_16),
.C2(n_13),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_13),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_286),
.B(n_6),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_307),
.B(n_296),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_14),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_295),
.B(n_297),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_302),
.C(n_308),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_310),
.B1(n_305),
.B2(n_4),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_4),
.B1(n_310),
.B2(n_305),
.Y(n_314)
);


endmodule