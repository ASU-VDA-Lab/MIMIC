module fake_jpeg_6281_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_35),
.A2(n_39),
.B(n_45),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_19),
.B1(n_33),
.B2(n_32),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_2),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_49),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_3),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_20),
.B(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_5),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_27),
.B1(n_22),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_52),
.A2(n_73),
.B1(n_93),
.B2(n_97),
.Y(n_126)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_58),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_56),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_57),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_64),
.Y(n_105)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_70),
.Y(n_109)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_27),
.B1(n_28),
.B2(n_22),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_89),
.B(n_7),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_94),
.Y(n_108)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_90),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_45),
.B(n_6),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_42),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_16),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_30),
.B1(n_21),
.B2(n_25),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_21),
.B(n_34),
.C(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_89),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_25),
.B(n_34),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_25),
.C(n_16),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_120),
.Y(n_129)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_16),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_97),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_16),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_60),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_73),
.B1(n_104),
.B2(n_123),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_93),
.B1(n_52),
.B2(n_84),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_55),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_139),
.B(n_100),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_88),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_8),
.B(n_11),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_70),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_60),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_59),
.B1(n_86),
.B2(n_82),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_54),
.B1(n_59),
.B2(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_156),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_114),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_147),
.B1(n_148),
.B2(n_155),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_53),
.B1(n_18),
.B2(n_23),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_112),
.B1(n_110),
.B2(n_100),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_29),
.A3(n_23),
.B1(n_18),
.B2(n_10),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_157),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_66),
.B1(n_18),
.B2(n_29),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_29),
.B1(n_23),
.B2(n_65),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_99),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_7),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_8),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_120),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_109),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_74),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_74),
.B1(n_9),
.B2(n_11),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_8),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_12),
.CI(n_13),
.CON(n_178),
.SN(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_168),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_163),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_115),
.B(n_113),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_166),
.A2(n_175),
.B(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_103),
.C(n_113),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_169),
.C(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_117),
.C(n_99),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_176),
.Y(n_189)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_13),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_14),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_14),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_158),
.B(n_134),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_127),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_192),
.Y(n_214)
);

XOR2x2_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_134),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_143),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_195),
.C(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_140),
.C(n_129),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_181),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_145),
.B1(n_137),
.B2(n_139),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_139),
.B1(n_148),
.B2(n_153),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_183),
.Y(n_206)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_159),
.B(n_175),
.C(n_186),
.D(n_176),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_155),
.C(n_146),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_162),
.C(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_191),
.A3(n_165),
.B1(n_204),
.B2(n_193),
.C1(n_199),
.C2(n_188),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_195),
.Y(n_231)
);

NAND2x1_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_166),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_209),
.B(n_210),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_171),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_220),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_168),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_221),
.B(n_196),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_219),
.C(n_194),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_179),
.B1(n_163),
.B2(n_161),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_170),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_162),
.C(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

XOR2x1_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_187),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_227),
.B(n_229),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_189),
.B1(n_219),
.B2(n_146),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_232),
.C(n_214),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_213),
.B1(n_217),
.B2(n_211),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_212),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_212),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_221),
.B(n_189),
.C(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_213),
.B1(n_210),
.B2(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_201),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_237),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_232),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_223),
.B(n_228),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_226),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_190),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_243),
.Y(n_251)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_239),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_247),
.B(n_230),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_174),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_249),
.B(n_250),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_233),
.B1(n_230),
.B2(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_174),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_231),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_245),
.B(n_236),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_249),
.C(n_185),
.Y(n_258)
);

OAI221xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_255),
.B1(n_258),
.B2(n_164),
.C(n_172),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_178),
.Y(n_261)
);


endmodule