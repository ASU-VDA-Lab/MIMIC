module fake_aes_3380_n_546 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_546);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_546;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g78 ( .A(n_75), .Y(n_78) );
INVx3_ASAP7_75t_L g79 ( .A(n_39), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_58), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_17), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_61), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_6), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_0), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_31), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_6), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_32), .Y(n_87) );
OR2x2_ASAP7_75t_L g88 ( .A(n_48), .B(n_14), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_25), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_21), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_24), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_67), .Y(n_92) );
OR2x2_ASAP7_75t_L g93 ( .A(n_22), .B(n_36), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_66), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_50), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_40), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_73), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_68), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_15), .Y(n_101) );
NOR2xp67_ASAP7_75t_L g102 ( .A(n_34), .B(n_41), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_64), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_43), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_42), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_18), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_77), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_45), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_55), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_3), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_11), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_112), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_83), .B(n_0), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_84), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_95), .B(n_1), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_112), .Y(n_121) );
AND2x6_ASAP7_75t_L g122 ( .A(n_79), .B(n_37), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_107), .B(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_79), .Y(n_126) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_85), .A2(n_38), .B(n_74), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_113), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_128) );
INVx2_ASAP7_75t_SL g129 ( .A(n_78), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_86), .B(n_114), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_86), .B(n_4), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_101), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_101), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_88), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_119), .B(n_100), .Y(n_139) );
INVx4_ASAP7_75t_SL g140 ( .A(n_122), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_130), .B(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_126), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_117), .A2(n_87), .B1(n_110), .B2(n_109), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_119), .B(n_82), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_124), .B(n_90), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_124), .B(n_90), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_122), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_125), .B(n_111), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_122), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_125), .B(n_110), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_129), .B(n_99), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_116), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_122), .A2(n_101), .B1(n_104), .B2(n_96), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_117), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_134), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_123), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_129), .B(n_109), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_141), .A2(n_122), .B1(n_123), .B2(n_133), .Y(n_164) );
NOR2xp33_ASAP7_75t_SL g165 ( .A(n_141), .B(n_91), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_141), .A2(n_133), .B1(n_132), .B2(n_120), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_146), .B(n_133), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_145), .B(n_131), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
OR2x6_ASAP7_75t_L g172 ( .A(n_141), .B(n_128), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_151), .A2(n_132), .B1(n_137), .B2(n_136), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_127), .B(n_121), .C(n_115), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_148), .B(n_103), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_139), .B(n_103), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_140), .B(n_115), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_127), .B(n_121), .C(n_97), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_163), .B(n_91), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_152), .B(n_92), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_142), .B(n_92), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_151), .B(n_94), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_153), .B(n_94), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_161), .B(n_106), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
AO22x1_ASAP7_75t_L g195 ( .A1(n_151), .A2(n_118), .B1(n_106), .B2(n_98), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_159), .A2(n_101), .B1(n_105), .B2(n_108), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_166), .B(n_159), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_172), .B(n_128), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_173), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_172), .A2(n_157), .B1(n_144), .B2(n_156), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_192), .A2(n_159), .B(n_140), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_192), .A2(n_159), .B(n_140), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_166), .B(n_144), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_182), .B(n_93), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_164), .A2(n_102), .B1(n_140), .B2(n_135), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_173), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_170), .B(n_8), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_173), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_174), .Y(n_211) );
NOR2xp33_ASAP7_75t_R g212 ( .A(n_165), .B(n_9), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_181), .B(n_9), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_193), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_174), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_175), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_169), .A2(n_162), .B(n_160), .C(n_147), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_165), .B(n_135), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_171), .B(n_135), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_175), .A2(n_135), .B1(n_134), .B2(n_147), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_171), .B(n_135), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_194), .B(n_134), .Y(n_226) );
NOR2xp67_ASAP7_75t_L g227 ( .A(n_189), .B(n_10), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_172), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_181), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_209), .A2(n_172), .B(n_178), .C(n_180), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_229), .B(n_195), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_202), .A2(n_192), .B(n_184), .Y(n_232) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_220), .A2(n_185), .B(n_186), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_208), .B(n_183), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_200), .A2(n_172), .B1(n_177), .B2(n_185), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_203), .A2(n_190), .B(n_187), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_214), .A2(n_191), .B(n_188), .C(n_186), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_208), .Y(n_238) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_220), .A2(n_179), .B(n_176), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_204), .B(n_195), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_219), .A2(n_183), .B(n_176), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_207), .A2(n_179), .B(n_167), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_198), .A2(n_196), .B(n_182), .C(n_194), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_210), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_212), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_228), .A2(n_182), .B1(n_194), .B2(n_168), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_198), .A2(n_182), .B1(n_168), .B2(n_162), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_198), .A2(n_168), .B1(n_160), .B2(n_12), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_204), .B(n_168), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_217), .A2(n_221), .B(n_225), .C(n_226), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_221), .B(n_168), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_216), .A2(n_168), .B1(n_11), .B2(n_13), .Y(n_255) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_225), .A2(n_10), .A3(n_13), .B(n_14), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_231), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_234), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_230), .A2(n_222), .B(n_226), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_224), .B(n_222), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_243), .A2(n_227), .B(n_199), .C(n_215), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
OAI21xp33_ASAP7_75t_SL g264 ( .A1(n_233), .A2(n_201), .B(n_205), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_238), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_247), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_246), .B(n_212), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_244), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_232), .A2(n_224), .B(n_199), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_245), .B(n_215), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_241), .A2(n_201), .B(n_223), .Y(n_275) );
OAI221xp5_ASAP7_75t_L g276 ( .A1(n_235), .A2(n_206), .B1(n_197), .B2(n_213), .C(n_15), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_240), .A2(n_213), .B(n_206), .C(n_197), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_246), .A2(n_213), .B1(n_16), .B2(n_20), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_256), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_274), .A2(n_241), .B(n_233), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_270), .B(n_256), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_270), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_268), .Y(n_287) );
AOI21xp5_ASAP7_75t_SL g288 ( .A1(n_277), .A2(n_251), .B(n_255), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_266), .B(n_242), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_268), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_276), .A2(n_242), .B(n_236), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_262), .A2(n_250), .B(n_254), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_258), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_271), .B(n_249), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_261), .A2(n_254), .B(n_248), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_267), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_258), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_257), .B(n_16), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_258), .A2(n_239), .B1(n_213), .B2(n_256), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_269), .B(n_253), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_300), .B(n_279), .C(n_274), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_298), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_296), .B(n_279), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_280), .B(n_267), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_256), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_284), .B(n_263), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_290), .B(n_271), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_282), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_280), .B(n_259), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_296), .B(n_259), .Y(n_315) );
NOR2x1_ASAP7_75t_SL g316 ( .A(n_283), .B(n_278), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_293), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_287), .B(n_273), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_283), .B(n_273), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_285), .B(n_264), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_293), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_290), .B(n_264), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_285), .B(n_275), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_286), .B(n_275), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_299), .A2(n_278), .B1(n_260), .B2(n_275), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_286), .B(n_275), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_282), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_281), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_281), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_308), .B(n_281), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_308), .B(n_297), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_312), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_308), .B(n_289), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_310), .B(n_289), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_310), .B(n_289), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_310), .B(n_289), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_330), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_320), .B(n_289), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_305), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_306), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_320), .B(n_281), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_304), .B(n_294), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_323), .B(n_291), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_305), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_323), .B(n_295), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_306), .B(n_301), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_304), .B(n_288), .Y(n_350) );
NOR2x1p5_ASAP7_75t_L g351 ( .A(n_327), .B(n_288), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_309), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_324), .B(n_239), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_324), .B(n_292), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_326), .B(n_292), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_326), .B(n_239), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_272), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_330), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_328), .B(n_19), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_322), .B(n_26), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_311), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_319), .B(n_27), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_311), .B(n_28), .Y(n_366) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_314), .B(n_29), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_303), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_319), .B(n_30), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_327), .B(n_35), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
NOR2x1_ASAP7_75t_L g372 ( .A(n_303), .B(n_44), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_307), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_332), .B(n_331), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_344), .B(n_330), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_357), .B(n_318), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_332), .B(n_321), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_332), .B(n_321), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_344), .B(n_327), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_357), .B(n_307), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_341), .B(n_317), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_364), .B(n_302), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_375), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_333), .B(n_318), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_341), .B(n_317), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_340), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_340), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_364), .B(n_302), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_375), .B(n_313), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_367), .A2(n_325), .B(n_313), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_346), .B(n_314), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_334), .Y(n_394) );
AOI22x1_ASAP7_75t_L g395 ( .A1(n_351), .A2(n_315), .B1(n_316), .B2(n_325), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_368), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_346), .B(n_316), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_356), .A2(n_315), .B1(n_47), .B2(n_49), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_346), .B(n_46), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_348), .B(n_51), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_348), .B(n_53), .Y(n_402) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_372), .B(n_54), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_348), .B(n_56), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_356), .B(n_358), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_334), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_358), .B(n_57), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_343), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_367), .A2(n_59), .B1(n_60), .B2(n_62), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_335), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_340), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_340), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_345), .B(n_63), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_374), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_343), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g416 ( .A1(n_367), .A2(n_65), .B(n_69), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_333), .B(n_71), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_335), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_353), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_361), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_345), .B(n_72), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_361), .Y(n_424) );
NOR2x1p5_ASAP7_75t_L g425 ( .A(n_350), .B(n_337), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_371), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_383), .B(n_336), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_426), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_376), .B(n_373), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_419), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_422), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_376), .B(n_373), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_392), .A2(n_350), .B1(n_337), .B2(n_372), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_425), .B(n_336), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_414), .B(n_349), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_425), .B(n_338), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_422), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_418), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_405), .B(n_349), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g442 ( .A1(n_392), .A2(n_366), .B(n_361), .C(n_355), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_405), .B(n_355), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_416), .B(n_363), .C(n_366), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_408), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_386), .B(n_338), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_417), .A2(n_351), .B1(n_339), .B2(n_369), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_383), .B(n_339), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_386), .B(n_354), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_403), .B(n_370), .Y(n_451) );
CKINVDCx14_ASAP7_75t_R g452 ( .A(n_387), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_415), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_387), .B(n_354), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_394), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_384), .B(n_354), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_382), .B(n_359), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_398), .A2(n_369), .B1(n_365), .B2(n_363), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_384), .B(n_361), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_393), .B(n_359), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_393), .B(n_359), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_379), .B(n_359), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_379), .B(n_360), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_382), .B(n_378), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_378), .B(n_342), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_390), .B(n_342), .Y(n_468) );
AOI211xp5_ASAP7_75t_L g469 ( .A1(n_416), .A2(n_398), .B(n_423), .C(n_413), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_390), .B(n_342), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_391), .B(n_360), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_466), .B(n_397), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_457), .B(n_385), .Y(n_474) );
NOR4xp25_ASAP7_75t_L g475 ( .A(n_442), .B(n_396), .C(n_407), .D(n_410), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_452), .B(n_396), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_460), .A2(n_395), .B1(n_381), .B2(n_417), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_467), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_448), .A2(n_395), .B1(n_381), .B2(n_402), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_435), .B(n_381), .Y(n_483) );
OAI21xp5_ASAP7_75t_SL g484 ( .A1(n_448), .A2(n_409), .B(n_403), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_469), .A2(n_391), .B1(n_406), .B2(n_407), .C(n_399), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_433), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_440), .B(n_377), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_440), .B(n_381), .Y(n_489) );
NAND2xp33_ASAP7_75t_SL g490 ( .A(n_435), .B(n_401), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_439), .B(n_377), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_429), .Y(n_492) );
OAI31xp33_ASAP7_75t_L g493 ( .A1(n_434), .A2(n_401), .A3(n_402), .B(n_404), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_457), .B(n_377), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_443), .B(n_377), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_443), .A2(n_380), .B1(n_394), .B2(n_406), .C(n_410), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
AOI211x1_ASAP7_75t_L g500 ( .A1(n_432), .A2(n_404), .B(n_400), .C(n_380), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_454), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_437), .B(n_385), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_488), .Y(n_503) );
AOI211xp5_ASAP7_75t_SL g504 ( .A1(n_478), .A2(n_445), .B(n_400), .C(n_453), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_480), .B(n_438), .Y(n_505) );
AOI21xp33_ASAP7_75t_SL g506 ( .A1(n_478), .A2(n_451), .B(n_453), .Y(n_506) );
AOI221x1_ASAP7_75t_L g507 ( .A1(n_476), .A2(n_431), .B1(n_444), .B2(n_461), .C(n_468), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_479), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_481), .B(n_461), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_490), .A2(n_437), .B(n_447), .C(n_450), .Y(n_510) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_492), .A2(n_470), .B(n_468), .C(n_472), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_482), .A2(n_451), .B1(n_470), .B2(n_458), .C(n_406), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g513 ( .A1(n_484), .A2(n_365), .B(n_463), .C(n_462), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_485), .A2(n_465), .B1(n_464), .B2(n_471), .Y(n_514) );
OAI21xp33_ASAP7_75t_L g515 ( .A1(n_475), .A2(n_428), .B(n_449), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_494), .A2(n_370), .B(n_459), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_493), .A2(n_415), .B(n_420), .C(n_370), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_489), .A2(n_455), .B(n_370), .C(n_420), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_497), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_486), .B(n_389), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_504), .A2(n_498), .B1(n_473), .B2(n_477), .C(n_474), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_506), .A2(n_500), .B1(n_487), .B2(n_474), .C(n_491), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_514), .B(n_501), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_512), .B(n_499), .C(n_496), .Y(n_524) );
AOI21xp33_ASAP7_75t_SL g525 ( .A1(n_517), .A2(n_502), .B(n_483), .Y(n_525) );
NOR2x1_ASAP7_75t_L g526 ( .A(n_510), .B(n_502), .Y(n_526) );
NOR2xp33_ASAP7_75t_SL g527 ( .A(n_508), .B(n_495), .Y(n_527) );
NOR2xp33_ASAP7_75t_R g528 ( .A(n_514), .B(n_76), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g529 ( .A1(n_515), .A2(n_389), .B1(n_421), .B2(n_412), .C1(n_388), .C2(n_424), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_513), .A2(n_389), .B1(n_421), .B2(n_412), .C(n_388), .Y(n_530) );
OAI211xp5_ASAP7_75t_SL g531 ( .A1(n_529), .A2(n_511), .B(n_518), .C(n_516), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_521), .A2(n_511), .B1(n_503), .B2(n_519), .C(n_505), .Y(n_532) );
NOR3xp33_ASAP7_75t_L g533 ( .A(n_525), .B(n_509), .C(n_520), .Y(n_533) );
OR5x1_ASAP7_75t_L g534 ( .A(n_526), .B(n_507), .C(n_411), .D(n_388), .E(n_412), .Y(n_534) );
NOR2xp67_ASAP7_75t_L g535 ( .A(n_523), .B(n_411), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_534), .Y(n_536) );
AND3x2_ASAP7_75t_L g537 ( .A(n_532), .B(n_527), .C(n_524), .Y(n_537) );
NAND4xp75_ASAP7_75t_L g538 ( .A(n_535), .B(n_522), .C(n_530), .D(n_528), .Y(n_538) );
NOR3xp33_ASAP7_75t_SL g539 ( .A(n_538), .B(n_531), .C(n_533), .Y(n_539) );
NAND3xp33_ASAP7_75t_SL g540 ( .A(n_536), .B(n_362), .C(n_411), .Y(n_540) );
OAI22x1_ASAP7_75t_L g541 ( .A1(n_539), .A2(n_537), .B1(n_362), .B2(n_421), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_541), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_542), .A2(n_540), .B(n_424), .Y(n_543) );
AOI21xp5_ASAP7_75t_SL g544 ( .A1(n_543), .A2(n_424), .B(n_347), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_544), .A2(n_347), .B(n_352), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_545), .A2(n_347), .B1(n_352), .B2(n_540), .Y(n_546) );
endmodule