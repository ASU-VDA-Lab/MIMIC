module fake_jpeg_444_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_18),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_82),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_54),
.B1(n_55),
.B2(n_52),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_54),
.B1(n_55),
.B2(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_62),
.Y(n_102)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_80),
.B1(n_50),
.B2(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_64),
.B(n_63),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_57),
.B(n_58),
.Y(n_118)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_0),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_52),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_111),
.B1(n_57),
.B2(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_50),
.B1(n_77),
.B2(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_21),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_3),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_139),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_3),
.B(n_4),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_15),
.B(n_16),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_22),
.C(n_44),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_135),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_8),
.B(n_9),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_39),
.Y(n_157)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_29),
.B1(n_41),
.B2(n_40),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_19),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_146),
.C(n_122),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_10),
.B(n_11),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_14),
.Y(n_151)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_32),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_153),
.B(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_17),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_24),
.C(n_33),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_37),
.C(n_38),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_169),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_129),
.B1(n_135),
.B2(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_128),
.B1(n_137),
.B2(n_132),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_173),
.B(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_162),
.B1(n_161),
.B2(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_179),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_152),
.B(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_178),
.B(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_174),
.B(n_175),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_182),
.B(n_164),
.Y(n_184)
);

OAI31xp33_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_147),
.A3(n_149),
.B(n_166),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_166),
.Y(n_186)
);


endmodule