module fake_netlist_5_1365_n_188 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_188);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_188;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_122;
wire n_82;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_136;
wire n_146;
wire n_86;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_123;
wire n_38;
wire n_113;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_64;
wire n_106;
wire n_102;
wire n_77;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_141;
wire n_97;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_8),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

OAI22x1_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_0),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_46),
.C(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_4),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_40),
.C(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_57),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_48),
.B1(n_45),
.B2(n_32),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_24),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR4xp25_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_71),
.C(n_61),
.D(n_62),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_85),
.B(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_83),
.Y(n_94)
);

NAND3x1_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_71),
.C(n_68),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_56),
.Y(n_96)
);

AO31x2_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_55),
.A3(n_68),
.B(n_62),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_66),
.B(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_72),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_54),
.B(n_60),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_66),
.C(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

OR2x6_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_80),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_75),
.B(n_87),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_79),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_87),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_76),
.B(n_84),
.Y(n_111)
);

OAI221xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_80),
.B1(n_92),
.B2(n_98),
.C(n_102),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_93),
.B(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_110),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_102),
.B1(n_98),
.B2(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_95),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_106),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_105),
.B1(n_106),
.B2(n_110),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_112),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_82),
.C(n_74),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_116),
.Y(n_140)
);

OAI322xp33_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_82),
.A3(n_67),
.B1(n_65),
.B2(n_96),
.C1(n_63),
.C2(n_77),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

AOI211xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_73),
.B(n_67),
.C(n_124),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_63),
.B1(n_55),
.B2(n_78),
.C(n_77),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_113),
.B(n_127),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_55),
.A3(n_95),
.B1(n_58),
.B2(n_60),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_97),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_58),
.A3(n_60),
.B1(n_78),
.B2(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_91),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_101),
.B1(n_89),
.B2(n_104),
.C(n_116),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_127),
.B(n_126),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_128),
.B(n_132),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_138),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_152),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_139),
.C(n_140),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_139),
.Y(n_161)
);

NOR3x1_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_10),
.C(n_11),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_138),
.Y(n_163)
);

NAND3x1_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_140),
.C(n_13),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_12),
.Y(n_166)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

NAND5xp2_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_101),
.C(n_14),
.D(n_16),
.E(n_17),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_97),
.B1(n_14),
.B2(n_12),
.C(n_19),
.Y(n_169)
);

NAND4xp75_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_97),
.C(n_90),
.D(n_107),
.Y(n_170)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_156),
.A3(n_159),
.B1(n_161),
.B2(n_97),
.C1(n_103),
.C2(n_88),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_97),
.Y(n_172)
);

OAI221xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_97),
.B1(n_88),
.B2(n_103),
.C(n_93),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_97),
.Y(n_174)
);

OAI322xp33_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_162),
.A3(n_168),
.B1(n_164),
.B2(n_170),
.C1(n_166),
.C2(n_103),
.Y(n_175)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_86),
.A3(n_88),
.B1(n_93),
.B2(n_109),
.C1(n_156),
.C2(n_69),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_109),
.B1(n_88),
.B2(n_86),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_109),
.B1(n_88),
.B2(n_86),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_88),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_86),
.B1(n_88),
.B2(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_86),
.B1(n_171),
.B2(n_177),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_179),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_177),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_184),
.B1(n_187),
.B2(n_183),
.Y(n_188)
);


endmodule