module fake_jpeg_13321_n_133 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_1),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_23),
.B1(n_17),
.B2(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_59),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_67),
.B1(n_28),
.B2(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_36),
.B1(n_34),
.B2(n_28),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_46),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_73),
.C(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_39),
.C(n_25),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_79),
.B1(n_42),
.B2(n_53),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_16),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_62),
.B1(n_22),
.B2(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_12),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_8),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_66),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_60),
.B1(n_57),
.B2(n_52),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_91),
.B1(n_68),
.B2(n_77),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_16),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_8),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_15),
.C(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_24),
.C(n_15),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_49),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_78),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_104),
.C(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_71),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_90),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_85),
.C(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_99),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_99),
.C(n_103),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_71),
.C(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_101),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_97),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_118),
.B(n_120),
.Y(n_122)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_110),
.B(n_106),
.C(n_107),
.D(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_116),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_9),
.B(n_27),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_22),
.A3(n_27),
.B1(n_51),
.B2(n_4),
.C1(n_1),
.C2(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_125),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_128),
.B(n_14),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_14),
.B(n_3),
.C(n_4),
.D(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_37),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_14),
.B1(n_4),
.B2(n_2),
.Y(n_131)
);

XNOR2x2_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);


endmodule