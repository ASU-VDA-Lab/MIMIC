module fake_jpeg_5235_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_13),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_13),
.B1(n_20),
.B2(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_44),
.B1(n_15),
.B2(n_18),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_45),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_28),
.B1(n_20),
.B2(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_33),
.B1(n_36),
.B2(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_68),
.B1(n_4),
.B2(n_9),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_32),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_25),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_25),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_17),
.B1(n_14),
.B2(n_33),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_81),
.B1(n_51),
.B2(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_24),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_36),
.B1(n_24),
.B2(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_1),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_54),
.B(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_66),
.B1(n_72),
.B2(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_72),
.B1(n_69),
.B2(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_74),
.B1(n_73),
.B2(n_70),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_74),
.B1(n_69),
.B2(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_110),
.B1(n_97),
.B2(n_90),
.Y(n_113)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_98),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_113),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_97),
.C(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.Y(n_120)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_56),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_110),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_111),
.B1(n_115),
.B2(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_70),
.B1(n_113),
.B2(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_85),
.Y(n_129)
);

OA21x2_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_100),
.B(n_104),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_120),
.C(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_133),
.C(n_12),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_106),
.B(n_4),
.C(n_11),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_129),
.C(n_112),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_135),
.B(n_136),
.C(n_1),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_12),
.B(n_2),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_2),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_2),
.Y(n_140)
);


endmodule