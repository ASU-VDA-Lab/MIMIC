module fake_jpeg_10894_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_87),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_1),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_0),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_85),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_48),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_86),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_0),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_1),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_19),
.Y(n_105)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_20),
.B1(n_46),
.B2(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_124),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_109),
.A2(n_96),
.B1(n_94),
.B2(n_84),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_31),
.B(n_21),
.C(n_24),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_17),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_53),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_118),
.A2(n_126),
.B1(n_131),
.B2(n_150),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_137),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_38),
.B1(n_47),
.B2(n_49),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_89),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_63),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_48),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_101),
.A2(n_49),
.B1(n_30),
.B2(n_20),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_49),
.B1(n_46),
.B2(n_31),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_151),
.A2(n_158),
.B1(n_162),
.B2(n_54),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_79),
.A2(n_46),
.B1(n_95),
.B2(n_19),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_99),
.A2(n_41),
.B1(n_21),
.B2(n_42),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_25),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_164),
.B(n_178),
.Y(n_253)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_23),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_169),
.A2(n_216),
.B(n_114),
.Y(n_225)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_79),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_173),
.B(n_183),
.Y(n_230)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_207),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_25),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_119),
.A2(n_24),
.B1(n_36),
.B2(n_37),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_179),
.A2(n_186),
.B1(n_196),
.B2(n_215),
.Y(n_239)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_119),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_187),
.A2(n_197),
.B1(n_208),
.B2(n_143),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_46),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_188),
.B(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_192),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_103),
.B(n_45),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_193),
.B(n_199),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_129),
.A2(n_45),
.B1(n_23),
.B2(n_19),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_150),
.A2(n_82),
.B1(n_74),
.B2(n_66),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

AO22x1_ASAP7_75t_SL g199 ( 
.A1(n_107),
.A2(n_23),
.B1(n_45),
.B2(n_60),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_109),
.A2(n_62),
.B1(n_61),
.B2(n_56),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_200),
.B(n_204),
.Y(n_275)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_46),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_1),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_205),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_1),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_218),
.C(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_118),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_158),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_213),
.Y(n_235)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_155),
.A2(n_51),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_2),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_112),
.Y(n_220)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_138),
.B1(n_147),
.B2(n_159),
.Y(n_250)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_117),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_153),
.B(n_2),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_225),
.B(n_17),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_168),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_242),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_166),
.B(n_130),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_243),
.B(n_246),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_166),
.B(n_130),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_185),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_164),
.A2(n_126),
.B1(n_151),
.B2(n_131),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_189),
.B1(n_200),
.B2(n_167),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_178),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_257),
.B(n_258),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_104),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_216),
.B(n_160),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_174),
.B(n_123),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_204),
.B(n_143),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_273),
.A2(n_149),
.B1(n_146),
.B2(n_144),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_216),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_7),
.Y(n_317)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_193),
.A3(n_223),
.B1(n_218),
.B2(n_206),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_284),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_181),
.C(n_170),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_169),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_283),
.A2(n_316),
.B1(n_262),
.B2(n_224),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_199),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_285),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_265),
.B1(n_273),
.B2(n_200),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_300),
.B1(n_303),
.B2(n_307),
.Y(n_339)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_211),
.B(n_222),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_293),
.B(n_227),
.Y(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g290 ( 
.A1(n_226),
.A2(n_199),
.B1(n_180),
.B2(n_214),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_291),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_192),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_239),
.A2(n_194),
.B(n_219),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_165),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_247),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_217),
.B1(n_194),
.B2(n_203),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_247),
.B(n_177),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_321),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_230),
.A2(n_221),
.B1(n_149),
.B2(n_146),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_240),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_313),
.B1(n_262),
.B2(n_233),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_229),
.A2(n_220),
.B1(n_212),
.B2(n_172),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_267),
.A2(n_172),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g342 ( 
.A1(n_310),
.A2(n_322),
.B1(n_316),
.B2(n_307),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_311),
.A2(n_234),
.B(n_261),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_241),
.B(n_2),
.C(n_5),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_231),
.CI(n_227),
.CON(n_329),
.SN(n_329)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_241),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_252),
.B(n_267),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_314),
.B(n_315),
.Y(n_345)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_266),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_317),
.B(n_312),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_232),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_318),
.A2(n_13),
.B1(n_16),
.B2(n_295),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_272),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_320),
.B(n_323),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_228),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_232),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_338),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_331),
.B1(n_354),
.B2(n_297),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_286),
.A2(n_233),
.B1(n_238),
.B2(n_236),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_236),
.A3(n_238),
.B1(n_234),
.B2(n_228),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_343),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_342),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_288),
.A2(n_261),
.B(n_260),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_337),
.B(n_350),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_245),
.B(n_256),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_294),
.B(n_260),
.CI(n_255),
.CON(n_338),
.SN(n_338)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_349),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_291),
.A2(n_264),
.A3(n_255),
.B1(n_256),
.B2(n_245),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_301),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_264),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_299),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_358),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_283),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_295),
.A2(n_11),
.B(n_12),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_356),
.A2(n_363),
.B(n_285),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_292),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_359),
.A2(n_360),
.B1(n_309),
.B2(n_300),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_278),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_362),
.A2(n_311),
.B1(n_313),
.B2(n_297),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_293),
.A2(n_311),
.B(n_281),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_280),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_341),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_368),
.B(n_373),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_369),
.A2(n_371),
.B1(n_383),
.B2(n_399),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_324),
.B(n_277),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_378),
.C(n_387),
.Y(n_409)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_315),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_340),
.A2(n_306),
.B1(n_290),
.B2(n_276),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_379),
.A2(n_350),
.B(n_356),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_392),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_339),
.A2(n_290),
.B1(n_279),
.B2(n_296),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_290),
.Y(n_385)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_282),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_308),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_388),
.B(n_394),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_289),
.Y(n_389)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_321),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_320),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_393),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_326),
.B(n_303),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_323),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_395),
.Y(n_402)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_396),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_397),
.A2(n_384),
.B(n_325),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_337),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_400),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_339),
.A2(n_287),
.B1(n_330),
.B2(n_331),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_343),
.B(n_332),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_416),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_386),
.A2(n_354),
.B1(n_350),
.B2(n_338),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_404),
.A2(n_427),
.B1(n_430),
.B2(n_397),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_372),
.A2(n_353),
.B1(n_358),
.B2(n_364),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_379),
.B1(n_382),
.B2(n_371),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_392),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_408),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_390),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_345),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_394),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_414),
.A2(n_431),
.B(n_385),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g415 ( 
.A(n_373),
.B(n_338),
.CI(n_329),
.CON(n_415),
.SN(n_415)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_415),
.B(n_359),
.CI(n_380),
.CON(n_457),
.SN(n_457)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_375),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_429),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_386),
.A2(n_348),
.B1(n_329),
.B2(n_336),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_383),
.A2(n_327),
.B1(n_336),
.B2(n_362),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_367),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_386),
.A2(n_364),
.B1(n_346),
.B2(n_355),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_384),
.A2(n_363),
.B(n_335),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_432),
.A2(n_439),
.B1(n_441),
.B2(n_449),
.Y(n_463)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_412),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_444),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_374),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_451),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_387),
.C(n_388),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_440),
.C(n_446),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_422),
.A2(n_399),
.B1(n_369),
.B2(n_400),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_376),
.C(n_370),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_389),
.Y(n_442)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_443),
.B(n_445),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_410),
.B(n_381),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_377),
.C(n_395),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_393),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_403),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_401),
.A2(n_367),
.B(n_366),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_419),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_365),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_361),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_456),
.Y(n_474)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_453),
.Y(n_468)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_396),
.C(n_391),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_425),
.C(n_426),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_360),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_415),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_457),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_357),
.Y(n_461)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_455),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_465),
.B(n_447),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_431),
.C(n_423),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_472),
.C(n_475),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_436),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_470),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_428),
.B1(n_420),
.B2(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_420),
.C(n_430),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_414),
.C(n_424),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_478),
.Y(n_488)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_446),
.B(n_415),
.CI(n_421),
.CON(n_478),
.SN(n_478)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_494),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_440),
.C(n_434),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_481),
.B(n_486),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_434),
.C(n_450),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_474),
.C(n_465),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_487),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_469),
.A2(n_441),
.B1(n_429),
.B2(n_424),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_491),
.B1(n_493),
.B2(n_488),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_448),
.C(n_445),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_452),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_464),
.Y(n_489)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_475),
.A2(n_466),
.B1(n_458),
.B2(n_467),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_444),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_457),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_495),
.Y(n_498)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_497),
.Y(n_514)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_501),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_463),
.C(n_474),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_503),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_477),
.C(n_456),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_473),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_346),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_477),
.C(n_442),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_425),
.C(n_426),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_507),
.A2(n_488),
.B(n_494),
.Y(n_509)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_509),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_496),
.A2(n_404),
.B1(n_402),
.B2(n_480),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_511),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_468),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_512),
.A2(n_515),
.B(n_499),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_512),
.B1(n_516),
.B2(n_503),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_490),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_521),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_517),
.A2(n_498),
.B(n_514),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_509),
.A2(n_500),
.B1(n_501),
.B2(n_505),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_522),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_522),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_511),
.C(n_520),
.Y(n_527)
);

A2O1A1O1Ixp25_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_528),
.B(n_524),
.C(n_508),
.D(n_347),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_SL g528 ( 
.A1(n_525),
.A2(n_518),
.B(n_510),
.C(n_508),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_355),
.B(n_333),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_333),
.B(n_347),
.Y(n_531)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_531),
.A2(n_334),
.B(n_342),
.C(n_357),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_342),
.Y(n_533)
);


endmodule