module real_aes_18245_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_850, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_850;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_626;
wire n_292;
wire n_400;
wire n_539;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AND2x4_ASAP7_75t_L g120 ( .A(n_0), .B(n_121), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_1), .A2(n_3), .B1(n_143), .B2(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_2), .A2(n_46), .B1(n_150), .B2(n_256), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_4), .A2(n_27), .B1(n_221), .B2(n_256), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_5), .A2(n_17), .B1(n_140), .B2(n_189), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_6), .A2(n_63), .B1(n_168), .B2(n_223), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_7), .A2(n_18), .B1(n_150), .B2(n_172), .Y(n_534) );
INVx1_ASAP7_75t_L g121 ( .A(n_8), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_9), .A2(n_38), .B1(n_559), .B2(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_9), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_10), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_11), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_12), .A2(n_20), .B1(n_167), .B2(n_170), .Y(n_166) );
OR2x2_ASAP7_75t_L g111 ( .A(n_13), .B(n_42), .Y(n_111) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_15), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_16), .Y(n_838) );
OAI22xp5_ASAP7_75t_SL g811 ( .A1(n_19), .A2(n_75), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_19), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_21), .B(n_819), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_22), .A2(n_101), .B1(n_140), .B2(n_143), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_23), .A2(n_43), .B1(n_184), .B2(n_186), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_24), .B(n_141), .Y(n_234) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_25), .A2(n_59), .B(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_26), .A2(n_799), .B1(n_803), .B2(n_804), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_26), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_28), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_29), .Y(n_629) );
INVx4_ASAP7_75t_R g546 ( .A(n_30), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_31), .B(n_147), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_32), .A2(n_50), .B1(n_200), .B2(n_202), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_33), .A2(n_70), .B1(n_801), .B2(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_33), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_34), .A2(n_56), .B1(n_140), .B2(n_202), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_35), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_36), .B(n_184), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_37), .Y(n_247) );
INVx1_ASAP7_75t_L g559 ( .A(n_38), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_39), .B(n_256), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_SL g495 ( .A1(n_40), .A2(n_146), .B(n_150), .C(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_41), .A2(n_57), .B1(n_150), .B2(n_202), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_44), .A2(n_89), .B1(n_150), .B2(n_220), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_45), .A2(n_49), .B1(n_150), .B2(n_172), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_47), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_48), .A2(n_61), .B1(n_140), .B2(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g581 ( .A(n_51), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_52), .B(n_150), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_53), .Y(n_521) );
INVx2_ASAP7_75t_L g119 ( .A(n_54), .Y(n_119) );
BUFx3_ASAP7_75t_L g110 ( .A(n_55), .Y(n_110) );
INVx1_ASAP7_75t_L g822 ( .A(n_55), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_58), .A2(n_90), .B1(n_150), .B2(n_202), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_60), .Y(n_547) );
XNOR2xp5_ASAP7_75t_SL g799 ( .A(n_62), .B(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_64), .A2(n_78), .B1(n_149), .B2(n_200), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_65), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_66), .A2(n_80), .B1(n_150), .B2(n_172), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_67), .A2(n_100), .B1(n_140), .B2(n_170), .Y(n_244) );
AND2x4_ASAP7_75t_L g136 ( .A(n_68), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g159 ( .A(n_69), .Y(n_159) );
INVx1_ASAP7_75t_L g801 ( .A(n_70), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_71), .A2(n_92), .B1(n_200), .B2(n_202), .Y(n_555) );
AO22x1_ASAP7_75t_L g512 ( .A1(n_72), .A2(n_79), .B1(n_186), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g137 ( .A(n_73), .Y(n_137) );
AND2x2_ASAP7_75t_L g499 ( .A(n_74), .B(n_240), .Y(n_499) );
INVx1_ASAP7_75t_L g812 ( .A(n_75), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_76), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_77), .B(n_223), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_81), .B(n_256), .Y(n_522) );
INVx2_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_83), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_84), .B(n_240), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_85), .A2(n_99), .B1(n_202), .B2(n_223), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_86), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_87), .B(n_157), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_88), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_91), .B(n_240), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_93), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_94), .B(n_240), .Y(n_518) );
INVx1_ASAP7_75t_L g115 ( .A(n_95), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_95), .B(n_821), .Y(n_820) );
NAND2xp33_ASAP7_75t_L g237 ( .A(n_96), .B(n_141), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_97), .A2(n_174), .B(n_223), .C(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g548 ( .A(n_98), .B(n_549), .Y(n_548) );
NAND2xp33_ASAP7_75t_L g526 ( .A(n_102), .B(n_185), .Y(n_526) );
AOI211xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_122), .B(n_807), .C(n_837), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx4_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx4f_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_112), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g113 ( .A(n_109), .B(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g823 ( .A(n_111), .Y(n_823) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
AND2x2_ASAP7_75t_L g840 ( .A(n_113), .B(n_841), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_114), .Y(n_797) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g479 ( .A(n_115), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_116), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_117), .B(n_120), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_118), .B(n_835), .Y(n_834) );
INVx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_119), .B(n_848), .Y(n_847) );
INVx2_ASAP7_75t_SL g836 ( .A(n_120), .Y(n_836) );
INVxp67_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_798), .B1(n_805), .B2(n_806), .Y(n_123) );
INVx1_ASAP7_75t_L g805 ( .A(n_124), .Y(n_805) );
OAI22x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_477), .B1(n_480), .B2(n_797), .Y(n_124) );
INVx2_ASAP7_75t_L g814 ( .A(n_125), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_125), .B(n_816), .Y(n_815) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_386), .Y(n_125) );
NOR2x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_325), .Y(n_126) );
NAND4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_276), .C(n_295), .D(n_306), .Y(n_127) );
O2A1O1Ixp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_207), .B(n_214), .C(n_248), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_179), .Y(n_129) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_130), .B(n_341), .C(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g422 ( .A(n_130), .B(n_304), .Y(n_422) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
AND2x2_ASAP7_75t_L g266 ( .A(n_131), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g284 ( .A(n_131), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g301 ( .A(n_131), .Y(n_301) );
AND2x2_ASAP7_75t_L g346 ( .A(n_131), .B(n_181), .Y(n_346) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g211 ( .A(n_132), .Y(n_211) );
AND2x4_ASAP7_75t_L g294 ( .A(n_132), .B(n_285), .Y(n_294) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .A3(n_154), .B(n_160), .Y(n_132) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_133), .A2(n_175), .A3(n_243), .B(n_246), .Y(n_242) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_134), .A2(n_541), .B(n_544), .Y(n_540) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AO31x2_ASAP7_75t_L g164 ( .A1(n_135), .A2(n_165), .A3(n_175), .B(n_177), .Y(n_164) );
AO31x2_ASAP7_75t_L g181 ( .A1(n_135), .A2(n_182), .A3(n_191), .B(n_193), .Y(n_181) );
AO31x2_ASAP7_75t_L g253 ( .A1(n_135), .A2(n_254), .A3(n_258), .B(n_259), .Y(n_253) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_135), .A2(n_162), .A3(n_533), .B(n_536), .Y(n_532) );
BUFx10_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
INVx1_ASAP7_75t_L g498 ( .A(n_136), .Y(n_498) );
BUFx10_ASAP7_75t_L g530 ( .A(n_136), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B1(n_148), .B2(n_151), .Y(n_138) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_141), .Y(n_513) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g144 ( .A(n_142), .Y(n_144) );
INVx3_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
INVx1_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
INVx1_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_142), .Y(n_202) );
INVx2_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
INVx1_ASAP7_75t_L g223 ( .A(n_142), .Y(n_223) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_142), .Y(n_256) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_144), .B(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_145), .A2(n_166), .B1(n_171), .B2(n_173), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_145), .A2(n_151), .B1(n_183), .B2(n_188), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_145), .A2(n_151), .B1(n_199), .B2(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_145), .A2(n_219), .B1(n_222), .B2(n_224), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_145), .A2(n_236), .B(n_237), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_145), .A2(n_173), .B1(n_244), .B2(n_245), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_145), .A2(n_151), .B1(n_255), .B2(n_257), .Y(n_254) );
OAI22x1_ASAP7_75t_L g533 ( .A1(n_145), .A2(n_224), .B1(n_534), .B2(n_535), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_145), .A2(n_224), .B1(n_555), .B2(n_556), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_145), .A2(n_508), .B1(n_626), .B2(n_627), .Y(n_625) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_146), .A2(n_172), .B(n_233), .C(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_146), .B(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_146), .A2(n_526), .B(n_527), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_146), .A2(n_507), .B(n_512), .C(n_515), .Y(n_567) );
BUFx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx1_ASAP7_75t_L g494 ( .A(n_147), .Y(n_494) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVx4_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g508 ( .A(n_152), .Y(n_508) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g524 ( .A(n_153), .Y(n_524) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_154), .A2(n_198), .A3(n_203), .B(n_205), .Y(n_197) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_154), .A2(n_540), .B(n_548), .Y(n_539) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_SL g177 ( .A(n_156), .B(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_156), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
INVx2_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
OAI21xp33_ASAP7_75t_L g515 ( .A1(n_157), .A2(n_498), .B(n_510), .Y(n_515) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_162), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g212 ( .A(n_163), .B(n_213), .Y(n_212) );
AND2x4_ASAP7_75t_L g269 ( .A(n_163), .B(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_163), .Y(n_292) );
INVx1_ASAP7_75t_L g303 ( .A(n_163), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_163), .B(n_195), .Y(n_312) );
INVx2_ASAP7_75t_L g319 ( .A(n_163), .Y(n_319) );
INVx4_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g264 ( .A(n_164), .B(n_181), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_164), .B(n_271), .Y(n_337) );
AND2x2_ASAP7_75t_L g345 ( .A(n_164), .B(n_197), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_164), .B(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g398 ( .A(n_164), .Y(n_398) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_169), .B(n_543), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_172), .A2(n_521), .B(n_522), .C(n_523), .Y(n_520) );
INVx1_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g224 ( .A(n_174), .Y(n_224) );
AOI21x1_ASAP7_75t_L g486 ( .A1(n_175), .A2(n_487), .B(n_499), .Y(n_486) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_175), .A2(n_203), .A3(n_554), .B(n_558), .Y(n_553) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_176), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g549 ( .A(n_176), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_176), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_176), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g414 ( .A(n_180), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_195), .Y(n_180) );
INVx1_ASAP7_75t_L g213 ( .A(n_181), .Y(n_213) );
INVx1_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
INVx2_ASAP7_75t_L g305 ( .A(n_181), .Y(n_305) );
OR2x2_ASAP7_75t_L g309 ( .A(n_181), .B(n_197), .Y(n_309) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_181), .Y(n_358) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g200 ( .A(n_185), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_185), .A2(n_190), .B1(n_546), .B2(n_547), .Y(n_545) );
OAI21xp33_ASAP7_75t_SL g577 ( .A1(n_186), .A2(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_191), .A2(n_203), .A3(n_218), .B(n_225), .Y(n_217) );
BUFx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_192), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_SL g230 ( .A(n_192), .Y(n_230) );
INVx4_ASAP7_75t_L g240 ( .A(n_192), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_192), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_192), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g585 ( .A(n_192), .B(n_530), .Y(n_585) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g331 ( .A(n_196), .B(n_211), .Y(n_331) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
INVx2_ASAP7_75t_L g285 ( .A(n_197), .Y(n_285) );
AND2x4_ASAP7_75t_L g304 ( .A(n_197), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g392 ( .A(n_197), .Y(n_392) );
INVx2_ASAP7_75t_L g557 ( .A(n_202), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_202), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_SL g238 ( .A(n_204), .Y(n_238) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g310 ( .A(n_210), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_210), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g373 ( .A(n_211), .Y(n_373) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2x1_ASAP7_75t_L g215 ( .A(n_216), .B(n_227), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_216), .B(n_228), .Y(n_323) );
INVx1_ASAP7_75t_L g421 ( .A(n_216), .Y(n_421) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g261 ( .A(n_217), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g275 ( .A(n_217), .B(n_253), .Y(n_275) );
AND2x4_ASAP7_75t_L g298 ( .A(n_217), .B(n_241), .Y(n_298) );
INVx2_ASAP7_75t_L g315 ( .A(n_217), .Y(n_315) );
AND2x2_ASAP7_75t_L g341 ( .A(n_217), .B(n_242), .Y(n_341) );
INVx1_ASAP7_75t_L g406 ( .A(n_217), .Y(n_406) );
INVx2_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_221), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_224), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g366 ( .A(n_227), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
AND2x2_ASAP7_75t_L g332 ( .A(n_228), .B(n_289), .Y(n_332) );
AND2x4_ASAP7_75t_L g348 ( .A(n_228), .B(n_315), .Y(n_348) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g342 ( .A(n_229), .Y(n_342) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_263) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_235), .B(n_238), .Y(n_231) );
INVx2_ASAP7_75t_L g258 ( .A(n_240), .Y(n_258) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_240), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g274 ( .A(n_241), .Y(n_274) );
INVx3_ASAP7_75t_L g280 ( .A(n_241), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_241), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_241), .B(n_409), .Y(n_408) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g314 ( .A(n_242), .B(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g438 ( .A(n_242), .Y(n_438) );
OAI33xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_264), .A3(n_265), .B1(n_266), .B2(n_268), .B3(n_272), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NOR2x1_ASAP7_75t_L g250 ( .A(n_251), .B(n_261), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g372 ( .A(n_252), .B(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g281 ( .A(n_253), .B(n_263), .Y(n_281) );
INVx2_ASAP7_75t_L g289 ( .A(n_253), .Y(n_289) );
INVx1_ASAP7_75t_L g297 ( .A(n_253), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_256), .B(n_490), .Y(n_489) );
AO31x2_ASAP7_75t_L g624 ( .A1(n_258), .A2(n_530), .A3(n_625), .B(n_628), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_261), .A2(n_317), .B1(n_320), .B2(n_324), .Y(n_316) );
OR2x2_ASAP7_75t_L g456 ( .A(n_261), .B(n_274), .Y(n_456) );
AND2x4_ASAP7_75t_L g360 ( .A(n_262), .B(n_322), .Y(n_360) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_263), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_264), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g324 ( .A(n_264), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_264), .B(n_300), .Y(n_402) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g375 ( .A(n_266), .Y(n_375) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g433 ( .A(n_269), .B(n_301), .Y(n_433) );
NAND2x1_ASAP7_75t_L g451 ( .A(n_269), .B(n_300), .Y(n_451) );
AND2x2_ASAP7_75t_L g475 ( .A(n_269), .B(n_294), .Y(n_475) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g465 ( .A(n_273), .B(n_342), .Y(n_465) );
NOR2x1p5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g399 ( .A(n_274), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g367 ( .A(n_275), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_282), .B1(n_286), .B2(n_290), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g374 ( .A(n_279), .B(n_342), .Y(n_374) );
AND2x2_ASAP7_75t_L g411 ( .A(n_279), .B(n_360), .Y(n_411) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g286 ( .A(n_280), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_280), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g452 ( .A(n_280), .B(n_281), .Y(n_452) );
AND2x2_ASAP7_75t_L g313 ( .A(n_281), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g432 ( .A(n_281), .B(n_298), .Y(n_432) );
AND2x2_ASAP7_75t_L g476 ( .A(n_281), .B(n_341), .Y(n_476) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_286), .A2(n_411), .B1(n_412), .B2(n_415), .C1(n_417), .C2(n_418), .Y(n_410) );
AND2x2_ASAP7_75t_L g333 ( .A(n_287), .B(n_301), .Y(n_333) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g364 ( .A(n_288), .Y(n_364) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_288), .Y(n_409) );
INVx2_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g379 ( .A(n_292), .Y(n_379) );
INVx2_ASAP7_75t_L g385 ( .A(n_293), .Y(n_385) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g369 ( .A(n_294), .B(n_358), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x4_ASAP7_75t_L g400 ( .A(n_297), .B(n_348), .Y(n_400) );
INVx2_ASAP7_75t_L g447 ( .A(n_297), .Y(n_447) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g390 ( .A(n_301), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g424 ( .A(n_301), .B(n_309), .Y(n_424) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_304), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g436 ( .A(n_304), .B(n_352), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .B(n_313), .C(n_316), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OR2x2_ASAP7_75t_L g317 ( .A(n_309), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g353 ( .A(n_309), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_310), .B(n_345), .Y(n_449) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g425 ( .A(n_312), .B(n_394), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_314), .B(n_364), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_314), .A2(n_330), .B1(n_372), .B2(n_374), .Y(n_371) );
AND2x2_ASAP7_75t_L g377 ( .A(n_314), .B(n_342), .Y(n_377) );
AND2x2_ASAP7_75t_L g446 ( .A(n_314), .B(n_447), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_317), .A2(n_419), .B(n_440), .C(n_443), .Y(n_439) );
INVx2_ASAP7_75t_L g352 ( .A(n_319), .Y(n_352) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g430 ( .A(n_322), .Y(n_430) );
INVx1_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_324), .A2(n_371), .B1(n_375), .B2(n_376), .Y(n_370) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_338), .C(n_361), .Y(n_325) );
AO22x1_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_332), .B1(n_333), .B2(n_334), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_331), .Y(n_464) );
OR2x2_ASAP7_75t_L g471 ( .A(n_331), .B(n_352), .Y(n_471) );
AND2x2_ASAP7_75t_L g383 ( .A(n_332), .B(n_341), .Y(n_383) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g459 ( .A(n_337), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_343), .C(n_349), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
AND2x4_ASAP7_75t_SL g417 ( .A(n_341), .B(n_360), .Y(n_417) );
INVx1_ASAP7_75t_SL g428 ( .A(n_341), .Y(n_428) );
OR2x2_ASAP7_75t_L g380 ( .A(n_342), .B(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x4_ASAP7_75t_L g357 ( .A(n_345), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g415 ( .A(n_346), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g437 ( .A(n_348), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g462 ( .A(n_348), .B(n_442), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B1(n_356), .B2(n_359), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x4_ASAP7_75t_L g397 ( .A(n_353), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g419 ( .A(n_353), .Y(n_419) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g474 ( .A(n_357), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_370), .C(n_378), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_368), .Y(n_362) );
INVx1_ASAP7_75t_L g443 ( .A(n_364), .Y(n_443) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_369), .A2(n_467), .B1(n_470), .B2(n_472), .C1(n_474), .C2(n_476), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_372), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_382), .C(n_384), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_444), .Y(n_386) );
NAND4xp25_ASAP7_75t_L g387 ( .A(n_388), .B(n_410), .C(n_420), .D(n_431), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_399), .B1(n_401), .B2(n_403), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .C(n_396), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_390), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_394), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g441 ( .A(n_406), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_408), .Y(n_473) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g468 ( .A(n_417), .Y(n_468) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_423), .C(n_429), .Y(n_420) );
AOI21xp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_425), .B(n_426), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_424), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_434), .B2(n_437), .C(n_439), .Y(n_431) );
INVx1_ASAP7_75t_L g469 ( .A(n_432), .Y(n_469) );
AOI31xp33_ASAP7_75t_L g453 ( .A1(n_435), .A2(n_454), .A3(n_455), .B(n_456), .Y(n_453) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_438), .Y(n_442) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_457), .C(n_466), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_450), .B2(n_452), .C(n_453), .Y(n_445) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g454 ( .A(n_452), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B1(n_463), .B2(n_465), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_697), .Y(n_481) );
NAND3xp33_ASAP7_75t_SL g482 ( .A(n_483), .B(n_600), .C(n_659), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_500), .B1(n_587), .B2(n_593), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g656 ( .A(n_485), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_485), .B(n_574), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_485), .B(n_620), .Y(n_767) );
AND2x2_ASAP7_75t_L g773 ( .A(n_485), .B(n_599), .Y(n_773) );
INVxp67_ASAP7_75t_L g778 ( .A(n_485), .Y(n_778) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g591 ( .A(n_486), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_495), .B(n_498), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_491), .B(n_493), .Y(n_488) );
BUFx4f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_494), .B(n_581), .Y(n_580) );
OAI21xp5_ASAP7_75t_SL g500 ( .A1(n_501), .A2(n_550), .B(n_560), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_531), .Y(n_502) );
INVx1_ASAP7_75t_L g694 ( .A(n_503), .Y(n_694) );
AND2x2_ASAP7_75t_L g723 ( .A(n_503), .B(n_685), .Y(n_723) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_516), .Y(n_503) );
AND2x2_ASAP7_75t_L g617 ( .A(n_504), .B(n_539), .Y(n_617) );
INVx1_ASAP7_75t_L g672 ( .A(n_504), .Y(n_672) );
AND2x2_ASAP7_75t_L g722 ( .A(n_504), .B(n_538), .Y(n_722) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g597 ( .A(n_505), .B(n_538), .Y(n_597) );
AND2x4_ASAP7_75t_L g741 ( .A(n_505), .B(n_539), .Y(n_741) );
AOI21x1_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_511), .B(n_514), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI21x1_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_510), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_508), .A2(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g666 ( .A(n_516), .Y(n_666) );
AND2x2_ASAP7_75t_L g735 ( .A(n_516), .B(n_539), .Y(n_735) );
AND2x2_ASAP7_75t_L g742 ( .A(n_516), .B(n_568), .Y(n_742) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
BUFx3_ASAP7_75t_L g599 ( .A(n_517), .Y(n_599) );
AND2x2_ASAP7_75t_L g610 ( .A(n_517), .B(n_596), .Y(n_610) );
AND2x2_ASAP7_75t_L g673 ( .A(n_517), .B(n_532), .Y(n_673) );
AND2x2_ASAP7_75t_L g678 ( .A(n_517), .B(n_539), .Y(n_678) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_525), .B(n_528), .Y(n_519) );
INVx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_531), .B(n_684), .Y(n_786) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_538), .Y(n_531) );
INVx2_ASAP7_75t_L g568 ( .A(n_532), .Y(n_568) );
OR2x2_ASAP7_75t_L g571 ( .A(n_532), .B(n_539), .Y(n_571) );
INVx2_ASAP7_75t_L g596 ( .A(n_532), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_532), .B(n_566), .Y(n_612) );
AND2x2_ASAP7_75t_L g685 ( .A(n_532), .B(n_539), .Y(n_685) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g613 ( .A(n_539), .Y(n_613) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_551), .B(n_648), .Y(n_794) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g606 ( .A(n_552), .Y(n_606) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g586 ( .A(n_553), .Y(n_586) );
AND2x2_ASAP7_75t_L g592 ( .A(n_553), .B(n_574), .Y(n_592) );
INVx1_ASAP7_75t_L g640 ( .A(n_553), .Y(n_640) );
OR2x2_ASAP7_75t_L g645 ( .A(n_553), .B(n_624), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_553), .B(n_624), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_553), .B(n_623), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_553), .B(n_591), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_559), .A2(n_838), .B1(n_839), .B2(n_844), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_569), .B(n_572), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
OR2x2_ASAP7_75t_L g570 ( .A(n_563), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g721 ( .A(n_563), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g751 ( .A(n_563), .B(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_564), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g719 ( .A(n_564), .Y(n_719) );
OR2x2_ASAP7_75t_L g632 ( .A(n_565), .B(n_633), .Y(n_632) );
INVxp33_ASAP7_75t_L g750 ( .A(n_565), .Y(n_750) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx2_ASAP7_75t_L g654 ( .A(n_566), .Y(n_654) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g716 ( .A1(n_570), .A2(n_641), .B1(n_646), .B2(n_717), .C(n_720), .Y(n_716) );
OR2x2_ASAP7_75t_L g703 ( .A(n_571), .B(n_654), .Y(n_703) );
INVx2_ASAP7_75t_L g752 ( .A(n_571), .Y(n_752) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g652 ( .A(n_573), .Y(n_652) );
OR2x2_ASAP7_75t_L g655 ( .A(n_573), .B(n_656), .Y(n_655) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_573), .Y(n_696) );
OR2x2_ASAP7_75t_L g709 ( .A(n_573), .B(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_586), .Y(n_573) );
NAND2x1p5_ASAP7_75t_SL g605 ( .A(n_574), .B(n_590), .Y(n_605) );
INVx3_ASAP7_75t_L g620 ( .A(n_574), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_574), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
AND2x2_ASAP7_75t_L g724 ( .A(n_574), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g731 ( .A(n_574), .B(n_638), .Y(n_731) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_582), .B(n_585), .Y(n_576) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
AND2x2_ASAP7_75t_L g783 ( .A(n_588), .B(n_642), .Y(n_783) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g687 ( .A(n_590), .B(n_657), .Y(n_687) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g622 ( .A(n_591), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g648 ( .A(n_591), .B(n_624), .Y(n_648) );
AND2x4_ASAP7_75t_L g745 ( .A(n_592), .B(n_715), .Y(n_745) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_598), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g664 ( .A(n_597), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_598), .B(n_685), .Y(n_769) );
AND2x2_ASAP7_75t_L g776 ( .A(n_598), .B(n_736), .Y(n_776) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx2_ASAP7_75t_L g701 ( .A(n_599), .Y(n_701) );
AOI321xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_614), .A3(n_630), .B1(n_631), .B2(n_634), .C(n_649), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_611), .Y(n_601) );
AOI21xp33_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_607), .B(n_609), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_604), .A2(n_615), .B(n_618), .Y(n_614) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OR2x2_ASAP7_75t_L g713 ( .A(n_605), .B(n_645), .Y(n_713) );
INVx1_ASAP7_75t_L g705 ( .A(n_606), .Y(n_705) );
INVx2_ASAP7_75t_L g690 ( .A(n_607), .Y(n_690) );
OAI32xp33_ASAP7_75t_L g793 ( .A1(n_607), .A2(n_755), .A3(n_766), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g708 ( .A(n_608), .Y(n_708) );
INVx1_ASAP7_75t_L g658 ( .A(n_609), .Y(n_658) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_SL g746 ( .A(n_610), .B(n_653), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_611), .B(n_615), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_611), .A2(n_687), .B1(n_748), .B2(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g736 ( .A(n_612), .Y(n_736) );
INVx1_ASAP7_75t_L g633 ( .A(n_613), .Y(n_633) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g718 ( .A(n_617), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_618), .B(n_635), .C(n_641), .D(n_646), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVxp67_ASAP7_75t_L g660 ( .A(n_619), .Y(n_660) );
AND2x2_ASAP7_75t_L g739 ( .A(n_619), .B(n_648), .Y(n_739) );
OR2x2_ASAP7_75t_L g748 ( .A(n_619), .B(n_622), .Y(n_748) );
AND2x2_ASAP7_75t_L g772 ( .A(n_619), .B(n_644), .Y(n_772) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g686 ( .A(n_620), .B(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_L g693 ( .A(n_620), .B(n_640), .Y(n_693) );
INVx1_ASAP7_75t_L g757 ( .A(n_621), .Y(n_757) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g665 ( .A(n_622), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g715 ( .A(n_622), .Y(n_715) );
INVx1_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g638 ( .A(n_624), .Y(n_638) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AND2x4_ASAP7_75t_L g651 ( .A(n_637), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g692 ( .A(n_637), .Y(n_692) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_639), .Y(n_756) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_643), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g733 ( .A(n_645), .Y(n_733) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g710 ( .A(n_648), .Y(n_710) );
AND2x2_ASAP7_75t_L g753 ( .A(n_648), .B(n_693), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_653), .B(n_655), .C(n_658), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g764 ( .A(n_653), .B(n_742), .Y(n_764) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g668 ( .A(n_656), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B(n_674), .C(n_688), .Y(n_659) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_667), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_663), .A2(n_771), .B(n_774), .Y(n_770) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g684 ( .A(n_666), .Y(n_684) );
AND2x2_ASAP7_75t_L g744 ( .A(n_666), .B(n_741), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g763 ( .A(n_671), .Y(n_763) );
AND2x2_ASAP7_75t_L g789 ( .A(n_671), .B(n_752), .Y(n_789) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_672), .Y(n_677) );
INVx2_ASAP7_75t_L g728 ( .A(n_673), .Y(n_728) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_673), .B(n_763), .Y(n_762) );
AOI33xp33_ASAP7_75t_L g780 ( .A1(n_673), .A2(n_693), .A3(n_731), .B1(n_741), .B2(n_773), .B3(n_850), .Y(n_780) );
OAI22xp33_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_679), .B1(n_682), .B2(n_686), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x2_ASAP7_75t_L g707 ( .A(n_678), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_679), .B(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
OR2x2_ASAP7_75t_L g792 ( .A(n_681), .B(n_726), .Y(n_792) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
OAI22xp33_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_691), .B1(n_694), .B2(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_692), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_692), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g714 ( .A(n_693), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g779 ( .A(n_693), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_758), .Y(n_697) );
NOR4xp25_ASAP7_75t_L g698 ( .A(n_699), .B(n_716), .C(n_737), .D(n_754), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B1(n_706), .B2(n_709), .C(n_711), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_SL g754 ( .A1(n_700), .A2(n_755), .B(n_756), .C(n_757), .Y(n_754) );
NAND2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g787 ( .A(n_703), .Y(n_787) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_707), .A2(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_723), .B(n_724), .C(n_727), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g766 ( .A(n_726), .B(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_726), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_732), .B2(n_734), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
OAI211xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B(n_743), .C(n_749), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g788 ( .A1(n_741), .A2(n_789), .B1(n_790), .B2(n_791), .C(n_793), .Y(n_788) );
INVx3_ASAP7_75t_L g796 ( .A(n_741), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_743) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g755 ( .A(n_752), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_781), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_770), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_764), .B(n_765), .C(n_768), .Y(n_760) );
INVx2_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_764), .B(n_785), .C(n_787), .Y(n_784) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_777), .B(n_780), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OR2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B(n_788), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g806 ( .A(n_798), .Y(n_806) );
INVx1_ASAP7_75t_L g804 ( .A(n_799), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_830), .Y(n_807) );
NOR2x1_ASAP7_75t_L g808 ( .A(n_809), .B(n_827), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_817), .B(n_826), .Y(n_809) );
AOI21x1_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_814), .B(n_815), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_811), .Y(n_816) );
AOI211xp5_ASAP7_75t_SL g827 ( .A1(n_811), .A2(n_814), .B(n_815), .C(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_824), .Y(n_817) );
INVx4_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_819), .B(n_824), .Y(n_829) );
CKINVDCx8_ASAP7_75t_R g843 ( .A(n_819), .Y(n_843) );
INVx3_ASAP7_75t_L g848 ( .A(n_819), .Y(n_848) );
AND2x6_ASAP7_75t_SL g819 ( .A(n_820), .B(n_823), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
INVx4_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
BUFx3_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OR2x4_ASAP7_75t_L g846 ( .A(n_835), .B(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx3_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
CKINVDCx6p67_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
BUFx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
endmodule