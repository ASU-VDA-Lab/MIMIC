module fake_jpeg_7784_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_8),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_33),
.Y(n_71)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_19),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_63),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_29),
.B1(n_35),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_59),
.B1(n_64),
.B2(n_78),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_29),
.B1(n_35),
.B2(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_73),
.B(n_47),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_36),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_83),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_33),
.B1(n_21),
.B2(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_34),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_27),
.B1(n_32),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_85),
.B1(n_28),
.B2(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_22),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_28),
.B(n_22),
.C(n_44),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_46),
.B1(n_48),
.B2(n_45),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_88),
.A2(n_125),
.B1(n_4),
.B2(n_5),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_102),
.Y(n_137)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_100),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_18),
.B1(n_65),
.B2(n_80),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_111),
.B(n_22),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_24),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_104),
.Y(n_148)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_120),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_12),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_112),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_49),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_0),
.C(n_1),
.Y(n_145)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_10),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_2),
.Y(n_154)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_65),
.Y(n_119)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_30),
.B1(n_31),
.B2(n_22),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_70),
.A2(n_68),
.B1(n_74),
.B2(n_54),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_31),
.B1(n_30),
.B2(n_2),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_68),
.B1(n_74),
.B2(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_22),
.B(n_31),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_133),
.A2(n_136),
.B(n_145),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_151),
.B1(n_104),
.B2(n_119),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_0),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_150),
.Y(n_169)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_149),
.Y(n_163)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_0),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_89),
.A2(n_111),
.B1(n_121),
.B2(n_114),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_100),
.B1(n_114),
.B2(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_4),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_107),
.B1(n_93),
.B2(n_87),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_191),
.B1(n_153),
.B2(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_161),
.B(n_170),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_92),
.B(n_127),
.Y(n_162)
);

XOR2x1_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_150),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_164),
.B(n_142),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_178),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_173),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_167),
.A2(n_182),
.B1(n_7),
.B2(n_9),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_99),
.B1(n_93),
.B2(n_118),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_174),
.B(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_172),
.B(n_175),
.Y(n_220)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_96),
.B(n_115),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_112),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_108),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_88),
.B1(n_107),
.B2(n_91),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_101),
.B1(n_94),
.B2(n_6),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_131),
.B1(n_138),
.B2(n_132),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_193),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_198),
.A2(n_169),
.B(n_164),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_216),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_217),
.B(n_177),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_154),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_207),
.C(n_213),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_142),
.C(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_208),
.B(n_218),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_186),
.B1(n_178),
.B2(n_173),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_190),
.B1(n_183),
.B2(n_181),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_192),
.B1(n_176),
.B2(n_191),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_130),
.C(n_5),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_182),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_185),
.B(n_163),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_169),
.B(n_4),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_15),
.C(n_11),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_6),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_241)
);

XOR2x1_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_245),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_197),
.Y(n_273)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_230),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_242),
.C(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_241),
.B1(n_250),
.B2(n_251),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_169),
.B(n_162),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_240),
.B(n_214),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_166),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_7),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_194),
.A2(n_11),
.B(n_13),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_221),
.B(n_219),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_14),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_14),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_14),
.B1(n_200),
.B2(n_194),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_200),
.A2(n_196),
.B1(n_198),
.B2(n_210),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_231),
.B1(n_250),
.B2(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_263),
.C(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_227),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_216),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_207),
.C(n_199),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_224),
.C(n_225),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_232),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_226),
.C(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_252),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_280),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_255),
.A2(n_235),
.B1(n_251),
.B2(n_231),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_287),
.B1(n_253),
.B2(n_271),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_259),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_242),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_288),
.C(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_212),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_234),
.B1(n_209),
.B2(n_223),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_244),
.C(n_245),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_258),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_216),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_272),
.C(n_256),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_257),
.B1(n_271),
.B2(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_262),
.B(n_260),
.C(n_269),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_294),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_259),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_274),
.C(n_277),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_305),
.C(n_274),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_297),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_275),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_285),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_258),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_298),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_300),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_322),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_321),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_299),
.B(n_279),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_264),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_313),
.B(n_288),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_329),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_305),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_318),
.A2(n_293),
.B1(n_313),
.B2(n_311),
.Y(n_329)
);

XOR2x2_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_319),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_332),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_330),
.B(n_317),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_334),
.A2(n_331),
.B(n_329),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_335),
.B1(n_328),
.B2(n_331),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_294),
.C(n_327),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_294),
.Y(n_340)
);


endmodule