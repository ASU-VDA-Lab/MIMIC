module fake_netlist_5_149_n_626 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_626);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_626;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_611;
wire n_444;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_280;
wire n_590;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_77),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_24),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

BUFx2_ASAP7_75t_SL g140 ( 
.A(n_75),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_67),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_26),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_12),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_20),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_22),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_110),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_61),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_80),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_44),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_38),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_21),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_46),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_49),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_4),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

INVxp33_ASAP7_75t_SL g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

BUFx8_ASAP7_75t_SL g171 ( 
.A(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_27),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_39),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_91),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_51),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_10),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_71),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_70),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_0),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_14),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_69),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_13),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_74),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_54),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_11),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_48),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_18),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_47),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_137),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_145),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g216 ( 
.A(n_165),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g217 ( 
.A(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_151),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_146),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_148),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_153),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_156),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_138),
.B(n_2),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_157),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_159),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_162),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_R g248 ( 
.A(n_154),
.B(n_15),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_175),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_182),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_184),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_138),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_214),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_150),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_160),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_161),
.Y(n_269)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_152),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_161),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_140),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_150),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_189),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_192),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_248),
.B(n_192),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_211),
.B(n_172),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_217),
.B(n_152),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_204),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_227),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_233),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_205),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_281),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_194),
.B1(n_197),
.B2(n_202),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_185),
.B1(n_203),
.B2(n_201),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_164),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_253),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_198),
.Y(n_309)
);

BUFx6f_ASAP7_75t_SL g310 ( 
.A(n_302),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_263),
.A2(n_180),
.B(n_200),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_251),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_252),
.B(n_251),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_166),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_173),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

BUFx4f_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

AND3x4_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_2),
.C(n_3),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_263),
.Y(n_327)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_195),
.B1(n_193),
.B2(n_187),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_181),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_281),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_274),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_16),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_287),
.B(n_6),
.Y(n_345)
);

NAND2xp33_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_276),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_6),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_268),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_268),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_267),
.B(n_269),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_267),
.B(n_19),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_290),
.B(n_7),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_254),
.Y(n_353)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_289),
.B(n_7),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_270),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_278),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_269),
.B(n_8),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_260),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_294),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

OR2x6_ASAP7_75t_SL g369 ( 
.A(n_304),
.B(n_295),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_301),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_353),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_326),
.A2(n_300),
.B1(n_299),
.B2(n_298),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_300),
.B1(n_299),
.B2(n_298),
.Y(n_375)
);

BUFx6f_ASAP7_75t_SL g376 ( 
.A(n_358),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_257),
.B1(n_279),
.B2(n_283),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_272),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_301),
.Y(n_379)
);

AO22x2_ASAP7_75t_L g380 ( 
.A1(n_311),
.A2(n_290),
.B1(n_303),
.B2(n_296),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_327),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_309),
.A2(n_296),
.B1(n_272),
.B2(n_288),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_288),
.Y(n_383)
);

NAND2x1p5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_260),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_321),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_319),
.B(n_293),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

AO22x2_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

AO22x2_ASAP7_75t_L g402 ( 
.A1(n_365),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

AO22x2_ASAP7_75t_L g404 ( 
.A1(n_306),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_315),
.A2(n_270),
.B1(n_30),
.B2(n_31),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_270),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

NAND2x1p5_ASAP7_75t_L g411 ( 
.A(n_324),
.B(n_29),
.Y(n_411)
);

OAI221xp5_ASAP7_75t_L g412 ( 
.A1(n_345),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.C(n_35),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_330),
.B(n_307),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_367),
.Y(n_414)
);

OAI221xp5_ASAP7_75t_L g415 ( 
.A1(n_347),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.C(n_41),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_334),
.B(n_42),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_336),
.B(n_322),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_322),
.B(n_43),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_318),
.B(n_45),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_342),
.B(n_50),
.Y(n_424)
);

AO22x2_ASAP7_75t_L g425 ( 
.A1(n_329),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_358),
.Y(n_426)
);

OR2x6_ASAP7_75t_L g427 ( 
.A(n_354),
.B(n_56),
.Y(n_427)
);

OAI221xp5_ASAP7_75t_L g428 ( 
.A1(n_356),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.C(n_65),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_310),
.Y(n_430)
);

NAND2x1p5_ASAP7_75t_L g431 ( 
.A(n_325),
.B(n_68),
.Y(n_431)
);

OAI221xp5_ASAP7_75t_L g432 ( 
.A1(n_314),
.A2(n_357),
.B1(n_325),
.B2(n_359),
.C(n_368),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_SL g433 ( 
.A(n_376),
.B(n_359),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_413),
.B(n_367),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_357),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_421),
.B(n_368),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g437 ( 
.A(n_426),
.B(n_344),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_378),
.B(n_305),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_379),
.B(n_362),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_370),
.B(n_410),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_414),
.B(n_344),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_377),
.B(n_362),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_392),
.B(n_362),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_386),
.B(n_360),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_374),
.B(n_360),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_385),
.B(n_360),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_387),
.B(n_328),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_388),
.B(n_344),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_389),
.B(n_328),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_390),
.B(n_393),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_417),
.B(n_73),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_409),
.B(n_79),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_370),
.B(n_83),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_419),
.B(n_84),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_394),
.B(n_85),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_396),
.B(n_86),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_397),
.B(n_88),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_430),
.B(n_89),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_370),
.B(n_90),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_384),
.B(n_92),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_398),
.B(n_94),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_429),
.B(n_95),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_399),
.B(n_96),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_423),
.B(n_100),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g465 ( 
.A(n_400),
.B(n_101),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_383),
.B(n_103),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_371),
.B(n_104),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_373),
.B(n_108),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_383),
.B(n_111),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_112),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_403),
.B(n_113),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_418),
.B(n_114),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_408),
.B(n_416),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_436),
.A2(n_432),
.B(n_420),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_380),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_438),
.A2(n_462),
.B(n_471),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

AO31x2_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_422),
.A3(n_391),
.B(n_406),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_462),
.A2(n_412),
.B(n_401),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_434),
.B(n_380),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_382),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g483 ( 
.A1(n_451),
.A2(n_375),
.B(n_372),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_411),
.B(n_431),
.Y(n_485)
);

O2A1O1Ixp5_ASAP7_75t_SL g486 ( 
.A1(n_443),
.A2(n_382),
.B(n_428),
.C(n_415),
.Y(n_486)
);

A2O1A1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_454),
.A2(n_405),
.B(n_407),
.C(n_375),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_442),
.A2(n_427),
.B1(n_369),
.B2(n_402),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_466),
.A2(n_404),
.B(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_437),
.B(n_427),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_459),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_R g495 ( 
.A(n_469),
.B(n_470),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_425),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_395),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_447),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_467),
.A2(n_424),
.B(n_116),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_476),
.A2(n_456),
.B(n_455),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_449),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_478),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

OAI221xp5_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_458),
.B1(n_465),
.B2(n_441),
.C(n_457),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

O2A1O1Ixp33_ASAP7_75t_L g508 ( 
.A1(n_481),
.A2(n_463),
.B(n_461),
.C(n_452),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_501),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

OAI21x1_ASAP7_75t_SL g511 ( 
.A1(n_482),
.A2(n_468),
.B(n_395),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_500),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_115),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_L g516 ( 
.A1(n_497),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_123),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_474),
.A2(n_124),
.B(n_125),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_492),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_126),
.B(n_127),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_480),
.A2(n_128),
.B(n_129),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_483),
.A2(n_132),
.B(n_135),
.C(n_490),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_479),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_486),
.A2(n_493),
.B(n_499),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_494),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_479),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_495),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_505),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_514),
.B(n_487),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_515),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_512),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_526),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_515),
.A2(n_523),
.B(n_522),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_512),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_524),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_520),
.A2(n_518),
.B(n_521),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_513),
.B(n_519),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_507),
.B(n_525),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_525),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_525),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_509),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_512),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_503),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_517),
.Y(n_549)
);

OAI21x1_ASAP7_75t_SL g550 ( 
.A1(n_508),
.A2(n_511),
.B(n_502),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_522),
.B(n_503),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_509),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_510),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_520),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_547),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_502),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_548),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_538),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_530),
.B(n_521),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_506),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_R g562 ( 
.A(n_531),
.B(n_551),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_534),
.B(n_516),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_R g564 ( 
.A(n_531),
.B(n_518),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_R g565 ( 
.A(n_551),
.B(n_539),
.Y(n_565)
);

CKINVDCx8_ASAP7_75t_R g566 ( 
.A(n_541),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_R g567 ( 
.A(n_527),
.B(n_549),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_529),
.B(n_552),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_R g569 ( 
.A(n_549),
.B(n_536),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_554),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_560),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_570),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_557),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_528),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_556),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_568),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_555),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_555),
.B(n_532),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_541),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_559),
.B(n_541),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_566),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_556),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_528),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_571),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_571),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_575),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_573),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_576),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_580),
.B(n_536),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_574),
.B(n_563),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_587),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_587),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_584),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_573),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_577),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_589),
.B(n_578),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_586),
.B(n_578),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_595),
.B(n_562),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_597),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_588),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_596),
.Y(n_601)
);

AO221x2_ASAP7_75t_L g602 ( 
.A1(n_592),
.A2(n_590),
.B1(n_581),
.B2(n_582),
.C(n_567),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_598),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_600),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_599),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_601),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_602),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_597),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_604),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_591),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_609),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_608),
.Y(n_612)
);

INVx5_ASAP7_75t_SL g613 ( 
.A(n_612),
.Y(n_613)
);

NAND4xp25_ASAP7_75t_L g614 ( 
.A(n_613),
.B(n_611),
.C(n_603),
.D(n_610),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_605),
.Y(n_615)
);

NAND4xp75_ASAP7_75t_L g616 ( 
.A(n_615),
.B(n_608),
.C(n_606),
.D(n_533),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_586),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_617),
.B(n_592),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_619),
.B(n_575),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_620),
.A2(n_575),
.B1(n_547),
.B2(n_546),
.Y(n_621)
);

OAI322xp33_ASAP7_75t_L g622 ( 
.A1(n_621),
.A2(n_533),
.A3(n_594),
.B1(n_575),
.B2(n_565),
.C1(n_569),
.C2(n_564),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_622),
.A2(n_546),
.B1(n_554),
.B2(n_537),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_623),
.Y(n_624)
);

OAI221xp5_ASAP7_75t_R g625 ( 
.A1(n_624),
.A2(n_550),
.B1(n_579),
.B2(n_537),
.C(n_540),
.Y(n_625)
);

AOI211xp5_ASAP7_75t_L g626 ( 
.A1(n_625),
.A2(n_537),
.B(n_540),
.C(n_535),
.Y(n_626)
);


endmodule