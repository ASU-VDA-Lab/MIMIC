module fake_jpeg_126_n_93 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_13),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_28),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_29),
.B1(n_27),
.B2(n_35),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_48),
.B1(n_29),
.B2(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_51),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_0),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_14),
.B(n_22),
.C(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g60 ( 
.A(n_54),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_47),
.C(n_45),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_64),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_8),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_70),
.B(n_3),
.C(n_4),
.D(n_7),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_53),
.B1(n_45),
.B2(n_5),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_45),
.B(n_4),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_71),
.C(n_76),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_67),
.B1(n_61),
.B2(n_6),
.C(n_7),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_81),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_8),
.B1(n_9),
.B2(n_15),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_9),
.B1(n_16),
.B2(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_73),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_84),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_82),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_77),
.B(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_18),
.B(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_73),
.Y(n_93)
);


endmodule