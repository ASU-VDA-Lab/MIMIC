module fake_netlist_1_5880_n_813 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_114, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_813);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_813;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_729;
wire n_519;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g115 ( .A(n_65), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_10), .B(n_110), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_45), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_13), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_31), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_75), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_18), .Y(n_121) );
BUFx10_ASAP7_75t_L g122 ( .A(n_55), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_47), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_18), .Y(n_124) );
BUFx10_ASAP7_75t_L g125 ( .A(n_5), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_20), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_17), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_90), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_100), .Y(n_130) );
INVxp33_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_76), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_101), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_52), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_46), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_22), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_74), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_6), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_4), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_68), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_23), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_25), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_35), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_114), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_113), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_103), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_0), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_32), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_57), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_70), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_30), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_16), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_109), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_37), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_24), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_50), .Y(n_162) );
AOI22x1_ASAP7_75t_SL g163 ( .A1(n_124), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_140), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_121), .B(n_3), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
AOI22x1_ASAP7_75t_SL g167 ( .A1(n_124), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_117), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_138), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
XNOR2xp5_ASAP7_75t_L g171 ( .A(n_126), .B(n_7), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_139), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_147), .B(n_8), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_122), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_115), .Y(n_175) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_141), .A2(n_58), .B(n_108), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
NOR2x1_ASAP7_75t_L g178 ( .A(n_144), .B(n_9), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_130), .B(n_10), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_157), .B(n_11), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_115), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_132), .B(n_11), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_174), .B(n_122), .Y(n_185) );
CKINVDCx6p67_ASAP7_75t_R g186 ( .A(n_181), .Y(n_186) );
INVxp33_ASAP7_75t_L g187 ( .A(n_181), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_175), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_174), .B(n_137), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_168), .B(n_141), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_175), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_168), .B(n_151), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_170), .B(n_151), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_170), .B(n_152), .C(n_155), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_184), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_174), .B(n_122), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_184), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_174), .B(n_119), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_184), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_173), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_183), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_177), .B(n_154), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_166), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_183), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_183), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_173), .B(n_119), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_173), .B(n_120), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_177), .B(n_154), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_173), .B(n_120), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_190), .B(n_182), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_204), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_204), .B(n_169), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_204), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_185), .B(n_182), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_188), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_208), .A2(n_179), .B1(n_158), .B2(n_129), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_201), .A2(n_158), .B1(n_129), .B2(n_136), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_190), .B(n_180), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_204), .B(n_123), .Y(n_228) );
BUFx8_ASAP7_75t_L g229 ( .A(n_186), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_214), .B(n_123), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_215), .B(n_145), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_188), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_217), .B(n_145), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_187), .B(n_125), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_208), .B(n_146), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_192), .A2(n_136), .B1(n_172), .B2(n_164), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_186), .B(n_171), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_202), .B(n_131), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_205), .B(n_146), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_211), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_192), .B(n_159), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_211), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_201), .A2(n_178), .B1(n_118), .B2(n_143), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g245 ( .A(n_200), .B(n_150), .C(n_178), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_196), .B(n_159), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_203), .B(n_199), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_199), .B(n_160), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_193), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_203), .B(n_160), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_216), .B(n_125), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_206), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_193), .B(n_166), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_206), .B(n_133), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_195), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_195), .B(n_149), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_207), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_200), .A2(n_163), .B1(n_167), .B2(n_125), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_198), .B(n_153), .Y(n_260) );
NAND3x1_ASAP7_75t_L g261 ( .A(n_198), .B(n_163), .C(n_167), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_248), .A2(n_216), .B(n_210), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_229), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_252), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_221), .A2(n_176), .B(n_161), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_221), .A2(n_176), .B(n_162), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_262), .B(n_171), .Y(n_268) );
NOR2x1_ASAP7_75t_R g269 ( .A(n_229), .B(n_156), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_224), .A2(n_176), .B(n_161), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_256), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_253), .A2(n_176), .B(n_162), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_253), .A2(n_213), .B(n_212), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_250), .B(n_116), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_224), .A2(n_213), .B(n_212), .Y(n_275) );
AO21x1_ASAP7_75t_L g276 ( .A1(n_247), .A2(n_213), .B(n_212), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_250), .B(n_143), .Y(n_277) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_259), .B(n_209), .C(n_197), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_256), .B(n_219), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_SL g280 ( .A1(n_218), .A2(n_209), .B(n_197), .C(n_194), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_252), .B(n_143), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_227), .B(n_143), .Y(n_282) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_235), .A2(n_132), .B(n_142), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
OR2x6_ASAP7_75t_L g285 ( .A(n_226), .B(n_142), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_219), .B(n_115), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_220), .B(n_12), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_257), .B(n_12), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_235), .B(n_13), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_237), .A2(n_115), .B1(n_135), .B2(n_183), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_232), .A2(n_209), .B(n_189), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_238), .B(n_14), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_232), .A2(n_197), .B(n_194), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_234), .A2(n_194), .B(n_191), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_238), .B(n_225), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_234), .A2(n_191), .B(n_189), .Y(n_298) );
NOR2x1p5_ASAP7_75t_SL g299 ( .A(n_243), .B(n_189), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_241), .A2(n_135), .B(n_183), .C(n_207), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_249), .B(n_14), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_228), .B(n_135), .Y(n_302) );
OAI21x1_ASAP7_75t_SL g303 ( .A1(n_276), .A2(n_243), .B(n_251), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_284), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_265), .B(n_241), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_268), .B(n_260), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_274), .B(n_242), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_290), .B(n_223), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_263), .A2(n_245), .B(n_239), .C(n_222), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_271), .B(n_244), .Y(n_311) );
INVx5_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
AOI21x1_ASAP7_75t_SL g313 ( .A1(n_289), .A2(n_246), .B(n_230), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_264), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_296), .B(n_231), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_272), .A2(n_236), .B(n_255), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_293), .B(n_233), .Y(n_319) );
AND2x6_ASAP7_75t_L g320 ( .A(n_297), .B(n_229), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_267), .A2(n_258), .B(n_191), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_267), .A2(n_240), .B(n_258), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_277), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_266), .A2(n_207), .B(n_261), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_285), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
AO21x1_ASAP7_75t_L g327 ( .A1(n_270), .A2(n_135), .B(n_261), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_285), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_285), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_275), .A2(n_207), .B(n_63), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_288), .B(n_15), .Y(n_331) );
INVx3_ASAP7_75t_SL g332 ( .A(n_288), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_321), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_322), .A2(n_280), .B(n_302), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_317), .B(n_283), .Y(n_335) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_327), .A2(n_278), .B(n_301), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_320), .Y(n_337) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_324), .A2(n_300), .B(n_282), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_324), .B(n_299), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_329), .A2(n_281), .B1(n_269), .B2(n_291), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_321), .A2(n_298), .B(n_295), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_316), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_304), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_307), .B(n_279), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_307), .B(n_292), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_298), .B(n_295), .Y(n_349) );
OA21x2_ASAP7_75t_L g350 ( .A1(n_303), .A2(n_294), .B(n_275), .Y(n_350) );
BUFx2_ASAP7_75t_R g351 ( .A(n_325), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_325), .A2(n_286), .B1(n_294), .B2(n_273), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_318), .A2(n_62), .B(n_107), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_306), .B(n_19), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_332), .B(n_19), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_306), .B(n_20), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_342), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_342), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_342), .B(n_332), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_341), .A2(n_330), .B(n_303), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_357), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_343), .B(n_347), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_333), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_344), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_351), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_348), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_333), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_337), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_337), .A2(n_320), .B1(n_328), .B2(n_314), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_355), .Y(n_378) );
NOR2x1_ASAP7_75t_R g379 ( .A(n_337), .B(n_314), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_335), .A2(n_319), .B(n_331), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_333), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_357), .B(n_332), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_366), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_367), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_364), .B(n_339), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_367), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_379), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_387), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_375), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_373), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_364), .B(n_339), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_383), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_383), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_369), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_363), .A2(n_356), .B1(n_354), .B2(n_357), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_380), .B(n_349), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_380), .B(n_349), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_362), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_368), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_382), .B(n_349), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_382), .B(n_349), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_371), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_372), .B(n_356), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_358), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_384), .B(n_349), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_386), .B(n_351), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_384), .B(n_349), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_359), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_359), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_385), .B(n_336), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_365), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_372), .B(n_354), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_374), .B(n_356), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_365), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_374), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_361), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_360), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_387), .B(n_336), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_375), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_361), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_389), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_389), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_392), .B(n_376), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_390), .B(n_378), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_390), .B(n_378), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_430), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_391), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_403), .B(n_360), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_388), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_391), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_408), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_403), .A2(n_386), .B1(n_340), .B2(n_335), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_408), .B(n_336), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_390), .B(n_336), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_399), .B(n_336), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_426), .B(n_347), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_426), .B(n_347), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_399), .B(n_350), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_432), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_426), .B(n_381), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_413), .B(n_346), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_397), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_432), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_432), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_399), .B(n_404), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_428), .B(n_350), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_395), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_397), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_428), .B(n_350), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_404), .B(n_350), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_429), .B(n_350), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_402), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_404), .B(n_350), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_402), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_405), .B(n_338), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_405), .B(n_338), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_406), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_392), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_388), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_429), .B(n_346), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_406), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_413), .B(n_346), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_407), .Y(n_479) );
NOR2xp33_ASAP7_75t_SL g480 ( .A(n_409), .B(n_320), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_395), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_433), .B(n_338), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_431), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_398), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_405), .B(n_338), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_407), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_410), .B(n_338), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_412), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_433), .B(n_338), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_410), .B(n_341), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_388), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_412), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_393), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_414), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_414), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_425), .B(n_340), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_415), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_393), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_425), .B(n_320), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_393), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_435), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_415), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_400), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_400), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_400), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_398), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_416), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_416), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_401), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_463), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_461), .B(n_394), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_456), .B(n_410), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_437), .B(n_411), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_461), .B(n_394), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_455), .B(n_411), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_438), .B(n_411), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_440), .B(n_418), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_440), .B(n_418), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_463), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_455), .B(n_421), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_438), .B(n_418), .Y(n_523) );
NAND2xp33_ASAP7_75t_L g524 ( .A(n_448), .B(n_320), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_459), .B(n_421), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_460), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_443), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_441), .B(n_420), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_441), .B(n_420), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_459), .B(n_422), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_460), .B(n_420), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_460), .B(n_435), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_443), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_446), .B(n_423), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_454), .B(n_396), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_454), .B(n_396), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_446), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_502), .B(n_396), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_490), .B(n_434), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_434), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_439), .A2(n_496), .B1(n_444), .B2(n_478), .C(n_457), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_476), .B(n_422), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_476), .B(n_427), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_447), .B(n_427), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_458), .B(n_464), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_474), .B(n_417), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_466), .B(n_434), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_447), .B(n_417), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_464), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_468), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_468), .Y(n_552) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_484), .B(n_419), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_470), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_474), .B(n_417), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_484), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_470), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_466), .B(n_423), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_469), .B(n_423), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_473), .B(n_425), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_473), .B(n_431), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_481), .B(n_424), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_477), .B(n_431), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_477), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
AND2x4_ASAP7_75t_SL g566 ( .A(n_480), .B(n_424), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_474), .B(n_424), .Y(n_567) );
OR2x6_ASAP7_75t_L g568 ( .A(n_462), .B(n_401), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_452), .B(n_401), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_436), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_450), .B(n_451), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_462), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_479), .Y(n_573) );
OAI32xp33_ASAP7_75t_L g574 ( .A1(n_465), .A2(n_430), .A3(n_308), .B1(n_323), .B2(n_320), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_450), .B(n_436), .Y(n_575) );
INVxp33_ASAP7_75t_L g576 ( .A(n_465), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_483), .Y(n_577) );
AND2x6_ASAP7_75t_SL g578 ( .A(n_500), .B(n_320), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_479), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_483), .B(n_430), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_486), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_488), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_488), .Y(n_584) );
BUFx2_ASAP7_75t_L g585 ( .A(n_467), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_492), .Y(n_586) );
OAI32xp33_ASAP7_75t_L g587 ( .A1(n_467), .A2(n_308), .A3(n_323), .B1(n_326), .B2(n_311), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_492), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_451), .B(n_453), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_494), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_445), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_483), .B(n_312), .Y(n_592) );
AND2x4_ASAP7_75t_SL g593 ( .A(n_508), .B(n_315), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_508), .B(n_21), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_509), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_471), .B(n_21), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_445), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_475), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_509), .B(n_22), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_572), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_524), .A2(n_353), .B(n_449), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_565), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_538), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_568), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_585), .B(n_449), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_572), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_513), .B(n_482), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_568), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_558), .B(n_471), .Y(n_610) );
OR2x6_ASAP7_75t_L g611 ( .A(n_526), .B(n_482), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_545), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_513), .B(n_489), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_589), .B(n_472), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_595), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_571), .B(n_472), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_516), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_512), .B(n_489), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_527), .Y(n_621) );
NOR2xp33_ASAP7_75t_R g622 ( .A(n_524), .B(n_23), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_533), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_541), .A2(n_487), .A3(n_485), .B1(n_499), .B2(n_503), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_541), .B(n_485), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_576), .A2(n_499), .B1(n_497), .B2(n_503), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_562), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_522), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_537), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_559), .B(n_487), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_519), .B(n_494), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_520), .B(n_497), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_546), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_528), .B(n_495), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_550), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_551), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_525), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_517), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_556), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_515), .B(n_499), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_529), .B(n_495), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_548), .B(n_475), .Y(n_643) );
OR2x6_ASAP7_75t_L g644 ( .A(n_526), .B(n_491), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_535), .B(n_491), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_592), .B(n_312), .Y(n_646) );
CKINVDCx16_ASAP7_75t_R g647 ( .A(n_596), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_552), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_539), .B(n_493), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_554), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_557), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_536), .B(n_493), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_517), .B(n_442), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_540), .B(n_498), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_514), .B(n_498), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_514), .B(n_501), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_553), .B(n_501), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_518), .B(n_504), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_530), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_564), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_532), .B(n_442), .Y(n_661) );
BUFx3_ASAP7_75t_L g662 ( .A(n_566), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_577), .B(n_442), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_531), .B(n_504), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_573), .Y(n_665) );
INVx3_ASAP7_75t_SL g666 ( .A(n_553), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_518), .B(n_505), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_570), .B(n_575), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_523), .B(n_505), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_544), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_523), .B(n_506), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_569), .B(n_506), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_579), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_578), .B(n_510), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_576), .B(n_510), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_534), .B(n_442), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g677 ( .A(n_594), .B(n_353), .C(n_334), .D(n_352), .Y(n_677) );
NAND2x1p5_ASAP7_75t_L g678 ( .A(n_592), .B(n_312), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_581), .Y(n_679) );
OR2x6_ASAP7_75t_L g680 ( .A(n_547), .B(n_330), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_625), .A2(n_534), .B1(n_511), .B2(n_560), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_602), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_639), .B(n_511), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_607), .B(n_549), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g685 ( .A1(n_666), .A2(n_547), .B(n_555), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_624), .B(n_521), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_644), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_662), .B(n_555), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_647), .A2(n_599), .B1(n_542), .B2(n_543), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_657), .A2(n_560), .B1(n_583), .B2(n_582), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_612), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_613), .Y(n_692) );
OAI322xp33_ASAP7_75t_L g693 ( .A1(n_670), .A2(n_588), .A3(n_584), .B1(n_590), .B2(n_586), .C1(n_563), .C2(n_561), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_623), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_614), .B(n_597), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_623), .Y(n_696) );
OAI22xp5_ASAP7_75t_SL g697 ( .A1(n_644), .A2(n_567), .B1(n_577), .B2(n_597), .Y(n_697) );
NAND2xp33_ASAP7_75t_L g698 ( .A(n_622), .B(n_561), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_604), .B(n_567), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_677), .B(n_574), .C(n_587), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_638), .Y(n_701) );
INVxp33_ASAP7_75t_L g702 ( .A(n_674), .Y(n_702) );
NOR2xp33_ASAP7_75t_SL g703 ( .A(n_611), .B(n_580), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_629), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_629), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_633), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_601), .A2(n_608), .B1(n_609), .B2(n_611), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_600), .B(n_563), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_626), .B(n_580), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_640), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_680), .A2(n_598), .B1(n_591), .B2(n_312), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_633), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_603), .B(n_593), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_600), .B(n_334), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_635), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_606), .B(n_617), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_610), .B(n_341), .Y(n_717) );
INVxp67_ASAP7_75t_L g718 ( .A(n_616), .Y(n_718) );
INVx1_ASAP7_75t_SL g719 ( .A(n_661), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_631), .B(n_312), .Y(n_720) );
OAI32xp33_ASAP7_75t_L g721 ( .A1(n_632), .A2(n_326), .A3(n_352), .B1(n_309), .B2(n_313), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_668), .B(n_312), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_635), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_646), .A2(n_310), .B(n_27), .Y(n_724) );
OAI32xp33_ASAP7_75t_L g725 ( .A1(n_634), .A2(n_26), .A3(n_28), .B1(n_29), .B2(n_33), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_636), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_636), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_630), .B(n_315), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_653), .A2(n_315), .B(n_36), .C(n_38), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_641), .B(n_34), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_648), .Y(n_731) );
INVx1_ASAP7_75t_SL g732 ( .A(n_661), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_648), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_606), .B(n_39), .Y(n_734) );
NAND2x1_ASAP7_75t_L g735 ( .A(n_653), .B(n_315), .Y(n_735) );
AOI321xp33_ASAP7_75t_L g736 ( .A1(n_689), .A2(n_605), .A3(n_675), .B1(n_637), .B2(n_659), .C(n_628), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_701), .Y(n_737) );
AOI31xp33_ASAP7_75t_L g738 ( .A1(n_688), .A2(n_678), .A3(n_620), .B(n_642), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_694), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_696), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_684), .B(n_627), .Y(n_741) );
OAI31xp33_ASAP7_75t_L g742 ( .A1(n_689), .A2(n_663), .A3(n_676), .B(n_650), .Y(n_742) );
OAI322xp33_ASAP7_75t_SL g743 ( .A1(n_686), .A2(n_618), .A3(n_615), .B1(n_643), .B2(n_649), .C1(n_655), .C2(n_669), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_704), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_735), .B(n_663), .Y(n_745) );
OA21x2_ASAP7_75t_SL g746 ( .A1(n_702), .A2(n_667), .B(n_654), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_718), .B(n_656), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_685), .B(n_672), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_693), .A2(n_660), .B1(n_651), .B2(n_619), .C(n_621), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_707), .B(n_679), .C(n_673), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_700), .A2(n_680), .B1(n_645), .B2(n_652), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_705), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_698), .A2(n_665), .B(n_673), .Y(n_753) );
NAND2x1_ASAP7_75t_L g754 ( .A(n_687), .B(n_664), .Y(n_754) );
INVx2_ASAP7_75t_SL g755 ( .A(n_710), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_706), .Y(n_756) );
OA21x2_ASAP7_75t_SL g757 ( .A1(n_719), .A2(n_671), .B(n_658), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_681), .B(n_679), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_703), .A2(n_315), .B1(n_41), .B2(n_42), .Y(n_759) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_734), .A2(n_40), .B(n_43), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_691), .B(n_44), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_695), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_712), .Y(n_763) );
AOI222xp33_ASAP7_75t_L g764 ( .A1(n_682), .A2(n_48), .B1(n_49), .B2(n_51), .C1(n_53), .C2(n_54), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_715), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_722), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_736), .B(n_709), .C(n_714), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_743), .A2(n_692), .B1(n_708), .B2(n_683), .C(n_732), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g769 ( .A1(n_738), .A2(n_729), .B(n_703), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_754), .A2(n_719), .B1(n_732), .B2(n_697), .Y(n_770) );
AOI22x1_ASAP7_75t_L g771 ( .A1(n_757), .A2(n_730), .B1(n_724), .B2(n_699), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_749), .B(n_690), .Y(n_772) );
OAI221xp5_ASAP7_75t_SL g773 ( .A1(n_742), .A2(n_713), .B1(n_711), .B2(n_720), .C(n_717), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_748), .A2(n_725), .B(n_716), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_751), .A2(n_733), .B1(n_731), .B2(n_723), .C(n_727), .Y(n_775) );
AOI21xp33_ASAP7_75t_SL g776 ( .A1(n_746), .A2(n_724), .B(n_721), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_737), .A2(n_726), .B(n_699), .C(n_728), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_753), .A2(n_56), .B(n_59), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_755), .A2(n_60), .B1(n_61), .B2(n_64), .Y(n_779) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_750), .A2(n_66), .B1(n_67), .B2(n_69), .C(n_71), .Y(n_780) );
OAI211xp5_ASAP7_75t_L g781 ( .A1(n_759), .A2(n_72), .B(n_73), .C(n_77), .Y(n_781) );
AOI322xp5_ASAP7_75t_L g782 ( .A1(n_747), .A2(n_80), .A3(n_82), .B1(n_83), .B2(n_84), .C1(n_85), .C2(n_86), .Y(n_782) );
AOI211x1_ASAP7_75t_L g783 ( .A1(n_758), .A2(n_739), .B(n_765), .C(n_763), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_770), .Y(n_784) );
NAND4xp25_ASAP7_75t_L g785 ( .A(n_769), .B(n_764), .C(n_760), .D(n_758), .Y(n_785) );
OAI211xp5_ASAP7_75t_SL g786 ( .A1(n_772), .A2(n_760), .B(n_761), .C(n_766), .Y(n_786) );
NOR3xp33_ASAP7_75t_L g787 ( .A(n_776), .B(n_761), .C(n_740), .Y(n_787) );
NOR3xp33_ASAP7_75t_L g788 ( .A(n_780), .B(n_756), .C(n_752), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_771), .A2(n_745), .B1(n_762), .B2(n_744), .C(n_741), .Y(n_789) );
OAI21xp33_ASAP7_75t_L g790 ( .A1(n_771), .A2(n_745), .B(n_89), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_774), .B(n_88), .Y(n_791) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_773), .B(n_91), .C(n_92), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_787), .B(n_783), .C(n_767), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_784), .B(n_768), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_788), .B(n_777), .Y(n_795) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_791), .B(n_781), .Y(n_796) );
NOR2x1_ASAP7_75t_L g797 ( .A(n_785), .B(n_779), .Y(n_797) );
OR2x6_ASAP7_75t_L g798 ( .A(n_797), .B(n_790), .Y(n_798) );
NAND2xp5_ASAP7_75t_SL g799 ( .A(n_794), .B(n_792), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_795), .B(n_778), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_798), .B(n_796), .Y(n_801) );
NAND2xp5_ASAP7_75t_SL g802 ( .A(n_799), .B(n_793), .Y(n_802) );
AO22x1_ASAP7_75t_L g803 ( .A1(n_801), .A2(n_800), .B1(n_789), .B2(n_786), .Y(n_803) );
BUFx2_ASAP7_75t_L g804 ( .A(n_802), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_804), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_803), .Y(n_806) );
AOI22x1_ASAP7_75t_L g807 ( .A1(n_806), .A2(n_782), .B1(n_775), .B2(n_96), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_805), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_808), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_809), .B(n_807), .Y(n_810) );
OAI21x1_ASAP7_75t_L g811 ( .A1(n_810), .A2(n_93), .B(n_94), .Y(n_811) );
OA22x2_ASAP7_75t_L g812 ( .A1(n_811), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_812), .A2(n_102), .B1(n_104), .B2(n_112), .Y(n_813) );
endmodule