module fake_netlist_6_3778_n_1827 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1827);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1827;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_SL g197 ( 
.A(n_60),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_93),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_37),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_18),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_196),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_77),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_95),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_23),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_146),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_62),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_23),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_38),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_122),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_57),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_182),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_27),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_46),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_103),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_195),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_76),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_26),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_74),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_84),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_35),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_87),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_133),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_111),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_89),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_154),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_25),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_33),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_123),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_193),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_110),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_2),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_96),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_156),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_71),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_56),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_29),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_69),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_140),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_24),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_38),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_131),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_91),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_166),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_10),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_136),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_150),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_142),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_40),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_165),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_152),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_27),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_97),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_47),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_88),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_41),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_2),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_1),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_162),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_190),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_189),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_11),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_178),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_132),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_86),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_44),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_167),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_81),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_4),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_7),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_28),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_113),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_73),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_117),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_181),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_109),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_36),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_41),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_54),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_20),
.Y(n_321)
);

BUFx8_ASAP7_75t_SL g322 ( 
.A(n_183),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_120),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_31),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_9),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_90),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_6),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_100),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_99),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_39),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_49),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_164),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_65),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_20),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_66),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_115),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_68),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_138),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_7),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_10),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_61),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_151),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_54),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_17),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_126),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_116),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_21),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_31),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_141),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_168),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_135),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_188),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_44),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_118),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_102),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_159),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_128),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_169),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_6),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_80),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_1),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_15),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_149),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_47),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_114),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_134),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_3),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_127),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_170),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_32),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_36),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_40),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_106),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_171),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_45),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_57),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_52),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_79),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_174),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_185),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_175),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_14),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_160),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_52),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_75),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_34),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_78),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_29),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_137),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_17),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_51),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_72),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_22),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_8),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_215),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_294),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_294),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_252),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_230),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_294),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_246),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_259),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_294),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_283),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_255),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_322),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_294),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_296),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_294),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_294),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_221),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_248),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_248),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_202),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_294),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_284),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_311),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_303),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_303),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_221),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_341),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_272),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_272),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_201),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_222),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_272),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_328),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_272),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_236),
.Y(n_429)
);

INVx4_ASAP7_75t_R g430 ( 
.A(n_265),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_272),
.Y(n_431)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_198),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_388),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_248),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_237),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_200),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_203),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_226),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_222),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_265),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_238),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_282),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_330),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_270),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_275),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_240),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_223),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_249),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_262),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_282),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_276),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_279),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_223),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_384),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_227),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_227),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_281),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_299),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_310),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_264),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_320),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_324),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_293),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_340),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_353),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_361),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_266),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_229),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_386),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_229),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_293),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_262),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_359),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_301),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_301),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_271),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_326),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_326),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_350),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g490 ( 
.A(n_359),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_280),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_350),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_362),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_199),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_206),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_286),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_207),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_211),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_434),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_498),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_424),
.B(n_197),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_197),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_397),
.A2(n_268),
.B(n_251),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_495),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_431),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_338),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_338),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_403),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

BUFx8_ASAP7_75t_L g520 ( 
.A(n_487),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_398),
.A2(n_371),
.B1(n_391),
.B2(n_390),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_410),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_351),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_455),
.A2(n_268),
.B(n_251),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_455),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_432),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_395),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_351),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_432),
.Y(n_538)
);

AND3x2_ASAP7_75t_L g539 ( 
.A(n_412),
.B(n_377),
.C(n_285),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_429),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_395),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_489),
.B(n_356),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_444),
.B(n_377),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_448),
.B(n_314),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_439),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_432),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_456),
.B(n_356),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_414),
.B(n_362),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_457),
.B(n_274),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_401),
.B(n_314),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_458),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_469),
.B(n_484),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_420),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_463),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_414),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_492),
.B(n_314),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_418),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_467),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_470),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_445),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_398),
.A2(n_292),
.B1(n_334),
.B2(n_390),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_419),
.B(n_204),
.Y(n_570)
);

BUFx8_ASAP7_75t_L g571 ( 
.A(n_436),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_399),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_482),
.B(n_329),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_471),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_406),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_427),
.B(n_204),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_452),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_500),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_574),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_533),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_499),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_517),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_454),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_510),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_517),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_574),
.B(n_421),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_556),
.B(n_506),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_512),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_572),
.B(n_446),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_572),
.B(n_460),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_544),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_466),
.C(n_454),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_500),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_501),
.B(n_462),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_503),
.B(n_411),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_512),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_518),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_500),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_549),
.A2(n_408),
.B1(n_405),
.B2(n_411),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_572),
.B(n_466),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

INVxp67_ASAP7_75t_R g607 ( 
.A(n_559),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_557),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_SL g609 ( 
.A(n_544),
.B(n_364),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_536),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_517),
.Y(n_611)
);

OAI221xp5_ASAP7_75t_L g612 ( 
.A1(n_514),
.A2(n_474),
.B1(n_481),
.B2(n_478),
.C(n_475),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_561),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_525),
.Y(n_614)
);

AOI21x1_ASAP7_75t_L g615 ( 
.A1(n_527),
.A2(n_505),
.B(n_525),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_512),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_506),
.B(n_476),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_548),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_562),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_543),
.B(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_562),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_500),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_541),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_562),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_549),
.A2(n_408),
.B1(n_453),
.B2(n_443),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_517),
.Y(n_627)
);

INVxp33_ASAP7_75t_SL g628 ( 
.A(n_579),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_572),
.B(n_486),
.Y(n_629)
);

BUFx4f_ASAP7_75t_L g630 ( 
.A(n_517),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_486),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_507),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_531),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_536),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_573),
.Y(n_635)
);

AND2x2_ASAP7_75t_SL g636 ( 
.A(n_504),
.B(n_274),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_560),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_531),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_501),
.B(n_413),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_508),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_511),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_504),
.B(n_491),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_511),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_R g644 ( 
.A(n_577),
.B(n_491),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_560),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_522),
.A2(n_289),
.B1(n_297),
.B2(n_298),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_571),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_543),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_504),
.A2(n_552),
.B1(n_505),
.B2(n_524),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_502),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_513),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_535),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_540),
.B(n_443),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_513),
.Y(n_654)
);

AND3x2_ASAP7_75t_L g655 ( 
.A(n_504),
.B(n_316),
.C(n_285),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_535),
.Y(n_656)
);

AND3x2_ASAP7_75t_L g657 ( 
.A(n_524),
.B(n_317),
.C(n_316),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_537),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_522),
.A2(n_453),
.B1(n_490),
.B2(n_496),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_551),
.B(n_317),
.Y(n_660)
);

AND2x6_ASAP7_75t_L g661 ( 
.A(n_538),
.B(n_333),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_547),
.B(n_496),
.Y(n_662)
);

INVx8_ASAP7_75t_L g663 ( 
.A(n_552),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_552),
.B(n_333),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_502),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_537),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_568),
.B(n_490),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_570),
.B(n_472),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_536),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_570),
.B(n_553),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_515),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_546),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_515),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_569),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_526),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_564),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_526),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_564),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_575),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_575),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_538),
.B(n_260),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_502),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_502),
.B(n_242),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_519),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_519),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g686 ( 
.A1(n_527),
.A2(n_214),
.B(n_212),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_519),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_524),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_519),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_516),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_521),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_521),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_563),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_552),
.A2(n_313),
.B1(n_213),
.B2(n_233),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_521),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_571),
.B(n_329),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_571),
.Y(n_699)
);

CKINVDCx16_ASAP7_75t_R g700 ( 
.A(n_569),
.Y(n_700)
);

INVxp67_ASAP7_75t_SL g701 ( 
.A(n_538),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_563),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_538),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_521),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_521),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_521),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_509),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_523),
.Y(n_708)
);

AND3x2_ASAP7_75t_L g709 ( 
.A(n_555),
.B(n_224),
.C(n_219),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_523),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_571),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_523),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_523),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_523),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_523),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_527),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_552),
.A2(n_315),
.B1(n_244),
.B2(n_263),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_536),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_534),
.B(n_459),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_520),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_636),
.B(n_566),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_639),
.B(n_534),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_633),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_649),
.B(n_250),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_636),
.B(n_260),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_707),
.B(n_459),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_602),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_592),
.B(n_566),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_688),
.B(n_566),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_668),
.B(n_461),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_596),
.B(n_520),
.Y(n_731)
);

INVx8_ASAP7_75t_L g732 ( 
.A(n_663),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_638),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_652),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_620),
.B(n_461),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_639),
.B(n_477),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_688),
.B(n_566),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_656),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_596),
.B(n_520),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_674),
.A2(n_505),
.B1(n_527),
.B2(n_336),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_670),
.A2(n_477),
.B1(n_479),
.B2(n_493),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_637),
.B(n_567),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_586),
.B(n_479),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_637),
.B(n_520),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_648),
.B(n_205),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_689),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_648),
.B(n_567),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_620),
.B(n_483),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_701),
.B(n_567),
.Y(n_749)
);

INVx8_ASAP7_75t_L g750 ( 
.A(n_663),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_582),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_658),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_703),
.B(n_567),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_690),
.B(n_576),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_581),
.Y(n_755)
);

BUFx5_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_581),
.B(n_600),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_692),
.A2(n_576),
.B(n_542),
.C(n_514),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_619),
.B(n_555),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_666),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_645),
.B(n_483),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_588),
.B(n_576),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_590),
.B(n_576),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_689),
.B(n_505),
.Y(n_764)
);

BUFx6f_ASAP7_75t_SL g765 ( 
.A(n_660),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_645),
.B(n_205),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_593),
.B(n_536),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_631),
.B(n_208),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_663),
.B(n_509),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_601),
.B(n_536),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_663),
.B(n_542),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_616),
.B(n_660),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_716),
.B(n_545),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_719),
.B(n_613),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_599),
.B(n_493),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_716),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_604),
.B(n_208),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_599),
.B(n_209),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_642),
.B(n_545),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_621),
.B(n_545),
.Y(n_780)
);

O2A1O1Ixp5_ASAP7_75t_L g781 ( 
.A1(n_615),
.A2(n_565),
.B(n_558),
.C(n_555),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_624),
.B(n_545),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_608),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_625),
.B(n_209),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_682),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_661),
.B(n_253),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_582),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_674),
.A2(n_336),
.B1(n_380),
.B2(n_260),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_661),
.A2(n_380),
.B1(n_336),
.B2(n_277),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_692),
.B(n_336),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_597),
.B(n_558),
.Y(n_791)
);

INVx6_ASAP7_75t_L g792 ( 
.A(n_664),
.Y(n_792)
);

BUFx6f_ASAP7_75t_SL g793 ( 
.A(n_672),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_694),
.B(n_336),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_694),
.A2(n_323),
.B(n_241),
.C(n_243),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_617),
.B(n_545),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_683),
.A2(n_530),
.B(n_528),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_676),
.B(n_678),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_679),
.B(n_545),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_661),
.A2(n_380),
.B1(n_269),
.B2(n_306),
.Y(n_800)
);

AND2x6_ASAP7_75t_SL g801 ( 
.A(n_653),
.B(n_239),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_609),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_607),
.B(n_558),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_680),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_609),
.A2(n_295),
.B1(n_254),
.B2(n_256),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_682),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_695),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_528),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_702),
.B(n_530),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_684),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_684),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_700),
.A2(n_364),
.B1(n_367),
.B2(n_370),
.Y(n_812)
);

NOR2x1p5_ASAP7_75t_L g813 ( 
.A(n_720),
.B(n_367),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_685),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_650),
.B(n_532),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_591),
.B(n_210),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_650),
.B(n_532),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_659),
.B(n_210),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_605),
.B(n_216),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_685),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_583),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_629),
.B(n_216),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_583),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_665),
.B(n_532),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_607),
.B(n_565),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_646),
.B(n_217),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_632),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_717),
.A2(n_291),
.B1(n_305),
.B2(n_304),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_665),
.B(n_554),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_664),
.B(n_245),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_696),
.A2(n_290),
.B1(n_261),
.B2(n_273),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_594),
.A2(n_300),
.B1(n_288),
.B2(n_309),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_687),
.B(n_554),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_687),
.B(n_554),
.Y(n_834)
);

OAI221xp5_ASAP7_75t_L g835 ( 
.A1(n_612),
.A2(n_308),
.B1(n_302),
.B2(n_278),
.C(n_267),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_595),
.B(n_217),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_662),
.B(n_667),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_644),
.B(n_218),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_640),
.B(n_548),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_641),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_643),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_643),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_661),
.A2(n_380),
.B1(n_258),
.B2(n_257),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_651),
.B(n_548),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_623),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_720),
.B(n_628),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_651),
.B(n_548),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_SL g848 ( 
.A1(n_623),
.A2(n_402),
.B1(n_404),
.B2(n_416),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_698),
.B(n_218),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_654),
.B(n_548),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_654),
.B(n_247),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_628),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_664),
.B(n_539),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_618),
.B(n_337),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_587),
.Y(n_855)
);

AND3x1_ASAP7_75t_L g856 ( 
.A(n_671),
.B(n_358),
.C(n_373),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_671),
.B(n_357),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_673),
.B(n_319),
.C(n_318),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_673),
.B(n_360),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_675),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_675),
.Y(n_861)
);

NAND2x1_ASAP7_75t_L g862 ( 
.A(n_661),
.B(n_430),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_677),
.B(n_384),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_677),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_691),
.B(n_380),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_584),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_584),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_614),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_691),
.B(n_363),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_693),
.B(n_704),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_693),
.B(n_704),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_614),
.A2(n_712),
.B(n_715),
.C(n_706),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_776),
.B(n_705),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_776),
.B(n_705),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_746),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_730),
.B(n_399),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_807),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_774),
.B(n_402),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_722),
.B(n_647),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_728),
.B(n_706),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_755),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_732),
.B(n_664),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_852),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_755),
.B(n_647),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_732),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_848),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_788),
.B(n_740),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_759),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_730),
.B(n_404),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_757),
.B(n_416),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_759),
.Y(n_891)
);

CKINVDCx11_ASAP7_75t_R g892 ( 
.A(n_801),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_853),
.B(n_723),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_783),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_785),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_827),
.Y(n_896)
);

AND2x2_ASAP7_75t_SL g897 ( 
.A(n_826),
.B(n_788),
.Y(n_897)
);

NOR3x1_ASAP7_75t_L g898 ( 
.A(n_818),
.B(n_389),
.C(n_368),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_785),
.Y(n_899)
);

BUFx4f_ASAP7_75t_L g900 ( 
.A(n_792),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_751),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_740),
.B(n_757),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_726),
.B(n_417),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_787),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_842),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_845),
.Y(n_906)
);

AND2x4_ASAP7_75t_SL g907 ( 
.A(n_769),
.B(n_635),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_842),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_840),
.B(n_708),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_806),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_732),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_853),
.B(n_655),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_726),
.B(n_417),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_761),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_733),
.B(n_657),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_741),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_743),
.B(n_449),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_743),
.B(n_449),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_724),
.B(n_699),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_803),
.B(n_699),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_840),
.B(n_708),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_750),
.B(n_635),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_736),
.B(n_711),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_810),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_793),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_735),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_811),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_736),
.B(n_711),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_750),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_748),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_864),
.B(n_710),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_864),
.B(n_779),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_837),
.A2(n_779),
.B1(n_791),
.B2(n_772),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_775),
.B(n_802),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_814),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_820),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_750),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_813),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_825),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_747),
.B(n_796),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_796),
.B(n_710),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_837),
.A2(n_714),
.B1(n_713),
.B2(n_718),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_863),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_734),
.B(n_738),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_792),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_819),
.B(n_822),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_841),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_866),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_752),
.B(n_712),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_754),
.B(n_758),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_742),
.B(n_715),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_721),
.B(n_627),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_802),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_861),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_821),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_830),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_792),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_823),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_769),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_819),
.B(n_822),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_775),
.B(n_585),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_855),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_760),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_773),
.B(n_627),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_749),
.B(n_627),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_778),
.B(n_370),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_727),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_769),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_830),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_765),
.B(n_615),
.Y(n_971)
);

AND2x2_ASAP7_75t_SL g972 ( 
.A(n_826),
.B(n_392),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_816),
.B(n_371),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_753),
.B(n_804),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_828),
.B(n_287),
.C(n_228),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_765),
.B(n_686),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_798),
.B(n_697),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_729),
.B(n_697),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_766),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_836),
.B(n_589),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_867),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_816),
.B(n_836),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_868),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_830),
.B(n_622),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_745),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_849),
.B(n_589),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_856),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_725),
.A2(n_697),
.B1(n_681),
.B2(n_622),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_771),
.Y(n_989)
);

OR2x6_ASAP7_75t_SL g990 ( 
.A(n_858),
.B(n_391),
.Y(n_990)
);

INVx5_ASAP7_75t_L g991 ( 
.A(n_771),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_781),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_771),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_737),
.B(n_808),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_768),
.B(n_307),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_764),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_764),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_809),
.B(n_815),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_817),
.B(n_626),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_851),
.Y(n_1000)
);

AOI211xp5_ASAP7_75t_L g1001 ( 
.A1(n_812),
.A2(n_348),
.B(n_312),
.C(n_321),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_824),
.B(n_626),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_829),
.B(n_580),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_833),
.B(n_580),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_838),
.B(n_325),
.Y(n_1005)
);

AO22x1_ASAP7_75t_L g1006 ( 
.A1(n_812),
.A2(n_327),
.B1(n_331),
.B2(n_339),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_762),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_725),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_834),
.B(n_580),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_831),
.Y(n_1010)
);

INVxp33_ASAP7_75t_L g1011 ( 
.A(n_777),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_846),
.B(n_585),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_857),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_784),
.B(n_343),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_805),
.B(n_630),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_793),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_763),
.B(n_598),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_862),
.B(n_585),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_799),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_832),
.B(n_630),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_756),
.B(n_789),
.Y(n_1021)
);

BUFx4f_ASAP7_75t_L g1022 ( 
.A(n_854),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_870),
.B(n_598),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_767),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_731),
.B(n_344),
.Y(n_1026)
);

OR2x2_ASAP7_75t_SL g1027 ( 
.A(n_739),
.B(n_329),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_744),
.B(n_598),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_786),
.A2(n_611),
.B1(n_606),
.B2(n_603),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_795),
.A2(n_781),
.B(n_835),
.C(n_872),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_770),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_859),
.A2(n_681),
.B1(n_606),
.B2(n_603),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_797),
.B(n_611),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_780),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_869),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_782),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_871),
.B(n_611),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_789),
.B(n_871),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_756),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_839),
.B(n_220),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_756),
.B(n_618),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_844),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_847),
.B(n_220),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_850),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_982),
.B(n_756),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_964),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_893),
.B(n_790),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1039),
.A2(n_618),
.B(n_843),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1039),
.A2(n_618),
.B(n_843),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_902),
.B(n_800),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_934),
.B(n_347),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1039),
.A2(n_756),
.B(n_634),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1039),
.A2(n_634),
.B(n_669),
.Y(n_1053)
);

OR2x6_ASAP7_75t_SL g1054 ( 
.A(n_883),
.B(n_376),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_972),
.B(n_382),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_901),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_1035),
.B(n_225),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_887),
.A2(n_961),
.B1(n_1008),
.B2(n_933),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_904),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_958),
.B(n_794),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_980),
.A2(n_887),
.B(n_986),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_SL g1062 ( 
.A(n_885),
.B(n_225),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1008),
.A2(n_865),
.B(n_374),
.C(n_369),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_1016),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_906),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_890),
.B(n_394),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_875),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_907),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1021),
.A2(n_610),
.B(n_669),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_939),
.B(n_529),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_943),
.A2(n_973),
.B(n_962),
.C(n_917),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_939),
.B(n_681),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_881),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_1018),
.A2(n_669),
.B(n_634),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_881),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_918),
.A2(n_365),
.B(n_231),
.C(n_232),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_885),
.Y(n_1077)
);

BUFx10_ASAP7_75t_L g1078 ( 
.A(n_928),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_876),
.B(n_228),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_938),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_888),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_900),
.B(n_231),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_975),
.A2(n_709),
.B(n_3),
.C(n_4),
.Y(n_1083)
);

AO32x2_ASAP7_75t_L g1084 ( 
.A1(n_979),
.A2(n_0),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_998),
.A2(n_669),
.B(n_634),
.Y(n_1085)
);

NAND3xp33_ASAP7_75t_SL g1086 ( 
.A(n_889),
.B(n_232),
.C(n_234),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_891),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_894),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_932),
.A2(n_610),
.B1(n_634),
.B2(n_669),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_900),
.B(n_234),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_926),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_998),
.A2(n_610),
.B(n_550),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_1001),
.B(n_366),
.C(n_365),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_949),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_932),
.B(n_287),
.Y(n_1095)
);

BUFx8_ASAP7_75t_L g1096 ( 
.A(n_930),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_894),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_944),
.B(n_366),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_891),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_935),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_885),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_926),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_954),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_922),
.B(n_610),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_913),
.B(n_369),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_903),
.B(n_374),
.C(n_332),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1010),
.A2(n_378),
.B(n_342),
.C(n_387),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_940),
.A2(n_610),
.B(n_550),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_985),
.B(n_355),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_923),
.B(n_335),
.C(n_345),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_974),
.A2(n_379),
.B(n_385),
.C(n_383),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_1040),
.A2(n_346),
.B(n_354),
.C(n_352),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_974),
.A2(n_349),
.B1(n_550),
.B2(n_64),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_985),
.B(n_550),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1036),
.B(n_5),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_922),
.B(n_67),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_951),
.A2(n_550),
.B1(n_63),
.B2(n_70),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_975),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1118)
);

OAI22x1_ASAP7_75t_L g1119 ( 
.A1(n_886),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_954),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_879),
.A2(n_21),
.B(n_22),
.C(n_30),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_877),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_951),
.A2(n_33),
.B(n_34),
.C(n_39),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_935),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_878),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_994),
.A2(n_94),
.B(n_191),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_911),
.B(n_92),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_911),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_914),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_1011),
.A2(n_1014),
.B(n_967),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1005),
.B(n_42),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1018),
.A2(n_85),
.B(n_186),
.Y(n_1132)
);

NOR2x1_ASAP7_75t_L g1133 ( 
.A(n_884),
.B(n_83),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_911),
.Y(n_1134)
);

AO32x1_ASAP7_75t_L g1135 ( 
.A1(n_992),
.A2(n_42),
.A3(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_929),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_920),
.A2(n_43),
.B(n_48),
.C(n_49),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_873),
.A2(n_112),
.B1(n_184),
.B2(n_172),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1000),
.B(n_48),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_929),
.B(n_937),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_925),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_893),
.B(n_105),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_922),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_968),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1013),
.B(n_50),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1007),
.B(n_50),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_990),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_874),
.A2(n_98),
.B(n_157),
.Y(n_1148)
);

CKINVDCx11_ASAP7_75t_R g1149 ( 
.A(n_892),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1019),
.B(n_51),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_874),
.A2(n_82),
.B(n_124),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1038),
.A2(n_977),
.B1(n_953),
.B2(n_1015),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_977),
.A2(n_145),
.B1(n_194),
.B2(n_55),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_929),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1026),
.A2(n_58),
.B(n_989),
.C(n_947),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_996),
.A2(n_58),
.B1(n_997),
.B2(n_882),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_916),
.B(n_995),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1024),
.B(n_1016),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_937),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_1043),
.A2(n_1030),
.B(n_1037),
.C(n_941),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_996),
.A2(n_997),
.B1(n_882),
.B2(n_1034),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1030),
.A2(n_1025),
.B(n_1042),
.C(n_948),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_R g1163 ( 
.A(n_937),
.B(n_945),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_957),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_941),
.A2(n_1033),
.B(n_965),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_971),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_981),
.A2(n_983),
.B(n_1028),
.C(n_950),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_945),
.B(n_912),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_909),
.B(n_921),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_909),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_1020),
.A2(n_880),
.B(n_952),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_921),
.B(n_931),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_950),
.A2(n_963),
.B1(n_956),
.B2(n_959),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_996),
.A2(n_997),
.B1(n_882),
.B2(n_942),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1031),
.B(n_880),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_970),
.Y(n_1176)
);

INVx3_ASAP7_75t_SL g1177 ( 
.A(n_912),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_987),
.B(n_1027),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1031),
.B(n_965),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_993),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1046),
.Y(n_1181)
);

AOI211x1_ASAP7_75t_L g1182 ( 
.A1(n_1058),
.A2(n_1006),
.B(n_896),
.C(n_908),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1049),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1055),
.A2(n_915),
.B1(n_919),
.B2(n_993),
.C(n_960),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1051),
.A2(n_1071),
.B(n_1050),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1157),
.B(n_945),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1079),
.A2(n_991),
.B1(n_1028),
.B2(n_915),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1125),
.B(n_898),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1171),
.A2(n_1061),
.A3(n_1152),
.B(n_1162),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1091),
.B(n_984),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_1056),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1066),
.B(n_969),
.C(n_960),
.Y(n_1192)
);

AO22x1_ASAP7_75t_L g1193 ( 
.A1(n_1105),
.A2(n_991),
.B1(n_969),
.B2(n_960),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1089),
.A2(n_1033),
.A3(n_966),
.B(n_978),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1101),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1155),
.A2(n_1113),
.B(n_1093),
.C(n_1130),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1074),
.A2(n_978),
.B(n_1023),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1085),
.A2(n_966),
.B(n_1017),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1094),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1122),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1101),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1048),
.A2(n_1002),
.B(n_999),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1052),
.A2(n_1023),
.B(n_1017),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1170),
.B(n_955),
.Y(n_1204)
);

AOI211x1_ASAP7_75t_L g1205 ( 
.A1(n_1146),
.A2(n_1009),
.B(n_1004),
.C(n_1003),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1088),
.B(n_976),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1053),
.A2(n_1009),
.B(n_1029),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1169),
.A2(n_1022),
.B(n_1041),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1167),
.A2(n_905),
.B(n_895),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1168),
.B(n_993),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1132),
.A2(n_955),
.B(n_899),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1102),
.B(n_984),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1113),
.A2(n_910),
.B(n_924),
.C(n_927),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1108),
.A2(n_988),
.B(n_1032),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1095),
.B(n_1044),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1045),
.A2(n_936),
.B(n_1044),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1172),
.A2(n_1044),
.B(n_1012),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1073),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1092),
.A2(n_969),
.B(n_1179),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1168),
.B(n_1134),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1174),
.A2(n_1161),
.B(n_1117),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1131),
.B(n_1070),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1139),
.B(n_1145),
.Y(n_1223)
);

AO21x1_ASAP7_75t_L g1224 ( 
.A1(n_1153),
.A2(n_1138),
.B(n_1126),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1116),
.B(n_1104),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1150),
.B(n_1115),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1078),
.B(n_1103),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1065),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1166),
.B(n_1097),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1101),
.Y(n_1230)
);

NOR3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1178),
.B(n_1086),
.C(n_1110),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1123),
.A2(n_1063),
.A3(n_1111),
.B(n_1148),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1151),
.A2(n_1060),
.B(n_1173),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_SL g1234 ( 
.A1(n_1107),
.A2(n_1112),
.B(n_1142),
.C(n_1076),
.Y(n_1234)
);

AO22x2_ASAP7_75t_L g1235 ( 
.A1(n_1093),
.A2(n_1156),
.B1(n_1084),
.B2(n_1147),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1059),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1173),
.A2(n_1072),
.B(n_1114),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1144),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1096),
.Y(n_1239)
);

AOI21xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1119),
.A2(n_1098),
.B(n_1057),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1100),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1096),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1078),
.B(n_1081),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1047),
.B(n_1104),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1121),
.A2(n_1137),
.B(n_1083),
.C(n_1118),
.Y(n_1245)
);

O2A1O1Ixp5_ASAP7_75t_L g1246 ( 
.A1(n_1082),
.A2(n_1090),
.B(n_1062),
.C(n_1047),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1087),
.A2(n_1099),
.B(n_1124),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1075),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1133),
.A2(n_1127),
.B(n_1120),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1134),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1116),
.B(n_1104),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1077),
.A2(n_1136),
.B1(n_1116),
.B2(n_1129),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1077),
.A2(n_1136),
.B(n_1135),
.Y(n_1253)
);

OAI22x1_ASAP7_75t_L g1254 ( 
.A1(n_1176),
.A2(n_1177),
.B1(n_1136),
.B2(n_1077),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1128),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1140),
.A2(n_1180),
.B(n_1163),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1135),
.A2(n_1106),
.B(n_1158),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1135),
.A2(n_1158),
.B(n_1159),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_SL g1259 ( 
.A1(n_1084),
.A2(n_1180),
.B(n_1143),
.Y(n_1259)
);

CKINVDCx6p67_ASAP7_75t_R g1260 ( 
.A(n_1064),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1068),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1128),
.A2(n_1159),
.B(n_1154),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1084),
.Y(n_1263)
);

AND2x2_ASAP7_75t_SL g1264 ( 
.A(n_1128),
.B(n_1159),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1141),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1154),
.A2(n_1164),
.B(n_1080),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1054),
.A2(n_1152),
.B(n_1165),
.Y(n_1267)
);

NAND2xp33_ASAP7_75t_L g1268 ( 
.A(n_1149),
.B(n_982),
.Y(n_1268)
);

BUFx12f_ASAP7_75t_L g1269 ( 
.A(n_1080),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1067),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1074),
.A2(n_1069),
.B(n_1165),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1055),
.A2(n_897),
.B1(n_972),
.B2(n_982),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1125),
.B(n_926),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1051),
.B(n_982),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1051),
.B(n_982),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1066),
.B(n_730),
.C(n_982),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1046),
.Y(n_1277)
);

NAND3x1_ASAP7_75t_L g1278 ( 
.A(n_1055),
.B(n_730),
.C(n_876),
.Y(n_1278)
);

NOR2x1_ASAP7_75t_L g1279 ( 
.A(n_1175),
.B(n_1179),
.Y(n_1279)
);

O2A1O1Ixp5_ASAP7_75t_SL g1280 ( 
.A1(n_1058),
.A2(n_946),
.B(n_961),
.C(n_980),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1073),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1055),
.A2(n_730),
.B(n_982),
.Y(n_1282)
);

CKINVDCx8_ASAP7_75t_R g1283 ( 
.A(n_1056),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1074),
.A2(n_1069),
.B(n_1165),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1046),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1046),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1055),
.A2(n_982),
.B(n_730),
.C(n_961),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1073),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1116),
.B(n_732),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1171),
.A2(n_1061),
.A3(n_1152),
.B(n_1165),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1157),
.B(n_774),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1051),
.B(n_982),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1071),
.B(n_972),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1152),
.A2(n_1165),
.B(n_1058),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1168),
.B(n_893),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1055),
.A2(n_982),
.B(n_730),
.C(n_961),
.Y(n_1296)
);

INVx5_ASAP7_75t_L g1297 ( 
.A(n_1101),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1055),
.A2(n_982),
.B(n_730),
.C(n_961),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1051),
.B(n_982),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1171),
.A2(n_1061),
.A3(n_1152),
.B(n_1165),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1171),
.A2(n_1061),
.A3(n_1152),
.B(n_1165),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1071),
.A2(n_897),
.B1(n_972),
.B2(n_982),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1071),
.B(n_972),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1101),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1051),
.B(n_982),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1066),
.B(n_730),
.C(n_982),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1066),
.B(n_730),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1165),
.A2(n_1039),
.B(n_776),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1171),
.A2(n_1061),
.A3(n_1152),
.B(n_1165),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1051),
.B(n_982),
.Y(n_1310)
);

AO32x2_ASAP7_75t_L g1311 ( 
.A1(n_1058),
.A2(n_1152),
.A3(n_1174),
.B1(n_1156),
.B2(n_828),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1074),
.A2(n_1069),
.B(n_1165),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1051),
.B(n_982),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1051),
.B(n_982),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1185),
.B(n_1302),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1211),
.A2(n_1284),
.B(n_1271),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1276),
.C(n_1306),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1272),
.A2(n_1306),
.B1(n_1276),
.B2(n_1278),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1280),
.A2(n_1296),
.B(n_1287),
.Y(n_1319)
);

NAND2x1_ASAP7_75t_L g1320 ( 
.A(n_1221),
.B(n_1270),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1298),
.A2(n_1294),
.B(n_1293),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1225),
.B(n_1251),
.Y(n_1322)
);

CKINVDCx8_ASAP7_75t_R g1323 ( 
.A(n_1236),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1227),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1264),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1303),
.A2(n_1272),
.B(n_1267),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1283),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1282),
.A2(n_1196),
.B(n_1267),
.C(n_1310),
.Y(n_1328)
);

INVx6_ASAP7_75t_L g1329 ( 
.A(n_1191),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1291),
.A2(n_1314),
.B1(n_1299),
.B2(n_1305),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1261),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1312),
.A2(n_1207),
.B(n_1203),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1274),
.A2(n_1313),
.B1(n_1292),
.B2(n_1275),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1191),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1220),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1225),
.B(n_1251),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1244),
.A2(n_1258),
.B(n_1253),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1197),
.A2(n_1202),
.B(n_1308),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1199),
.Y(n_1339)
);

BUFx8_ASAP7_75t_SL g1340 ( 
.A(n_1269),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1200),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1279),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1217),
.A2(n_1245),
.B(n_1214),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1233),
.A2(n_1219),
.B(n_1216),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1239),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1231),
.A2(n_1226),
.B(n_1240),
.C(n_1246),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1240),
.A2(n_1223),
.B(n_1257),
.C(n_1222),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1247),
.A2(n_1198),
.B(n_1208),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1225),
.A2(n_1251),
.B1(n_1289),
.B2(n_1273),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1213),
.A2(n_1249),
.B(n_1215),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1192),
.A2(n_1234),
.B(n_1237),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1212),
.B(n_1190),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1235),
.A2(n_1188),
.B1(n_1259),
.B2(n_1187),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1237),
.A2(n_1270),
.B(n_1192),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1209),
.A2(n_1263),
.B(n_1204),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1266),
.A2(n_1262),
.B(n_1277),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1218),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1289),
.B(n_1193),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1285),
.A2(n_1286),
.B(n_1238),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1252),
.A2(n_1206),
.B(n_1281),
.C(n_1288),
.Y(n_1360)
);

AOI221xp5_ASAP7_75t_L g1361 ( 
.A1(n_1235),
.A2(n_1184),
.B1(n_1248),
.B2(n_1205),
.C(n_1268),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1241),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1243),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1289),
.A2(n_1194),
.B(n_1311),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1250),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1186),
.B(n_1229),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1256),
.A2(n_1250),
.B(n_1255),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1297),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1210),
.A2(n_1265),
.B(n_1311),
.C(n_1295),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1297),
.Y(n_1370)
);

OR2x6_ASAP7_75t_L g1371 ( 
.A(n_1182),
.B(n_1254),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1194),
.A2(n_1311),
.B(n_1309),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1265),
.B(n_1295),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1242),
.A2(n_1232),
.B(n_1189),
.C(n_1300),
.Y(n_1374)
);

AOI31xp33_ASAP7_75t_L g1375 ( 
.A1(n_1232),
.A2(n_1189),
.A3(n_1260),
.B(n_1290),
.Y(n_1375)
);

AOI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_1290),
.B(n_1301),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1195),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1189),
.B(n_1300),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1201),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1201),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1230),
.B(n_1304),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1267),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1307),
.A2(n_876),
.B1(n_889),
.B2(n_1278),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1185),
.B(n_897),
.Y(n_1384)
);

INVx4_ASAP7_75t_SL g1385 ( 
.A(n_1225),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1192),
.B(n_1056),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1306),
.C(n_1276),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1261),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1306),
.C(n_1276),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1181),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1307),
.B(n_1282),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1228),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1211),
.A2(n_1284),
.B(n_1271),
.Y(n_1396)
);

AOI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1307),
.A2(n_730),
.B1(n_1282),
.B2(n_876),
.C(n_889),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1181),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1211),
.A2(n_1284),
.B(n_1271),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1211),
.A2(n_1284),
.B(n_1271),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1185),
.A2(n_1280),
.B(n_961),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1211),
.A2(n_1284),
.B(n_1271),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1244),
.A2(n_1267),
.B(n_1258),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1211),
.A2(n_1284),
.B(n_1271),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1307),
.A2(n_897),
.B1(n_788),
.B2(n_972),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1185),
.A2(n_1280),
.B(n_961),
.Y(n_1407)
);

OAI211xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_730),
.C(n_1287),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1225),
.B(n_1251),
.Y(n_1409)
);

AO21x1_ASAP7_75t_L g1410 ( 
.A1(n_1293),
.A2(n_1303),
.B(n_1302),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1224),
.A2(n_1183),
.A3(n_1171),
.B(n_1061),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1224),
.A2(n_1183),
.A3(n_1171),
.B(n_1061),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1264),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1228),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1224),
.A2(n_1183),
.A3(n_1171),
.B(n_1061),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1307),
.A2(n_730),
.B1(n_1282),
.B2(n_876),
.C(n_889),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1185),
.B(n_897),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1181),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1306),
.C(n_1276),
.Y(n_1420)
);

AOI21xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1307),
.A2(n_730),
.B(n_876),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1228),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1185),
.A2(n_1280),
.B(n_961),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1306),
.C(n_1276),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1185),
.A2(n_1280),
.B(n_961),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1297),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1220),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1273),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1307),
.A2(n_972),
.B1(n_876),
.B2(n_889),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1181),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1307),
.A2(n_1272),
.B1(n_1282),
.B2(n_1276),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1185),
.A2(n_1280),
.B(n_961),
.Y(n_1433)
);

O2A1O1Ixp5_ASAP7_75t_L g1434 ( 
.A1(n_1321),
.A2(n_1319),
.B(n_1423),
.C(n_1425),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1421),
.B(n_1394),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1363),
.B(n_1330),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1384),
.B(n_1418),
.Y(n_1437)
);

CKINVDCx6p67_ASAP7_75t_R g1438 ( 
.A(n_1327),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1323),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1329),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1324),
.B(n_1429),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1351),
.A2(n_1319),
.B(n_1401),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1340),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1389),
.A2(n_1390),
.B1(n_1392),
.B2(n_1428),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1341),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1357),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1429),
.B(n_1418),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1346),
.A2(n_1417),
.B(n_1397),
.C(n_1391),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1397),
.A2(n_1417),
.B(n_1387),
.C(n_1420),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1317),
.A2(n_1424),
.B(n_1408),
.C(n_1406),
.Y(n_1450)
);

NOR2xp67_ASAP7_75t_L g1451 ( 
.A(n_1334),
.B(n_1373),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1403),
.A2(n_1430),
.B1(n_1412),
.B2(n_1406),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1383),
.A2(n_1333),
.B1(n_1315),
.B2(n_1328),
.Y(n_1453)
);

INVx3_ASAP7_75t_SL g1454 ( 
.A(n_1331),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1351),
.A2(n_1407),
.B(n_1401),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1369),
.A2(n_1432),
.B1(n_1321),
.B2(n_1318),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1326),
.A2(n_1408),
.B(n_1343),
.C(n_1318),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1329),
.Y(n_1458)
);

NOR2x1_ASAP7_75t_SL g1459 ( 
.A(n_1358),
.B(n_1322),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1388),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1358),
.B(n_1336),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1342),
.B(n_1415),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1347),
.A2(n_1433),
.B(n_1425),
.C(n_1423),
.Y(n_1463)
);

OA22x2_ASAP7_75t_L g1464 ( 
.A1(n_1336),
.A2(n_1409),
.B1(n_1371),
.B2(n_1382),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1369),
.A2(n_1353),
.B1(n_1409),
.B2(n_1343),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1342),
.B(n_1407),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1422),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1433),
.A2(n_1320),
.B(n_1364),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1409),
.A2(n_1361),
.B1(n_1414),
.B2(n_1325),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1410),
.B(n_1361),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1364),
.B(n_1374),
.Y(n_1471)
);

OA22x2_ASAP7_75t_L g1472 ( 
.A1(n_1371),
.A2(n_1358),
.B1(n_1404),
.B2(n_1370),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1360),
.A2(n_1375),
.B(n_1374),
.C(n_1350),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1395),
.Y(n_1474)
);

O2A1O1Ixp5_ASAP7_75t_L g1475 ( 
.A1(n_1350),
.A2(n_1376),
.B(n_1349),
.C(n_1378),
.Y(n_1475)
);

AOI211xp5_ASAP7_75t_L g1476 ( 
.A1(n_1386),
.A2(n_1360),
.B(n_1372),
.C(n_1431),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1325),
.A2(n_1414),
.B1(n_1393),
.B2(n_1339),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1375),
.A2(n_1371),
.B(n_1337),
.C(n_1398),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1372),
.B(n_1355),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1377),
.Y(n_1480)
);

OAI31xp33_ASAP7_75t_L g1481 ( 
.A1(n_1419),
.A2(n_1370),
.A3(n_1362),
.B(n_1427),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1345),
.B(n_1335),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1348),
.A2(n_1338),
.B(n_1332),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1316),
.A2(n_1402),
.B(n_1405),
.Y(n_1484)
);

AO21x1_ASAP7_75t_L g1485 ( 
.A1(n_1356),
.A2(n_1354),
.B(n_1368),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1411),
.B(n_1416),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1411),
.B(n_1413),
.Y(n_1487)
);

O2A1O1Ixp5_ASAP7_75t_L g1488 ( 
.A1(n_1368),
.A2(n_1365),
.B(n_1380),
.C(n_1379),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1367),
.B(n_1381),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1426),
.B(n_1344),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1396),
.A2(n_1399),
.B(n_1400),
.Y(n_1491)
);

A2O1A1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1397),
.A2(n_1307),
.B(n_1417),
.C(n_1282),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1421),
.A2(n_1307),
.B(n_1296),
.C(n_1298),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1385),
.B(n_1322),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1329),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1377),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1351),
.A2(n_1319),
.B(n_1401),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1406),
.A2(n_1307),
.B(n_1296),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1384),
.B(n_1418),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_1334),
.B(n_1056),
.Y(n_1500)
);

AOI221x1_ASAP7_75t_SL g1501 ( 
.A1(n_1432),
.A2(n_1307),
.B1(n_730),
.B2(n_1306),
.C(n_1276),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1359),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1429),
.B(n_1366),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1384),
.B(n_1418),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1352),
.B(n_1366),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1406),
.A2(n_1307),
.B(n_1296),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1429),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1385),
.B(n_1322),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1352),
.B(n_1366),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1429),
.B(n_1366),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1329),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1406),
.A2(n_1307),
.B(n_1296),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1384),
.B(n_1418),
.Y(n_1513)
);

O2A1O1Ixp5_ASAP7_75t_L g1514 ( 
.A1(n_1321),
.A2(n_1307),
.B(n_1303),
.C(n_1293),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1352),
.B(n_1366),
.Y(n_1515)
);

NOR2xp67_ASAP7_75t_L g1516 ( 
.A(n_1334),
.B(n_1056),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1466),
.B(n_1471),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1502),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1442),
.B(n_1497),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1489),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1461),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1507),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1489),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1461),
.B(n_1459),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1484),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1445),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1461),
.B(n_1490),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1434),
.A2(n_1468),
.B(n_1479),
.Y(n_1528)
);

BUFx4f_ASAP7_75t_SL g1529 ( 
.A(n_1460),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1484),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1466),
.B(n_1471),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1464),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1437),
.B(n_1499),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1497),
.B(n_1455),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1483),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1437),
.B(n_1499),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1491),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1447),
.B(n_1486),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1504),
.B(n_1513),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1491),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1487),
.B(n_1457),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1504),
.B(n_1513),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1475),
.B(n_1464),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1446),
.B(n_1436),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1470),
.A2(n_1514),
.B(n_1485),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1473),
.B(n_1478),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1507),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1456),
.B(n_1472),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1456),
.B(n_1472),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1462),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1501),
.B(n_1453),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1463),
.A2(n_1492),
.B(n_1498),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1488),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1438),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1476),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1476),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1450),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1477),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1465),
.A2(n_1469),
.B(n_1453),
.Y(n_1559)
);

BUFx4f_ASAP7_75t_SL g1560 ( 
.A(n_1480),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1465),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1501),
.B(n_1449),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1448),
.B(n_1503),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1510),
.B(n_1481),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1481),
.B(n_1435),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1508),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1441),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1534),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1517),
.B(n_1506),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1517),
.B(n_1512),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1524),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1531),
.B(n_1469),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1552),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1528),
.B(n_1494),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1562),
.A2(n_1444),
.B1(n_1452),
.B2(n_1493),
.C(n_1451),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1528),
.B(n_1515),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1565),
.B(n_1452),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1505),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1531),
.B(n_1467),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1528),
.B(n_1509),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1525),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1518),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1552),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1518),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1530),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1526),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1526),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1569),
.B(n_1523),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1569),
.B(n_1523),
.Y(n_1591)
);

OAI33xp33_ASAP7_75t_L g1592 ( 
.A1(n_1570),
.A2(n_1562),
.A3(n_1551),
.B1(n_1565),
.B2(n_1563),
.B3(n_1557),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1579),
.A2(n_1577),
.B1(n_1551),
.B2(n_1555),
.C(n_1556),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1577),
.A2(n_1546),
.B1(n_1555),
.B2(n_1556),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1579),
.B(n_1563),
.Y(n_1595)
);

AOI33xp33_ASAP7_75t_L g1596 ( 
.A1(n_1578),
.A2(n_1557),
.A3(n_1548),
.B1(n_1549),
.B2(n_1541),
.B3(n_1561),
.Y(n_1596)
);

AOI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1570),
.A2(n_1537),
.B(n_1540),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1523),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1577),
.A2(n_1552),
.B(n_1444),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1588),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1569),
.B(n_1523),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1567),
.B(n_1521),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1588),
.Y(n_1603)
);

OAI211xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1570),
.A2(n_1564),
.B(n_1542),
.C(n_1533),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1571),
.A2(n_1546),
.B1(n_1548),
.B2(n_1549),
.C(n_1561),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1575),
.B(n_1546),
.Y(n_1606)
);

NAND4xp25_ASAP7_75t_SL g1607 ( 
.A(n_1571),
.B(n_1548),
.C(n_1549),
.D(n_1543),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1581),
.B(n_1454),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1588),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1571),
.A2(n_1552),
.B1(n_1541),
.B2(n_1564),
.C(n_1550),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1575),
.A2(n_1559),
.B(n_1546),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1589),
.Y(n_1612)
);

OAI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1573),
.A2(n_1546),
.B1(n_1559),
.B2(n_1532),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1575),
.B(n_1522),
.C(n_1543),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1566),
.A2(n_1559),
.B1(n_1546),
.B2(n_1524),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1575),
.A2(n_1559),
.B1(n_1532),
.B2(n_1524),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1574),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1573),
.A2(n_1559),
.B1(n_1532),
.B2(n_1558),
.Y(n_1618)
);

INVx5_ASAP7_75t_L g1619 ( 
.A(n_1575),
.Y(n_1619)
);

AOI222xp33_ASAP7_75t_L g1620 ( 
.A1(n_1585),
.A2(n_1541),
.B1(n_1543),
.B2(n_1550),
.C1(n_1533),
.C2(n_1542),
.Y(n_1620)
);

AND2x4_ASAP7_75t_SL g1621 ( 
.A(n_1566),
.B(n_1527),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1585),
.A2(n_1544),
.B1(n_1536),
.B2(n_1539),
.C(n_1522),
.Y(n_1622)
);

OAI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1573),
.A2(n_1544),
.B(n_1545),
.C(n_1547),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1578),
.B(n_1538),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1600),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1603),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1611),
.A2(n_1597),
.B(n_1623),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1619),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1609),
.Y(n_1629)
);

INVx4_ASAP7_75t_SL g1630 ( 
.A(n_1606),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1596),
.B(n_1578),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1604),
.B(n_1553),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1619),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

AO21x1_ASAP7_75t_L g1635 ( 
.A1(n_1599),
.A2(n_1584),
.B(n_1586),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1617),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_SL g1637 ( 
.A(n_1610),
.B(n_1554),
.C(n_1581),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1597),
.A2(n_1587),
.B(n_1583),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1590),
.B(n_1576),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1592),
.B(n_1553),
.Y(n_1640)
);

OA21x2_ASAP7_75t_L g1641 ( 
.A1(n_1616),
.A2(n_1587),
.B(n_1583),
.Y(n_1641)
);

OR2x6_ASAP7_75t_L g1642 ( 
.A(n_1606),
.B(n_1527),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1606),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.B(n_1578),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1634),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1634),
.Y(n_1646)
);

AND2x2_ASAP7_75t_SL g1647 ( 
.A(n_1627),
.B(n_1596),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1638),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1625),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1632),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1640),
.A2(n_1595),
.B1(n_1631),
.B2(n_1627),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1632),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1643),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1631),
.B(n_1624),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1621),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1625),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1643),
.B(n_1621),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1628),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1626),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1626),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.B(n_1614),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1640),
.B(n_1620),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1593),
.C(n_1605),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1638),
.Y(n_1667)
);

AOI21xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1627),
.A2(n_1594),
.B(n_1443),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1601),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1637),
.A2(n_1615),
.B1(n_1608),
.B2(n_1622),
.C(n_1606),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1619),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1627),
.A2(n_1496),
.B1(n_1439),
.B2(n_1495),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1628),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1628),
.B(n_1619),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1629),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1628),
.B(n_1619),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1633),
.B(n_1607),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1660),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1680),
.B(n_1633),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1647),
.B(n_1642),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1642),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1675),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1675),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1618),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1662),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1649),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1649),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1656),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1665),
.A2(n_1633),
.B(n_1582),
.C(n_1580),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1656),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1665),
.B(n_1560),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1680),
.B(n_1642),
.Y(n_1695)
);

AOI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1663),
.A2(n_1635),
.B(n_1627),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1678),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1651),
.B(n_1567),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1653),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1653),
.B(n_1664),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1678),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1652),
.Y(n_1702)
);

NOR2xp67_ASAP7_75t_L g1703 ( 
.A(n_1658),
.B(n_1633),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1654),
.B(n_1644),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1645),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1645),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1663),
.A2(n_1641),
.B(n_1613),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1654),
.B(n_1664),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1655),
.B(n_1642),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1650),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1677),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1652),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1671),
.A2(n_1568),
.B1(n_1572),
.B2(n_1644),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1655),
.B(n_1636),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1646),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1657),
.B(n_1636),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1646),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1696),
.B(n_1668),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1712),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1671),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1699),
.B(n_1681),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1702),
.Y(n_1722)
);

CKINVDCx16_ASAP7_75t_R g1723 ( 
.A(n_1682),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1700),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1674),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1689),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1681),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1688),
.B(n_1674),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1707),
.A2(n_1635),
.B1(n_1666),
.B2(n_1659),
.Y(n_1731)
);

NOR2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1682),
.B(n_1496),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1689),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1685),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1677),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1690),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1690),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1695),
.B(n_1659),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1687),
.A2(n_1635),
.B1(n_1669),
.B2(n_1666),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1695),
.B(n_1661),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1708),
.B(n_1529),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1708),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1703),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1709),
.B(n_1661),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1727),
.B(n_1745),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1731),
.A2(n_1692),
.B1(n_1713),
.B2(n_1668),
.C(n_1698),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1718),
.A2(n_1673),
.B(n_1683),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1723),
.B(n_1727),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1729),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1729),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1723),
.B(n_1745),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1719),
.B(n_1686),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1729),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1738),
.B(n_1709),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1719),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1724),
.A2(n_1673),
.B1(n_1684),
.B2(n_1683),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1726),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1726),
.Y(n_1759)
);

OAI32xp33_ASAP7_75t_L g1760 ( 
.A1(n_1720),
.A2(n_1684),
.A3(n_1658),
.B1(n_1711),
.B2(n_1686),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1724),
.A2(n_1672),
.B1(n_1670),
.B2(n_1669),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1740),
.A2(n_1711),
.B1(n_1658),
.B2(n_1670),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1733),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1733),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_SL g1765 ( 
.A1(n_1722),
.A2(n_1715),
.B(n_1705),
.C(n_1706),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1738),
.B(n_1714),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1736),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1756),
.B(n_1742),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1749),
.B(n_1732),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1754),
.Y(n_1770)
);

XOR2x2_ASAP7_75t_L g1771 ( 
.A(n_1752),
.B(n_1721),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1749),
.B(n_1743),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1753),
.B(n_1722),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1754),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1750),
.B(n_1751),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1752),
.B(n_1721),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1758),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1746),
.B(n_1725),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1759),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1776),
.A2(n_1748),
.B(n_1747),
.C(n_1757),
.Y(n_1780)
);

AOI32xp33_ASAP7_75t_L g1781 ( 
.A1(n_1769),
.A2(n_1757),
.A3(n_1762),
.B1(n_1755),
.B2(n_1766),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1772),
.A2(n_1765),
.B1(n_1760),
.B2(n_1730),
.C(n_1767),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_SL g1783 ( 
.A(n_1773),
.B(n_1778),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1771),
.B(n_1766),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_SL g1785 ( 
.A(n_1768),
.B(n_1761),
.C(n_1744),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1775),
.A2(n_1765),
.B(n_1763),
.C(n_1764),
.Y(n_1786)
);

OAI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1775),
.A2(n_1658),
.B1(n_1735),
.B2(n_1770),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1777),
.A2(n_1732),
.B(n_1737),
.C(n_1736),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1774),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1779),
.B(n_1741),
.Y(n_1790)
);

OAI222xp33_ASAP7_75t_L g1791 ( 
.A1(n_1781),
.A2(n_1741),
.B1(n_1735),
.B2(n_1734),
.C1(n_1728),
.C2(n_1717),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1780),
.A2(n_1672),
.B(n_1728),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1783),
.Y(n_1793)
);

NOR4xp25_ASAP7_75t_L g1794 ( 
.A(n_1785),
.B(n_1782),
.C(n_1787),
.D(n_1784),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_1790),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1789),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1786),
.A2(n_1734),
.B1(n_1728),
.B2(n_1672),
.Y(n_1797)
);

NOR2x1_ASAP7_75t_L g1798 ( 
.A(n_1793),
.B(n_1788),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1796),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1797),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1794),
.B(n_1734),
.Y(n_1801)
);

NOR4xp25_ASAP7_75t_L g1802 ( 
.A(n_1791),
.B(n_1739),
.C(n_1737),
.D(n_1715),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1795),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1792),
.B(n_1496),
.Y(n_1804)
);

AOI222xp33_ASAP7_75t_L g1805 ( 
.A1(n_1801),
.A2(n_1739),
.B1(n_1697),
.B2(n_1691),
.C1(n_1701),
.C2(n_1693),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1798),
.Y(n_1806)
);

AOI211xp5_ASAP7_75t_L g1807 ( 
.A1(n_1802),
.A2(n_1500),
.B(n_1516),
.C(n_1672),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_SL g1808 ( 
.A(n_1803),
.B(n_1511),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1799),
.A2(n_1697),
.B(n_1693),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_R g1810 ( 
.A(n_1800),
.B(n_1676),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1806),
.B(n_1701),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1810),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1808),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1812),
.B(n_1804),
.Y(n_1814)
);

AOI322xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1813),
.A3(n_1805),
.B1(n_1811),
.B2(n_1809),
.C1(n_1807),
.C2(n_1676),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1815),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1815),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1816),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1817),
.B(n_1714),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1819),
.B(n_1716),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1818),
.A2(n_1440),
.B1(n_1458),
.B2(n_1474),
.Y(n_1821)
);

OAI22x1_ASAP7_75t_L g1822 ( 
.A1(n_1820),
.A2(n_1679),
.B1(n_1676),
.B2(n_1716),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1822),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1823),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1821),
.B1(n_1676),
.B2(n_1679),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1825),
.A2(n_1679),
.B1(n_1648),
.B2(n_1667),
.Y(n_1826)
);

AOI211xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1679),
.B(n_1482),
.C(n_1704),
.Y(n_1827)
);


endmodule