module fake_jpeg_21284_n_312 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_47),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_18),
.C(n_19),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_20),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_30),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_22),
.B1(n_18),
.B2(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_35),
.B1(n_25),
.B2(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_60),
.B1(n_53),
.B2(n_51),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_23),
.B1(n_22),
.B2(n_39),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_68),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_35),
.B1(n_32),
.B2(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_71),
.B1(n_54),
.B2(n_51),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_37),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_72),
.B(n_73),
.Y(n_88)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_75),
.Y(n_85)
);

AOI22x1_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_24),
.B1(n_34),
.B2(n_14),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_37),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_23),
.A3(n_37),
.B1(n_28),
.B2(n_15),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_25),
.C(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_53),
.Y(n_90)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_77),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_84),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_41),
.C(n_55),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_104),
.C(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_109),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_108),
.B1(n_69),
.B2(n_81),
.Y(n_132)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_61),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_64),
.C(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_77),
.B1(n_42),
.B2(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_62),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_44),
.B1(n_42),
.B2(n_34),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_21),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_84),
.B1(n_97),
.B2(n_109),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_123),
.B1(n_129),
.B2(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_100),
.B(n_96),
.Y(n_147)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_88),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_78),
.B1(n_57),
.B2(n_75),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_44),
.B(n_26),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_135),
.B(n_127),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_80),
.B(n_17),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_122),
.C(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_69),
.B1(n_81),
.B2(n_79),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_96),
.B1(n_102),
.B2(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_68),
.B1(n_34),
.B2(n_29),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_29),
.B1(n_26),
.B2(n_98),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_87),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_83),
.CI(n_90),
.CON(n_137),
.SN(n_137)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_129),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_152),
.B(n_125),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_24),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_143),
.C(n_111),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_85),
.B1(n_82),
.B2(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_162),
.B1(n_111),
.B2(n_115),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_108),
.C(n_85),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_93),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_146),
.B(n_151),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_124),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_164),
.B1(n_133),
.B2(n_110),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_92),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_99),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_13),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_95),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_95),
.B1(n_26),
.B2(n_19),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_113),
.B(n_12),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_11),
.B(n_1),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_167),
.B(n_2),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_170),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_137),
.B(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_115),
.B1(n_125),
.B2(n_120),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_186),
.B1(n_144),
.B2(n_158),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_178),
.B1(n_185),
.B2(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_180),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_146),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_176),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_177),
.C(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_113),
.C(n_121),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_110),
.B1(n_119),
.B2(n_19),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_14),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_14),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_159),
.B1(n_147),
.B2(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_148),
.A2(n_164),
.B1(n_160),
.B2(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_197),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_137),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_0),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_213),
.B1(n_217),
.B2(n_185),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_11),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_220),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_196),
.C(n_166),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_3),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_10),
.B(n_3),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_186),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_177),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_204),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_178),
.B1(n_190),
.B2(n_189),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_207),
.B1(n_211),
.B2(n_219),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_181),
.C(n_166),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_195),
.C(n_180),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_183),
.C(n_171),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_168),
.C(n_184),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_187),
.C(n_4),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_209),
.B1(n_198),
.B2(n_208),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_246),
.B1(n_256),
.B2(n_235),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_198),
.B1(n_215),
.B2(n_202),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_202),
.B1(n_215),
.B2(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_252),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_257),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_212),
.B1(n_222),
.B2(n_211),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_212),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_226),
.C(n_236),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_265),
.C(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_254),
.C(n_247),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_233),
.C(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_240),
.C(n_222),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_256),
.C(n_258),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_251),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_248),
.C(n_229),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_267),
.C(n_268),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_261),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_227),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_6),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_260),
.C(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_3),
.C(n_4),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_288),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_278),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

OA21x2_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_275),
.B(n_273),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_299),
.C(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_6),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_291),
.B(n_284),
.Y(n_303)
);

OA21x2_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_295),
.B(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_300),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_307),
.C(n_304),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_302),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_297),
.C(n_292),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_292),
.B(n_8),
.C(n_9),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_9),
.Y(n_312)
);


endmodule