module fake_netlist_6_339_n_3154 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_578, n_703, n_144, n_365, n_978, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_951, n_783, n_106, n_725, n_952, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_969, n_988, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_360, n_945, n_977, n_603, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_355, n_426, n_317, n_149, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3154);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_945;
input n_977;
input n_603;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3154;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_1923;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1517;
wire n_1867;
wire n_1393;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3107;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_1658;
wire n_2593;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_1543;
wire n_2811;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_1873;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1605;
wire n_1330;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_2908;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3069;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_1214;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3153;
wire n_1188;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_2377;
wire n_2178;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_1369;
wire n_2271;
wire n_1008;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_1208;
wire n_2775;
wire n_1627;
wire n_1164;
wire n_1295;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_2913;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_1952;
wire n_2573;
wire n_2646;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_3037;
wire n_1646;
wire n_1714;
wire n_1139;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_1913;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3148;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_1992;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_2990;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3109;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2315;
wire n_1733;
wire n_1077;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_2276;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_2327;
wire n_2201;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_1608;
wire n_2305;
wire n_2373;
wire n_1472;
wire n_2050;
wire n_2120;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_2872;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_2702;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_2649;
wire n_2721;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_2743;
wire n_1973;
wire n_2267;
wire n_3035;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3038;
wire n_2033;
wire n_3086;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_3130;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_1753;
wire n_3095;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_1322;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_3054;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_985),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_456),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_988),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_112),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_304),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_885),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_391),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_923),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_431),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_361),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_429),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_90),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_762),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_81),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_599),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_845),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_838),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_222),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_524),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_292),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_583),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_205),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_700),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_570),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_811),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_283),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_72),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_381),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_837),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_276),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_855),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_92),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_175),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_976),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_350),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_856),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_830),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_56),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_824),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_606),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_492),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_865),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_862),
.Y(n_1034)
);

BUFx10_ASAP7_75t_L g1035 ( 
.A(n_571),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_456),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_425),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_611),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_600),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_831),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_826),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_851),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_471),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_902),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_32),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_650),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_954),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_22),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_616),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_625),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_967),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_391),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_517),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_974),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_645),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_117),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_584),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_347),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_542),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_677),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_588),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_972),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_235),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_612),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_277),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_921),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_156),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_183),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_556),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_609),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_530),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_405),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_131),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_376),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_864),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_186),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_116),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_263),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_564),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_329),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_887),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_782),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_586),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_799),
.Y(n_1085)
);

BUFx10_ASAP7_75t_L g1086 ( 
.A(n_953),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_713),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_65),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_577),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_900),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_498),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_971),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_619),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_969),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_948),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_298),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_970),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_675),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_615),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_544),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_956),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_703),
.Y(n_1102)
);

BUFx5_ASAP7_75t_L g1103 ( 
.A(n_329),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_610),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_754),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_240),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_580),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_278),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_221),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_935),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_731),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_109),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_2),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_608),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_733),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_966),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_777),
.Y(n_1117)
);

BUFx5_ASAP7_75t_L g1118 ( 
.A(n_659),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_743),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_786),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_532),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_571),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_296),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_17),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_832),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_983),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_46),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_145),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_396),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_282),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_503),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_899),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_361),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_285),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_681),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_142),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_984),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_957),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_581),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_622),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_284),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_2),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_642),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_781),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_655),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_940),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_326),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_836),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_927),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_770),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_576),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_717),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_792),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_651),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_404),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_171),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_138),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_821),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_402),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_12),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_610),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_955),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_943),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_776),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_161),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_638),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_820),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_614),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_626),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_53),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_550),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_150),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_795),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_641),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_261),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_435),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_48),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_632),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_495),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_591),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_535),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_804),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_596),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_202),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_92),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_597),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_973),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_829),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_601),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_707),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_835),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_791),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_823),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_965),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_161),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_177),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_167),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_504),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_670),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_224),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_617),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_613),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_299),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_89),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_598),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_580),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_657),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_735),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_485),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_304),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_604),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_960),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_666),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_962),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_232),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_23),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_518),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_231),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_555),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_58),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_787),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_24),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_819),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_557),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_187),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_622),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_794),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_279),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_72),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_306),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_947),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_239),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_751),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_877),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_521),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_605),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_950),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_618),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_961),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_100),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_964),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_684),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_958),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_986),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_959),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_546),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_322),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_109),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_110),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_664),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_491),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_78),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_510),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_589),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_120),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_479),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_693),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_807),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_780),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_424),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_553),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_590),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_524),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_797),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_686),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_35),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_21),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_323),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_968),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_200),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_880),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_649),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_34),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_874),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_404),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_353),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_139),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_981),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_644),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_274),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_912),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_605),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_660),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_508),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_682),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_511),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_907),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_951),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_551),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_215),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_118),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_247),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_593),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_31),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_944),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_420),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_572),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_200),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_222),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_662),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_533),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_54),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_513),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_917),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_435),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_653),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_277),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_123),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_315),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_946),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_663),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_759),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_932),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_24),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_466),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_260),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_843),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_403),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_417),
.Y(n_1319)
);

CKINVDCx16_ASAP7_75t_R g1320 ( 
.A(n_949),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_893),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_280),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_918),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_415),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_81),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_727),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_812),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_463),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_234),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_621),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_904),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_745),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_48),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_490),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_555),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_513),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_128),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_100),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_879),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_114),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_295),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_469),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_630),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_209),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_639),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_529),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_20),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_269),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_945),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_99),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_661),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_167),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_478),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_687),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_80),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_499),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_117),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_592),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_678),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_602),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_275),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_281),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_579),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_606),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_769),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_410),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_989),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_387),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_578),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_526),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_336),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_243),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_445),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_916),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_883),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_351),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_83),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_552),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_765),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_509),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_221),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_911),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_152),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_778),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_768),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_157),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_462),
.Y(n_1387)
);

BUFx10_ASAP7_75t_L g1388 ( 
.A(n_4),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_705),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_629),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_643),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_464),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_587),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_91),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_975),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_977),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_519),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_496),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_241),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_540),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_603),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_291),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_784),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_395),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_352),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_585),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_147),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_216),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_108),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_138),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_616),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_528),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_895),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_132),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_582),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_245),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_607),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_405),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_889),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_106),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_325),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_594),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_210),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_246),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_560),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_654),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_264),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_398),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_939),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_148),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_177),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_231),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_108),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_896),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_963),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_595),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_903),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_256),
.Y(n_1438)
);

BUFx10_ASAP7_75t_L g1439 ( 
.A(n_343),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_328),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_88),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_515),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_620),
.Y(n_1443)
);

CKINVDCx16_ASAP7_75t_R g1444 ( 
.A(n_173),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_396),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_387),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1103),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1103),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1103),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_992),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1103),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1103),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_1186),
.Y(n_1453)
);

CKINVDCx16_ASAP7_75t_R g1454 ( 
.A(n_1444),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_994),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1024),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1024),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1004),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1061),
.Y(n_1459)
);

INVxp33_ASAP7_75t_L g1460 ( 
.A(n_1043),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1094),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1024),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_997),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1102),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1007),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1014),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1078),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1078),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1146),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1288),
.B(n_0),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1006),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1234),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_L g1473 ( 
.A(n_1288),
.B(n_1),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1078),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1079),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1025),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1079),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1079),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1310),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1364),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1364),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1407),
.B(n_1),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1364),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1311),
.B(n_3),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1027),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1300),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1380),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1327),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1044),
.B(n_4),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1326),
.B(n_6),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1035),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1380),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1380),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1391),
.B(n_6),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1359),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1020),
.B(n_5),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1030),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1029),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1031),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1118),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1128),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1155),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1226),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1235),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1260),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1290),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1303),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1382),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1334),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1009),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1010),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1011),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1040),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_999),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_1136),
.B(n_5),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1041),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1313),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1453),
.B(n_1193),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1456),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1457),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1489),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1462),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1450),
.B(n_1148),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1467),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1468),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1489),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1455),
.B(n_1213),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1475),
.Y(n_1529)
);

AND2x6_ASAP7_75t_L g1530 ( 
.A(n_1447),
.B(n_1187),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1477),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1478),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1463),
.B(n_1389),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1480),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1470),
.A2(n_1272),
.B(n_1082),
.Y(n_1535)
);

AO22x1_ASAP7_75t_L g1536 ( 
.A1(n_1490),
.A2(n_1017),
.B1(n_1141),
.B2(n_1012),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1481),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1483),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1487),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1465),
.B(n_1320),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1492),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1493),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1448),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1458),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1498),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1449),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1451),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1452),
.A2(n_1022),
.B(n_1016),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1514),
.B(n_1145),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1479),
.B(n_1259),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1511),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1499),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1501),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1502),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1466),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1503),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1504),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1505),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1506),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1454),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1507),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1500),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1476),
.B(n_1435),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1509),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1485),
.B(n_1008),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1497),
.B(n_1049),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1517),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1496),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1513),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1473),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1484),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1491),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1516),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1471),
.B(n_1028),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1549),
.B(n_1494),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1573),
.A2(n_1515),
.B1(n_1308),
.B2(n_1204),
.Y(n_1579)
);

AND2x6_ASAP7_75t_L g1580 ( 
.A(n_1571),
.B(n_1015),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_SL g1581 ( 
.A(n_1562),
.B(n_1426),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1567),
.B(n_1460),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1570),
.A2(n_1026),
.B1(n_1071),
.B2(n_1013),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1568),
.B(n_1459),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1521),
.B(n_1046),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1526),
.B(n_1047),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1556),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1538),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1569),
.B(n_1482),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1561),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1523),
.B(n_1461),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1554),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1552),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_L g1594 ( 
.A(n_1540),
.B(n_995),
.C(n_993),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1572),
.A2(n_1232),
.B1(n_1336),
.B2(n_1080),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1544),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1528),
.B(n_1464),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1535),
.B(n_1055),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1538),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1542),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1550),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1574),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1518),
.B(n_1355),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1533),
.B(n_1469),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1542),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1564),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1546),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1565),
.B(n_1472),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1547),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1543),
.B(n_1076),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1557),
.A2(n_998),
.B1(n_1000),
.B2(n_996),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1555),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1559),
.Y(n_1615)
);

BUFx10_ASAP7_75t_L g1616 ( 
.A(n_1574),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1560),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1536),
.A2(n_1023),
.B1(n_1037),
.B2(n_1001),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1575),
.B(n_1566),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1486),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1551),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1539),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1522),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_1083),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1524),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1525),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1530),
.B(n_1085),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1519),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1520),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1527),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1529),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1545),
.B(n_1086),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1558),
.Y(n_1633)
);

INVx5_ASAP7_75t_L g1634 ( 
.A(n_1563),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1534),
.B(n_1086),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1537),
.Y(n_1636)
);

AND2x6_ASAP7_75t_L g1637 ( 
.A(n_1531),
.B(n_1362),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1532),
.B(n_1163),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1541),
.Y(n_1639)
);

OR2x6_ASAP7_75t_L g1640 ( 
.A(n_1548),
.B(n_1057),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1530),
.B(n_1097),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1556),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1521),
.B(n_1160),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1538),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1552),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1573),
.B(n_1101),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1579),
.A2(n_1324),
.B1(n_1305),
.B2(n_1038),
.C(n_1054),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1593),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1597),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_SL g1650 ( 
.A(n_1605),
.B(n_1495),
.C(n_1488),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1645),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1623),
.Y(n_1652)
);

AO22x2_ASAP7_75t_L g1653 ( 
.A1(n_1618),
.A2(n_1405),
.B1(n_1404),
.B2(n_1224),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1582),
.B(n_1033),
.Y(n_1654)
);

AO22x2_ASAP7_75t_L g1655 ( 
.A1(n_1578),
.A2(n_1112),
.B1(n_1238),
.B2(n_1058),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1034),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1626),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1583),
.A2(n_1062),
.B1(n_1068),
.B2(n_1036),
.C(n_1018),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1630),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1603),
.A2(n_1508),
.B1(n_1119),
.B2(n_1120),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1596),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1636),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1614),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1592),
.B(n_1072),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1628),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1584),
.B(n_1002),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1588),
.B(n_1074),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1615),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1617),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1629),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1611),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1619),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1602),
.B(n_1099),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1646),
.A2(n_1108),
.B1(n_1121),
.B2(n_1113),
.C(n_1109),
.Y(n_1675)
);

OAI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1594),
.A2(n_1130),
.B1(n_1157),
.B2(n_1147),
.C(n_1133),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1621),
.Y(n_1677)
);

AO22x2_ASAP7_75t_L g1678 ( 
.A1(n_1613),
.A2(n_1280),
.B1(n_1297),
.B2(n_1273),
.Y(n_1678)
);

AO22x2_ASAP7_75t_L g1679 ( 
.A1(n_1635),
.A2(n_1291),
.B1(n_1329),
.B2(n_1282),
.Y(n_1679)
);

AO22x2_ASAP7_75t_L g1680 ( 
.A1(n_1632),
.A2(n_1348),
.B1(n_1366),
.B2(n_1319),
.Y(n_1680)
);

NAND2x1p5_ASAP7_75t_L g1681 ( 
.A(n_1577),
.B(n_1042),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1616),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1639),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1644),
.B(n_1159),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1577),
.B(n_1051),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1608),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1633),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1589),
.B(n_1035),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1585),
.A2(n_1176),
.B1(n_1179),
.B2(n_1175),
.C(n_1170),
.Y(n_1689)
);

AO22x2_ASAP7_75t_L g1690 ( 
.A1(n_1643),
.A2(n_1420),
.B1(n_1401),
.B2(n_1195),
.Y(n_1690)
);

AO22x2_ASAP7_75t_L g1691 ( 
.A1(n_1581),
.A2(n_1202),
.B1(n_1430),
.B2(n_1209),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1622),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1608),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1604),
.B(n_1180),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1631),
.Y(n_1695)
);

AO22x2_ASAP7_75t_L g1696 ( 
.A1(n_1638),
.A2(n_1315),
.B1(n_1377),
.B2(n_1251),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1631),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1591),
.B(n_1003),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1587),
.B(n_1590),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1590),
.B(n_1598),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1640),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1599),
.B(n_1185),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1607),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1606),
.A2(n_1126),
.B1(n_1132),
.B2(n_1117),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1598),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1642),
.B(n_1219),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1601),
.B(n_1607),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1586),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1600),
.Y(n_1709)
);

BUFx2_ASAP7_75t_SL g1710 ( 
.A(n_1634),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1610),
.B(n_1005),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1612),
.B(n_1052),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1624),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1637),
.Y(n_1714)
);

AO22x2_ASAP7_75t_L g1715 ( 
.A1(n_1595),
.A2(n_1381),
.B1(n_1421),
.B2(n_1261),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1627),
.B(n_1056),
.Y(n_1716)
);

AND2x6_ASAP7_75t_L g1717 ( 
.A(n_1620),
.B(n_1063),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1580),
.Y(n_1718)
);

AOI22x1_ASAP7_75t_L g1719 ( 
.A1(n_1641),
.A2(n_1152),
.B1(n_1207),
.B2(n_1090),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1582),
.B(n_1067),
.Y(n_1720)
);

AO22x2_ASAP7_75t_L g1721 ( 
.A1(n_1605),
.A2(n_1402),
.B1(n_1220),
.B2(n_1253),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1582),
.B(n_1087),
.Y(n_1722)
);

AO22x2_ASAP7_75t_L g1723 ( 
.A1(n_1605),
.A2(n_1409),
.B1(n_1256),
.B2(n_1263),
.Y(n_1723)
);

NAND2x1p5_ASAP7_75t_L g1724 ( 
.A(n_1592),
.B(n_1092),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1593),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1603),
.A2(n_1227),
.B1(n_1239),
.B2(n_1208),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1593),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1579),
.A2(n_1270),
.B1(n_1309),
.B2(n_1267),
.C(n_1246),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1582),
.B(n_1095),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1593),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1628),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1582),
.Y(n_1732)
);

NAND2x1_ASAP7_75t_L g1733 ( 
.A(n_1609),
.B(n_1187),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1582),
.B(n_1098),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1592),
.B(n_1105),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1593),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1579),
.A2(n_1335),
.B1(n_1360),
.B2(n_1330),
.C(n_1314),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1593),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1603),
.B(n_1361),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1616),
.Y(n_1740)
);

NAND2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1592),
.B(n_1110),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1628),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1640),
.A2(n_1403),
.B1(n_1279),
.B2(n_1115),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1582),
.B(n_1111),
.Y(n_1744)
);

AO22x2_ASAP7_75t_L g1745 ( 
.A1(n_1605),
.A2(n_1398),
.B1(n_1406),
.B2(n_1387),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1582),
.B(n_1185),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1593),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1603),
.A2(n_1125),
.B1(n_1137),
.B2(n_1116),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1616),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1640),
.A2(n_1138),
.B1(n_1150),
.B2(n_1149),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_L g1751 ( 
.A(n_1600),
.B(n_1135),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1582),
.B(n_1154),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1628),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1577),
.Y(n_1754)
);

AO22x2_ASAP7_75t_L g1755 ( 
.A1(n_1605),
.A2(n_1408),
.B1(n_1411),
.B2(n_1410),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1640),
.A2(n_1166),
.B1(n_1173),
.B2(n_1169),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1592),
.B(n_1415),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1628),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1603),
.A2(n_1143),
.B1(n_1153),
.B2(n_1144),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1582),
.B(n_1178),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1593),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1640),
.A2(n_1244),
.B1(n_1257),
.B2(n_1250),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1628),
.Y(n_1763)
);

AND2x2_ASAP7_75t_SL g1764 ( 
.A(n_1581),
.B(n_1075),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1593),
.Y(n_1765)
);

AO22x2_ASAP7_75t_L g1766 ( 
.A1(n_1605),
.A2(n_1425),
.B1(n_1428),
.B2(n_1422),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1580),
.A2(n_1089),
.B1(n_1091),
.B2(n_1053),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1592),
.B(n_1265),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1718),
.B(n_1107),
.Y(n_1769)
);

NAND2xp33_ASAP7_75t_SL g1770 ( 
.A(n_1714),
.B(n_1124),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1673),
.B(n_1764),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1708),
.B(n_1158),
.Y(n_1772)
);

NAND2xp33_ASAP7_75t_SL g1773 ( 
.A(n_1702),
.B(n_1168),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_SL g1774 ( 
.A(n_1746),
.B(n_1197),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1654),
.B(n_1162),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1720),
.B(n_1164),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1722),
.B(n_1167),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1729),
.B(n_1174),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1734),
.B(n_1182),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1744),
.B(n_1188),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1752),
.B(n_1190),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1760),
.B(n_1667),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1698),
.B(n_1711),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1713),
.B(n_1191),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1709),
.B(n_1192),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1648),
.B(n_1194),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1649),
.B(n_1651),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1652),
.B(n_1199),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1657),
.B(n_1212),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1658),
.B(n_1660),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1663),
.B(n_1214),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1664),
.B(n_1221),
.Y(n_1792)
);

NAND2xp33_ASAP7_75t_SL g1793 ( 
.A(n_1682),
.B(n_1749),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_SL g1794 ( 
.A(n_1701),
.B(n_1217),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1669),
.B(n_1223),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1662),
.B(n_1225),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1670),
.B(n_1274),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1672),
.B(n_1231),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1725),
.B(n_1233),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1727),
.B(n_1306),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1730),
.B(n_1312),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1736),
.B(n_1237),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1738),
.B(n_1242),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1747),
.B(n_1243),
.Y(n_1804)
);

NAND2xp33_ASAP7_75t_SL g1805 ( 
.A(n_1750),
.B(n_1248),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1761),
.B(n_1245),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1765),
.B(n_1258),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1688),
.B(n_1218),
.Y(n_1808)
);

NAND2xp33_ASAP7_75t_SL g1809 ( 
.A(n_1756),
.B(n_1268),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1687),
.B(n_1704),
.Y(n_1810)
);

NAND2xp33_ASAP7_75t_SL g1811 ( 
.A(n_1762),
.B(n_1307),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1661),
.B(n_1677),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1712),
.B(n_1666),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1743),
.B(n_1264),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1671),
.B(n_1323),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1739),
.B(n_1230),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1731),
.B(n_1332),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1692),
.B(n_1269),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1759),
.B(n_1271),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1700),
.B(n_1278),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1739),
.B(n_1230),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1686),
.B(n_1281),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1697),
.B(n_1283),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1742),
.B(n_1285),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1753),
.B(n_1287),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1758),
.B(n_1374),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1763),
.B(n_1295),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1683),
.B(n_1384),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1716),
.B(n_1304),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1693),
.B(n_1317),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1665),
.B(n_1388),
.Y(n_1831)
);

NAND2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1695),
.B(n_1341),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1757),
.B(n_1388),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1706),
.B(n_1439),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1656),
.B(n_1321),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1767),
.B(n_1331),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1699),
.B(n_1339),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1655),
.B(n_1717),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1705),
.B(n_1350),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1726),
.B(n_1345),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1748),
.B(n_1349),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1740),
.B(n_1354),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1754),
.B(n_1365),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1694),
.B(n_1367),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1703),
.B(n_1375),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1717),
.B(n_1385),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1668),
.B(n_1379),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1674),
.B(n_1390),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1684),
.B(n_1395),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1724),
.B(n_1396),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1751),
.B(n_1434),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1733),
.B(n_1438),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1735),
.B(n_1413),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1741),
.B(n_1419),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1721),
.B(n_1439),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1691),
.B(n_1429),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1768),
.B(n_1437),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1707),
.B(n_1163),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1723),
.B(n_1446),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1681),
.B(n_1343),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1745),
.B(n_1446),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1685),
.B(n_1187),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1719),
.B(n_1241),
.Y(n_1863)
);

NAND2xp33_ASAP7_75t_SL g1864 ( 
.A(n_1710),
.B(n_1019),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1650),
.B(n_1241),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1680),
.B(n_1241),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1679),
.B(n_1351),
.Y(n_1867)
);

NAND2xp33_ASAP7_75t_SL g1868 ( 
.A(n_1678),
.B(n_1021),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1755),
.B(n_1351),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1766),
.B(n_1351),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1696),
.B(n_1118),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1647),
.B(n_1032),
.Y(n_1872)
);

NAND2xp33_ASAP7_75t_SL g1873 ( 
.A(n_1728),
.B(n_1039),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1676),
.B(n_1045),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1737),
.B(n_1048),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1690),
.B(n_1050),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1715),
.B(n_1059),
.Y(n_1877)
);

NAND2xp33_ASAP7_75t_SL g1878 ( 
.A(n_1653),
.B(n_1060),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1675),
.B(n_1064),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1689),
.B(n_1065),
.Y(n_1880)
);

NAND2xp33_ASAP7_75t_SL g1881 ( 
.A(n_1659),
.B(n_1066),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1732),
.B(n_1069),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1732),
.B(n_1070),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1732),
.B(n_1073),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1732),
.B(n_1077),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_SL g1886 ( 
.A(n_1718),
.B(n_1081),
.Y(n_1886)
);

NAND2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1718),
.B(n_1084),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1732),
.B(n_1088),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1732),
.B(n_1093),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1732),
.B(n_1096),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1732),
.B(n_1104),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1732),
.B(n_1106),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1732),
.B(n_1114),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1732),
.B(n_1122),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1732),
.B(n_1123),
.Y(n_1895)
);

NAND2xp33_ASAP7_75t_SL g1896 ( 
.A(n_1718),
.B(n_1127),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1732),
.B(n_1129),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1732),
.B(n_1131),
.Y(n_1898)
);

NAND2xp33_ASAP7_75t_SL g1899 ( 
.A(n_1718),
.B(n_1134),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1732),
.B(n_1139),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1732),
.B(n_1140),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1732),
.B(n_1142),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1732),
.B(n_1156),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1732),
.B(n_1161),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1732),
.B(n_1165),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1732),
.B(n_1171),
.Y(n_1906)
);

XNOR2xp5_ASAP7_75t_L g1907 ( 
.A(n_1662),
.B(n_623),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1732),
.B(n_1172),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1732),
.B(n_1177),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1732),
.B(n_1181),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1718),
.B(n_1183),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1732),
.B(n_1184),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1732),
.B(n_1196),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1732),
.B(n_1198),
.Y(n_1914)
);

AND2x2_ASAP7_75t_SL g1915 ( 
.A(n_1764),
.B(n_1100),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1732),
.B(n_1200),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1732),
.B(n_1201),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1732),
.B(n_1203),
.Y(n_1918)
);

NAND2xp33_ASAP7_75t_SL g1919 ( 
.A(n_1718),
.B(n_1206),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1718),
.B(n_1210),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1732),
.B(n_1211),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1732),
.B(n_1215),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1732),
.B(n_1216),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1697),
.B(n_1151),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1732),
.B(n_1222),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1732),
.B(n_1228),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1732),
.B(n_1229),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1732),
.B(n_1236),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1732),
.B(n_1240),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1732),
.B(n_1247),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1732),
.B(n_1249),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1732),
.B(n_1252),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1732),
.B(n_1254),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1732),
.B(n_1255),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1732),
.B(n_1262),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1732),
.B(n_1266),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1732),
.B(n_1275),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1732),
.B(n_1276),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1732),
.B(n_1277),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1732),
.B(n_1286),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1732),
.B(n_1289),
.Y(n_1941)
);

NAND2xp33_ASAP7_75t_SL g1942 ( 
.A(n_1718),
.B(n_1292),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1796),
.Y(n_1943)
);

AOI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1805),
.A2(n_1296),
.B1(n_1298),
.B2(n_1294),
.C(n_1293),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1783),
.A2(n_1782),
.B(n_1813),
.Y(n_1945)
);

NAND3xp33_ASAP7_75t_SL g1946 ( 
.A(n_1773),
.B(n_1301),
.C(n_1299),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1790),
.Y(n_1947)
);

AO32x2_ASAP7_75t_L g1948 ( 
.A1(n_1838),
.A2(n_9),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1924),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_SL g1950 ( 
.A1(n_1846),
.A2(n_1205),
.B(n_1189),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1771),
.B(n_1928),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1787),
.Y(n_1952)
);

OA21x2_ASAP7_75t_L g1953 ( 
.A1(n_1828),
.A2(n_1302),
.B(n_1284),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1915),
.A2(n_1417),
.B(n_1440),
.C(n_1372),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1815),
.A2(n_1445),
.B(n_627),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1897),
.B(n_1909),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1883),
.B(n_1316),
.Y(n_1957)
);

O2A1O1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1812),
.A2(n_1322),
.B(n_1325),
.C(n_1318),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1834),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1888),
.B(n_1328),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1817),
.A2(n_628),
.B(n_624),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1901),
.B(n_1333),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1903),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1810),
.A2(n_1338),
.B(n_1337),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1826),
.A2(n_633),
.B(n_631),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1797),
.Y(n_1966)
);

INVx4_ASAP7_75t_L g1967 ( 
.A(n_1852),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1904),
.B(n_1913),
.Y(n_1968)
);

OAI21x1_ASAP7_75t_L g1969 ( 
.A1(n_1800),
.A2(n_635),
.B(n_634),
.Y(n_1969)
);

AO31x2_ASAP7_75t_L g1970 ( 
.A1(n_1851),
.A2(n_637),
.A3(n_640),
.B(n_636),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1918),
.A2(n_1342),
.B1(n_1344),
.B2(n_1340),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1852),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1922),
.B(n_1346),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1801),
.Y(n_1974)
);

NOR2xp67_ASAP7_75t_L g1975 ( 
.A(n_1925),
.B(n_646),
.Y(n_1975)
);

AO31x2_ASAP7_75t_L g1976 ( 
.A1(n_1856),
.A2(n_648),
.A3(n_652),
.B(n_647),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1863),
.A2(n_658),
.B(n_656),
.Y(n_1977)
);

OAI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1824),
.A2(n_667),
.B(n_665),
.Y(n_1978)
);

BUFx2_ASAP7_75t_L g1979 ( 
.A(n_1832),
.Y(n_1979)
);

NAND2x2_ASAP7_75t_L g1980 ( 
.A(n_1876),
.B(n_1347),
.Y(n_1980)
);

OAI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1933),
.A2(n_1353),
.B1(n_1356),
.B2(n_1352),
.Y(n_1981)
);

NAND3xp33_ASAP7_75t_L g1982 ( 
.A(n_1774),
.B(n_1358),
.C(n_1357),
.Y(n_1982)
);

OAI21x1_ASAP7_75t_L g1983 ( 
.A1(n_1825),
.A2(n_669),
.B(n_668),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1871),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1785),
.B(n_1772),
.Y(n_1985)
);

OAI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1827),
.A2(n_672),
.B(n_671),
.Y(n_1986)
);

OAI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1822),
.A2(n_674),
.B(n_673),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1808),
.B(n_1363),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1775),
.B(n_1368),
.Y(n_1989)
);

A2O1A1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1873),
.A2(n_1811),
.B(n_1809),
.C(n_1881),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1818),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1769),
.B(n_1369),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1907),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1867),
.Y(n_1994)
);

OA22x2_ASAP7_75t_L g1995 ( 
.A1(n_1855),
.A2(n_1371),
.B1(n_1373),
.B2(n_1370),
.Y(n_1995)
);

AO31x2_ASAP7_75t_L g1996 ( 
.A1(n_1865),
.A2(n_679),
.A3(n_680),
.B(n_676),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1784),
.A2(n_685),
.B(n_683),
.Y(n_1997)
);

NAND2x1_ASAP7_75t_L g1998 ( 
.A(n_1831),
.B(n_688),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1833),
.B(n_689),
.Y(n_1999)
);

NAND2x1p5_ASAP7_75t_L g2000 ( 
.A(n_1837),
.B(n_690),
.Y(n_2000)
);

AOI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1786),
.A2(n_1789),
.B(n_1788),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1776),
.A2(n_1378),
.B1(n_1383),
.B2(n_1376),
.Y(n_2002)
);

BUFx12f_ASAP7_75t_L g2003 ( 
.A(n_1816),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1820),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1777),
.B(n_1386),
.Y(n_2005)
);

AO31x2_ASAP7_75t_L g2006 ( 
.A1(n_1866),
.A2(n_692),
.A3(n_694),
.B(n_691),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1821),
.B(n_695),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1791),
.A2(n_697),
.B(n_696),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1792),
.A2(n_699),
.B(n_698),
.Y(n_2009)
);

AO31x2_ASAP7_75t_L g2010 ( 
.A1(n_1868),
.A2(n_702),
.A3(n_704),
.B(n_701),
.Y(n_2010)
);

AOI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1795),
.A2(n_708),
.B(n_706),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1882),
.B(n_1392),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1823),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1798),
.A2(n_710),
.B(n_709),
.Y(n_2014)
);

BUFx4_ASAP7_75t_SL g2015 ( 
.A(n_1793),
.Y(n_2015)
);

AOI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1799),
.A2(n_712),
.B(n_711),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1845),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1875),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1778),
.A2(n_1394),
.B(n_1393),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1802),
.Y(n_2020)
);

INVx2_ASAP7_75t_SL g2021 ( 
.A(n_1877),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1779),
.B(n_1397),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1859),
.Y(n_2023)
);

A2O1A1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_1770),
.A2(n_1400),
.B(n_1412),
.C(n_1399),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_SL g2025 ( 
.A1(n_1850),
.A2(n_715),
.B(n_714),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1803),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_1780),
.A2(n_1416),
.B1(n_1418),
.B2(n_1414),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1804),
.A2(n_718),
.B(n_716),
.Y(n_2028)
);

BUFx6f_ASAP7_75t_L g2029 ( 
.A(n_1842),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1806),
.Y(n_2030)
);

OAI21x1_ASAP7_75t_L g2031 ( 
.A1(n_1830),
.A2(n_720),
.B(n_719),
.Y(n_2031)
);

NAND3x1_ASAP7_75t_L g2032 ( 
.A(n_1861),
.B(n_1424),
.C(n_1423),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1807),
.A2(n_722),
.B(n_721),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1843),
.Y(n_2034)
);

OR2x6_ASAP7_75t_L g2035 ( 
.A(n_1869),
.B(n_7),
.Y(n_2035)
);

AO31x2_ASAP7_75t_L g2036 ( 
.A1(n_1781),
.A2(n_724),
.A3(n_725),
.B(n_723),
.Y(n_2036)
);

OAI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1835),
.A2(n_1829),
.B(n_1840),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1839),
.Y(n_2038)
);

AOI221x1_ASAP7_75t_L g2039 ( 
.A1(n_1878),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_1794),
.Y(n_2040)
);

OAI21x1_ASAP7_75t_L g2041 ( 
.A1(n_1819),
.A2(n_728),
.B(n_726),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1814),
.A2(n_730),
.B(n_729),
.Y(n_2042)
);

AO32x2_ASAP7_75t_L g2043 ( 
.A1(n_1870),
.A2(n_13),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1874),
.Y(n_2044)
);

AO21x1_ASAP7_75t_L g2045 ( 
.A1(n_1886),
.A2(n_1896),
.B(n_1887),
.Y(n_2045)
);

OAI21x1_ASAP7_75t_L g2046 ( 
.A1(n_1853),
.A2(n_734),
.B(n_732),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1872),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1847),
.A2(n_737),
.B(n_736),
.Y(n_2048)
);

OA21x2_ASAP7_75t_L g2049 ( 
.A1(n_1849),
.A2(n_1431),
.B(n_1427),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_1844),
.A2(n_739),
.B(n_738),
.Y(n_2050)
);

BUFx12f_ASAP7_75t_L g2051 ( 
.A(n_1864),
.Y(n_2051)
);

AO31x2_ASAP7_75t_L g2052 ( 
.A1(n_1899),
.A2(n_741),
.A3(n_742),
.B(n_740),
.Y(n_2052)
);

OR2x6_ASAP7_75t_L g2053 ( 
.A(n_1858),
.B(n_13),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1884),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1885),
.B(n_1432),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1848),
.A2(n_746),
.B(n_744),
.Y(n_2056)
);

BUFx12f_ASAP7_75t_L g2057 ( 
.A(n_1911),
.Y(n_2057)
);

OAI21x1_ASAP7_75t_L g2058 ( 
.A1(n_1854),
.A2(n_748),
.B(n_747),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1889),
.B(n_1433),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_SL g2060 ( 
.A1(n_1919),
.A2(n_1942),
.B(n_1920),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1879),
.Y(n_2061)
);

AO31x2_ASAP7_75t_L g2062 ( 
.A1(n_1880),
.A2(n_990),
.A3(n_991),
.B(n_987),
.Y(n_2062)
);

AO31x2_ASAP7_75t_L g2063 ( 
.A1(n_1841),
.A2(n_1857),
.A3(n_1836),
.B(n_1890),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1891),
.A2(n_750),
.B(n_749),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1892),
.B(n_1436),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_1862),
.A2(n_753),
.B(n_752),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_1893),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1894),
.A2(n_1442),
.B1(n_1443),
.B2(n_1441),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1895),
.A2(n_756),
.B(n_755),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1898),
.A2(n_758),
.B(n_757),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1900),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1902),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1905),
.A2(n_761),
.B(n_760),
.Y(n_2073)
);

INVx8_ASAP7_75t_L g2074 ( 
.A(n_2003),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1947),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1955),
.A2(n_2041),
.B(n_2037),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1951),
.A2(n_1941),
.B1(n_1940),
.B2(n_1906),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1952),
.Y(n_2078)
);

OAI21x1_ASAP7_75t_L g2079 ( 
.A1(n_1978),
.A2(n_1860),
.B(n_1908),
.Y(n_2079)
);

INVx4_ASAP7_75t_L g2080 ( 
.A(n_1972),
.Y(n_2080)
);

OAI21x1_ASAP7_75t_L g2081 ( 
.A1(n_1983),
.A2(n_1912),
.B(n_1910),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_1986),
.A2(n_1916),
.B(n_1914),
.Y(n_2082)
);

OR2x6_ASAP7_75t_L g2083 ( 
.A(n_1959),
.B(n_1917),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1956),
.B(n_1934),
.Y(n_2084)
);

CKINVDCx8_ASAP7_75t_R g2085 ( 
.A(n_1943),
.Y(n_2085)
);

BUFx2_ASAP7_75t_R g2086 ( 
.A(n_1993),
.Y(n_2086)
);

INVx1_ASAP7_75t_SL g2087 ( 
.A(n_2071),
.Y(n_2087)
);

OAI222xp33_ASAP7_75t_L g2088 ( 
.A1(n_2035),
.A2(n_1927),
.B1(n_1923),
.B2(n_1929),
.C1(n_1926),
.C2(n_1921),
.Y(n_2088)
);

INVxp67_ASAP7_75t_SL g2089 ( 
.A(n_1966),
.Y(n_2089)
);

OAI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_1968),
.A2(n_1931),
.B1(n_1932),
.B2(n_1930),
.Y(n_2090)
);

OAI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_1944),
.A2(n_1936),
.B(n_1937),
.C(n_1935),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_1987),
.A2(n_1965),
.B(n_1961),
.Y(n_2092)
);

OR2x6_ASAP7_75t_L g2093 ( 
.A(n_2021),
.B(n_1938),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1974),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_2012),
.A2(n_1939),
.B1(n_16),
.B2(n_14),
.Y(n_2095)
);

O2A1O1Ixp33_ASAP7_75t_SL g2096 ( 
.A1(n_1990),
.A2(n_1984),
.B(n_1985),
.C(n_2018),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1963),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1949),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_1967),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_2029),
.Y(n_2100)
);

OA21x2_ASAP7_75t_L g2101 ( 
.A1(n_1945),
.A2(n_764),
.B(n_763),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_2031),
.A2(n_767),
.B(n_766),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1969),
.A2(n_772),
.B(n_771),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_2044),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_SL g2105 ( 
.A1(n_2055),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_2023),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1994),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_2046),
.A2(n_774),
.B(n_773),
.Y(n_2108)
);

BUFx2_ASAP7_75t_SL g2109 ( 
.A(n_1999),
.Y(n_2109)
);

OAI21x1_ASAP7_75t_L g2110 ( 
.A1(n_2058),
.A2(n_1977),
.B(n_2066),
.Y(n_2110)
);

BUFx8_ASAP7_75t_L g2111 ( 
.A(n_2029),
.Y(n_2111)
);

NAND3xp33_ASAP7_75t_SL g2112 ( 
.A(n_1964),
.B(n_18),
.C(n_19),
.Y(n_2112)
);

NOR2xp67_ASAP7_75t_SL g2113 ( 
.A(n_2051),
.B(n_20),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2061),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2047),
.Y(n_2115)
);

AOI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_2001),
.A2(n_779),
.B(n_775),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1957),
.A2(n_785),
.B(n_783),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_SL g2118 ( 
.A1(n_1979),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2118)
);

BUFx3_ASAP7_75t_L g2119 ( 
.A(n_2004),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_2042),
.A2(n_789),
.B(n_788),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_1950),
.A2(n_793),
.B(n_790),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1988),
.B(n_25),
.Y(n_2122)
);

OR2x6_ASAP7_75t_L g2123 ( 
.A(n_2057),
.B(n_796),
.Y(n_2123)
);

AO21x1_ASAP7_75t_L g2124 ( 
.A1(n_1958),
.A2(n_28),
.B(n_27),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1953),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2043),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_2004),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_1997),
.A2(n_800),
.B(n_798),
.Y(n_2128)
);

OR2x6_ASAP7_75t_L g2129 ( 
.A(n_1998),
.B(n_801),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2043),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1960),
.A2(n_803),
.B(n_802),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2008),
.A2(n_806),
.B(n_805),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_SL g2133 ( 
.A1(n_2045),
.A2(n_2060),
.B(n_2050),
.Y(n_2133)
);

NOR2x1_ASAP7_75t_SL g2134 ( 
.A(n_2026),
.B(n_808),
.Y(n_2134)
);

O2A1O1Ixp33_ASAP7_75t_L g2135 ( 
.A1(n_2024),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2038),
.B(n_26),
.Y(n_2136)
);

OAI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_1962),
.A2(n_810),
.B(n_809),
.Y(n_2137)
);

AO31x2_ASAP7_75t_L g2138 ( 
.A1(n_2039),
.A2(n_814),
.A3(n_815),
.B(n_813),
.Y(n_2138)
);

OR2x6_ASAP7_75t_L g2139 ( 
.A(n_2007),
.B(n_816),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2020),
.Y(n_2140)
);

OAI21x1_ASAP7_75t_L g2141 ( 
.A1(n_2009),
.A2(n_818),
.B(n_817),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1972),
.B(n_822),
.Y(n_2142)
);

OAI21x1_ASAP7_75t_L g2143 ( 
.A1(n_2011),
.A2(n_827),
.B(n_825),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_2072),
.Y(n_2144)
);

AO31x2_ASAP7_75t_L g2145 ( 
.A1(n_1954),
.A2(n_833),
.A3(n_834),
.B(n_828),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1948),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1948),
.Y(n_2147)
);

OAI21x1_ASAP7_75t_L g2148 ( 
.A1(n_2014),
.A2(n_840),
.B(n_839),
.Y(n_2148)
);

OAI21x1_ASAP7_75t_L g2149 ( 
.A1(n_2016),
.A2(n_2033),
.B(n_2028),
.Y(n_2149)
);

AO31x2_ASAP7_75t_L g2150 ( 
.A1(n_2056),
.A2(n_842),
.A3(n_844),
.B(n_841),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_2048),
.A2(n_847),
.B(n_846),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_SL g2152 ( 
.A1(n_2064),
.A2(n_849),
.B(n_848),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2054),
.B(n_29),
.Y(n_2153)
);

OA21x2_ASAP7_75t_L g2154 ( 
.A1(n_2030),
.A2(n_852),
.B(n_850),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2067),
.B(n_853),
.Y(n_2155)
);

AOI21xp5_ASAP7_75t_L g2156 ( 
.A1(n_1973),
.A2(n_857),
.B(n_854),
.Y(n_2156)
);

BUFx3_ASAP7_75t_L g2157 ( 
.A(n_2034),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2013),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1991),
.Y(n_2159)
);

OA21x2_ASAP7_75t_L g2160 ( 
.A1(n_2017),
.A2(n_859),
.B(n_858),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2040),
.A2(n_2005),
.B1(n_2022),
.B2(n_1989),
.Y(n_2161)
);

AO21x2_ASAP7_75t_L g2162 ( 
.A1(n_1975),
.A2(n_861),
.B(n_860),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_1946),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2006),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2062),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2025),
.A2(n_866),
.B(n_863),
.Y(n_2166)
);

OAI21x1_ASAP7_75t_L g2167 ( 
.A1(n_2069),
.A2(n_868),
.B(n_867),
.Y(n_2167)
);

OAI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2059),
.A2(n_870),
.B(n_869),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_1982),
.B(n_871),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2062),
.Y(n_2170)
);

OR2x6_ASAP7_75t_L g2171 ( 
.A(n_2053),
.B(n_872),
.Y(n_2171)
);

AND2x2_ASAP7_75t_SL g2172 ( 
.A(n_2049),
.B(n_33),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_1992),
.B(n_873),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_2070),
.A2(n_876),
.B(n_875),
.Y(n_2174)
);

OAI21x1_ASAP7_75t_L g2175 ( 
.A1(n_2073),
.A2(n_881),
.B(n_878),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_2000),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2036),
.Y(n_2177)
);

INVx1_ASAP7_75t_SL g2178 ( 
.A(n_2015),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_SL g2179 ( 
.A1(n_1995),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_2179)
);

AO21x2_ASAP7_75t_L g2180 ( 
.A1(n_2019),
.A2(n_884),
.B(n_882),
.Y(n_2180)
);

NOR2xp67_ASAP7_75t_R g2181 ( 
.A(n_1980),
.B(n_37),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1996),
.Y(n_2182)
);

O2A1O1Ixp33_ASAP7_75t_L g2183 ( 
.A1(n_1971),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2063),
.B(n_886),
.Y(n_2184)
);

O2A1O1Ixp33_ASAP7_75t_L g2185 ( 
.A1(n_1981),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1996),
.Y(n_2186)
);

BUFx4_ASAP7_75t_SL g2187 ( 
.A(n_2032),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_L g2188 ( 
.A1(n_2065),
.A2(n_890),
.B(n_888),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_SL g2189 ( 
.A1(n_2010),
.A2(n_892),
.B(n_891),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_2002),
.A2(n_897),
.B(n_894),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_2027),
.A2(n_901),
.B(n_898),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_2068),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2192)
);

OAI21x1_ASAP7_75t_L g2193 ( 
.A1(n_1970),
.A2(n_906),
.B(n_905),
.Y(n_2193)
);

O2A1O1Ixp33_ASAP7_75t_L g2194 ( 
.A1(n_2010),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1976),
.B(n_44),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2052),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_2052),
.B(n_908),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_1970),
.A2(n_910),
.B(n_909),
.Y(n_2198)
);

AO31x2_ASAP7_75t_L g2199 ( 
.A1(n_1990),
.A2(n_914),
.A3(n_915),
.B(n_913),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1947),
.B(n_49),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_2021),
.Y(n_2201)
);

BUFx3_ASAP7_75t_L g2202 ( 
.A(n_2111),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_2100),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2122),
.B(n_50),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2075),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2094),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2078),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2089),
.B(n_51),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2136),
.B(n_51),
.Y(n_2209)
);

AO21x2_ASAP7_75t_L g2210 ( 
.A1(n_2133),
.A2(n_920),
.B(n_919),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2158),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2107),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2140),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2119),
.B(n_922),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2098),
.Y(n_2215)
);

INVx1_ASAP7_75t_SL g2216 ( 
.A(n_2087),
.Y(n_2216)
);

NAND3xp33_ASAP7_75t_L g2217 ( 
.A(n_2095),
.B(n_52),
.C(n_53),
.Y(n_2217)
);

INVxp67_ASAP7_75t_L g2218 ( 
.A(n_2201),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_2085),
.Y(n_2219)
);

INVx2_ASAP7_75t_SL g2220 ( 
.A(n_2074),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2159),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_2157),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2179),
.B(n_54),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2115),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2144),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2105),
.B(n_55),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2114),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2104),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2125),
.Y(n_2229)
);

OA21x2_ASAP7_75t_L g2230 ( 
.A1(n_2164),
.A2(n_925),
.B(n_924),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2200),
.Y(n_2231)
);

OR2x2_ASAP7_75t_L g2232 ( 
.A(n_2084),
.B(n_55),
.Y(n_2232)
);

OR2x6_ASAP7_75t_L g2233 ( 
.A(n_2109),
.B(n_2139),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2177),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2096),
.Y(n_2235)
);

INVx8_ASAP7_75t_L g2236 ( 
.A(n_2139),
.Y(n_2236)
);

OA21x2_ASAP7_75t_L g2237 ( 
.A1(n_2076),
.A2(n_2170),
.B(n_2182),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2184),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2090),
.B(n_56),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_2127),
.Y(n_2240)
);

OAI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2161),
.A2(n_57),
.B(n_58),
.Y(n_2241)
);

OAI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2077),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.C(n_61),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2081),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2126),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2130),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_2080),
.Y(n_2246)
);

OR2x2_ASAP7_75t_SL g2247 ( 
.A(n_2112),
.B(n_59),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2082),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2153),
.Y(n_2249)
);

BUFx2_ASAP7_75t_L g2250 ( 
.A(n_2083),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2195),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2091),
.B(n_61),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_2106),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2192),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2146),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2147),
.Y(n_2256)
);

BUFx2_ASAP7_75t_L g2257 ( 
.A(n_2083),
.Y(n_2257)
);

INVx2_ASAP7_75t_SL g2258 ( 
.A(n_2178),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2199),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2149),
.A2(n_979),
.B(n_978),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2138),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2151),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2124),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2117),
.A2(n_982),
.B(n_980),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2196),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2093),
.B(n_62),
.Y(n_2266)
);

BUFx2_ASAP7_75t_L g2267 ( 
.A(n_2093),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2097),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2194),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2172),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2086),
.Y(n_2271)
);

HB1xp67_ASAP7_75t_L g2272 ( 
.A(n_2155),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2167),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2174),
.Y(n_2274)
);

NOR2x1_ASAP7_75t_SL g2275 ( 
.A(n_2129),
.B(n_926),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_2171),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2188),
.Y(n_2277)
);

NAND2x1p5_ASAP7_75t_L g2278 ( 
.A(n_2099),
.B(n_928),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2175),
.Y(n_2279)
);

AO21x2_ASAP7_75t_L g2280 ( 
.A1(n_2165),
.A2(n_930),
.B(n_929),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_2132),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2141),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2253),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2205),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2233),
.B(n_2142),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_2203),
.Y(n_2286)
);

BUFx3_ASAP7_75t_L g2287 ( 
.A(n_2203),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2220),
.B(n_2173),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_R g2289 ( 
.A(n_2219),
.B(n_2176),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2231),
.B(n_2169),
.Y(n_2290)
);

NAND2xp33_ASAP7_75t_R g2291 ( 
.A(n_2276),
.B(n_2123),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2251),
.B(n_2163),
.Y(n_2292)
);

CKINVDCx6p67_ASAP7_75t_R g2293 ( 
.A(n_2202),
.Y(n_2293)
);

XNOR2xp5_ASAP7_75t_L g2294 ( 
.A(n_2271),
.B(n_2171),
.Y(n_2294)
);

NAND2xp33_ASAP7_75t_R g2295 ( 
.A(n_2250),
.B(n_2154),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2216),
.B(n_2088),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2222),
.B(n_2129),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2249),
.B(n_2118),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2239),
.B(n_2183),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_R g2300 ( 
.A(n_2236),
.B(n_2187),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2240),
.B(n_2134),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_R g2302 ( 
.A(n_2236),
.B(n_2246),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2270),
.B(n_2208),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2238),
.B(n_2145),
.Y(n_2304)
);

CKINVDCx16_ASAP7_75t_R g2305 ( 
.A(n_2258),
.Y(n_2305)
);

INVxp67_ASAP7_75t_L g2306 ( 
.A(n_2225),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_R g2307 ( 
.A(n_2257),
.B(n_2197),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_R g2308 ( 
.A(n_2267),
.B(n_931),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2228),
.B(n_2185),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2206),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_R g2311 ( 
.A(n_2272),
.B(n_2232),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2252),
.B(n_2135),
.Y(n_2312)
);

BUFx2_ASAP7_75t_L g2313 ( 
.A(n_2218),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2223),
.B(n_2168),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2226),
.B(n_2137),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2204),
.B(n_2180),
.Y(n_2316)
);

CKINVDCx20_ASAP7_75t_R g2317 ( 
.A(n_2209),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_R g2318 ( 
.A(n_2266),
.B(n_933),
.Y(n_2318)
);

NAND2xp33_ASAP7_75t_R g2319 ( 
.A(n_2214),
.B(n_2160),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_R g2320 ( 
.A(n_2265),
.B(n_934),
.Y(n_2320)
);

OR2x6_ASAP7_75t_L g2321 ( 
.A(n_2278),
.B(n_2166),
.Y(n_2321)
);

NAND2x1_ASAP7_75t_L g2322 ( 
.A(n_2235),
.B(n_2152),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2207),
.B(n_2145),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_R g2324 ( 
.A(n_2269),
.B(n_936),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_2213),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2221),
.Y(n_2326)
);

NAND2xp33_ASAP7_75t_SL g2327 ( 
.A(n_2241),
.B(n_2113),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2211),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2328),
.Y(n_2329)
);

INVx2_ASAP7_75t_SL g2330 ( 
.A(n_2286),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2303),
.B(n_2212),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2284),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2310),
.Y(n_2333)
);

INVxp67_ASAP7_75t_SL g2334 ( 
.A(n_2306),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2311),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2283),
.B(n_2244),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2316),
.B(n_2245),
.Y(n_2337)
);

INVxp67_ASAP7_75t_L g2338 ( 
.A(n_2313),
.Y(n_2338)
);

NOR2xp67_ASAP7_75t_L g2339 ( 
.A(n_2296),
.B(n_2224),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2326),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2323),
.Y(n_2341)
);

OR2x2_ASAP7_75t_L g2342 ( 
.A(n_2309),
.B(n_2255),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2290),
.B(n_2256),
.Y(n_2343)
);

AOI22xp33_ASAP7_75t_L g2344 ( 
.A1(n_2327),
.A2(n_2217),
.B1(n_2242),
.B2(n_2254),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2325),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2297),
.B(n_2234),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_2304),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2315),
.A2(n_2264),
.B1(n_2268),
.B2(n_2263),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2314),
.B(n_2227),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2325),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2301),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2292),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2322),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2312),
.Y(n_2354)
);

OAI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2299),
.A2(n_2247),
.B1(n_2215),
.B2(n_2156),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2305),
.B(n_2259),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2298),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_2289),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2294),
.A2(n_2247),
.B1(n_2131),
.B2(n_2116),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2285),
.B(n_2229),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2288),
.B(n_2261),
.Y(n_2361)
);

HB1xp67_ASAP7_75t_L g2362 ( 
.A(n_2319),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2286),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2318),
.B(n_2275),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2287),
.B(n_2277),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_2302),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2321),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2307),
.B(n_2243),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2320),
.B(n_2324),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2321),
.Y(n_2370)
);

OAI222xp33_ASAP7_75t_L g2371 ( 
.A1(n_2317),
.A2(n_2260),
.B1(n_2186),
.B2(n_2273),
.C1(n_2274),
.C2(n_2262),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2308),
.B(n_2181),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2293),
.Y(n_2373)
);

AOI22xp33_ASAP7_75t_L g2374 ( 
.A1(n_2300),
.A2(n_2189),
.B1(n_2210),
.B2(n_2162),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2295),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2291),
.B(n_2248),
.Y(n_2376)
);

BUFx2_ASAP7_75t_L g2377 ( 
.A(n_2351),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2332),
.Y(n_2378)
);

BUFx2_ASAP7_75t_L g2379 ( 
.A(n_2356),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2333),
.Y(n_2380)
);

OR2x2_ASAP7_75t_L g2381 ( 
.A(n_2337),
.B(n_2237),
.Y(n_2381)
);

BUFx3_ASAP7_75t_L g2382 ( 
.A(n_2358),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2329),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2336),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2345),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2340),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2343),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2354),
.B(n_2279),
.Y(n_2388)
);

INVx4_ASAP7_75t_L g2389 ( 
.A(n_2335),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2334),
.Y(n_2390)
);

AO21x2_ASAP7_75t_L g2391 ( 
.A1(n_2375),
.A2(n_2198),
.B(n_2193),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_2361),
.B(n_2281),
.Y(n_2392)
);

INVx5_ASAP7_75t_L g2393 ( 
.A(n_2330),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2341),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2344),
.A2(n_2230),
.B1(n_2282),
.B2(n_2101),
.Y(n_2395)
);

OR2x2_ASAP7_75t_L g2396 ( 
.A(n_2352),
.B(n_2150),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2342),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_2375),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2367),
.B(n_2280),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2349),
.Y(n_2400)
);

OAI33xp33_ASAP7_75t_L g2401 ( 
.A1(n_2357),
.A2(n_68),
.A3(n_70),
.B1(n_66),
.B2(n_67),
.B3(n_69),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2363),
.Y(n_2402)
);

INVx1_ASAP7_75t_SL g2403 ( 
.A(n_2366),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2362),
.Y(n_2404)
);

AOI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2359),
.A2(n_2355),
.B(n_2348),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2347),
.B(n_2376),
.Y(n_2406)
);

AOI211xp5_ASAP7_75t_L g2407 ( 
.A1(n_2369),
.A2(n_2190),
.B(n_2191),
.C(n_2079),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2331),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2350),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2338),
.B(n_2121),
.Y(n_2410)
);

OAI221xp5_ASAP7_75t_L g2411 ( 
.A1(n_2372),
.A2(n_2364),
.B1(n_2339),
.B2(n_2370),
.C(n_2374),
.Y(n_2411)
);

INVx4_ASAP7_75t_L g2412 ( 
.A(n_2365),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2346),
.B(n_2092),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2353),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2360),
.B(n_2103),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2346),
.Y(n_2416)
);

AOI22xp33_ASAP7_75t_SL g2417 ( 
.A1(n_2373),
.A2(n_2120),
.B1(n_2148),
.B2(n_2143),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2371),
.Y(n_2418)
);

AO21x2_ASAP7_75t_L g2419 ( 
.A1(n_2375),
.A2(n_2110),
.B(n_2108),
.Y(n_2419)
);

AND2x4_ASAP7_75t_SL g2420 ( 
.A(n_2368),
.B(n_2128),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2332),
.Y(n_2421)
);

OR2x2_ASAP7_75t_SL g2422 ( 
.A(n_2362),
.B(n_67),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2332),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2352),
.B(n_2102),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2352),
.B(n_68),
.Y(n_2425)
);

OAI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2369),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2332),
.Y(n_2427)
);

AO21x2_ASAP7_75t_L g2428 ( 
.A1(n_2375),
.A2(n_71),
.B(n_73),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2352),
.B(n_73),
.Y(n_2429)
);

NAND2xp33_ASAP7_75t_L g2430 ( 
.A(n_2369),
.B(n_74),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2344),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_2361),
.B(n_937),
.Y(n_2432)
);

OAI31xp33_ASAP7_75t_L g2433 ( 
.A1(n_2359),
.A2(n_77),
.A3(n_75),
.B(n_76),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2333),
.Y(n_2434)
);

INVx4_ASAP7_75t_L g2435 ( 
.A(n_2358),
.Y(n_2435)
);

INVx5_ASAP7_75t_L g2436 ( 
.A(n_2358),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2332),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2330),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2380),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2436),
.Y(n_2440)
);

OR2x2_ASAP7_75t_L g2441 ( 
.A(n_2398),
.B(n_79),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2384),
.B(n_80),
.Y(n_2442)
);

NAND2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2436),
.B(n_938),
.Y(n_2443)
);

INVx2_ASAP7_75t_SL g2444 ( 
.A(n_2393),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2406),
.B(n_82),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_2412),
.Y(n_2446)
);

OR2x2_ASAP7_75t_L g2447 ( 
.A(n_2404),
.B(n_82),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2434),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2386),
.Y(n_2449)
);

AOI21xp33_ASAP7_75t_SL g2450 ( 
.A1(n_2405),
.A2(n_84),
.B(n_85),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2387),
.B(n_84),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2378),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2389),
.B(n_85),
.Y(n_2453)
);

NAND2x1p5_ASAP7_75t_L g2454 ( 
.A(n_2393),
.B(n_941),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2390),
.B(n_86),
.Y(n_2455)
);

BUFx2_ASAP7_75t_SL g2456 ( 
.A(n_2435),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2414),
.Y(n_2457)
);

OAI21xp33_ASAP7_75t_L g2458 ( 
.A1(n_2431),
.A2(n_87),
.B(n_88),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2377),
.B(n_89),
.Y(n_2459)
);

AND2x4_ASAP7_75t_SL g2460 ( 
.A(n_2438),
.B(n_2432),
.Y(n_2460)
);

NOR2x1p5_ASAP7_75t_L g2461 ( 
.A(n_2382),
.B(n_90),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2421),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2423),
.Y(n_2463)
);

INVxp67_ASAP7_75t_L g2464 ( 
.A(n_2409),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2427),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2437),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2394),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2400),
.B(n_93),
.Y(n_2468)
);

OR2x2_ASAP7_75t_L g2469 ( 
.A(n_2381),
.B(n_94),
.Y(n_2469)
);

AND2x4_ASAP7_75t_L g2470 ( 
.A(n_2416),
.B(n_94),
.Y(n_2470)
);

INVxp67_ASAP7_75t_L g2471 ( 
.A(n_2402),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2383),
.B(n_95),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2408),
.B(n_2385),
.Y(n_2473)
);

NAND2xp67_ASAP7_75t_L g2474 ( 
.A(n_2425),
.B(n_95),
.Y(n_2474)
);

INVx1_ASAP7_75t_SL g2475 ( 
.A(n_2403),
.Y(n_2475)
);

INVxp67_ASAP7_75t_L g2476 ( 
.A(n_2411),
.Y(n_2476)
);

NAND3xp33_ASAP7_75t_L g2477 ( 
.A(n_2433),
.B(n_96),
.C(n_97),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2392),
.B(n_96),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2410),
.B(n_98),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2388),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2424),
.B(n_99),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2413),
.B(n_101),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2396),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2415),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2438),
.B(n_102),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2429),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2418),
.B(n_103),
.Y(n_2487)
);

NAND2x1p5_ASAP7_75t_L g2488 ( 
.A(n_2399),
.B(n_942),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2419),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2428),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2391),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2420),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2422),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2395),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2407),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2430),
.B(n_2417),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2401),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2426),
.B(n_104),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2412),
.B(n_104),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2379),
.B(n_105),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2380),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2380),
.Y(n_2502)
);

INVxp67_ASAP7_75t_SL g2503 ( 
.A(n_2404),
.Y(n_2503)
);

OR2x2_ASAP7_75t_L g2504 ( 
.A(n_2397),
.B(n_107),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2379),
.B(n_107),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2398),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2380),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2414),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2380),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2398),
.B(n_110),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2380),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2380),
.Y(n_2512)
);

INVx4_ASAP7_75t_L g2513 ( 
.A(n_2436),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2380),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2397),
.B(n_111),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_2412),
.B(n_113),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2380),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2414),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_2513),
.Y(n_2519)
);

AO221x1_ASAP7_75t_L g2520 ( 
.A1(n_2495),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.C(n_118),
.Y(n_2520)
);

NOR2x1_ASAP7_75t_L g2521 ( 
.A(n_2456),
.B(n_115),
.Y(n_2521)
);

AOI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2496),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_2522)
);

NOR4xp25_ASAP7_75t_SL g2523 ( 
.A(n_2490),
.B(n_125),
.C(n_119),
.D(n_124),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2456),
.Y(n_2524)
);

AO221x2_ASAP7_75t_L g2525 ( 
.A1(n_2477),
.A2(n_128),
.B1(n_130),
.B2(n_127),
.C(n_129),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2439),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2444),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2476),
.B(n_126),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2480),
.B(n_127),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_2475),
.Y(n_2530)
);

CKINVDCx20_ASAP7_75t_R g2531 ( 
.A(n_2460),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2508),
.Y(n_2532)
);

AOI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2494),
.A2(n_2497),
.B1(n_2458),
.B2(n_2498),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2448),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2483),
.B(n_133),
.Y(n_2535)
);

INVx2_ASAP7_75t_SL g2536 ( 
.A(n_2506),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2469),
.B(n_133),
.Y(n_2537)
);

AO221x2_ASAP7_75t_L g2538 ( 
.A1(n_2455),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.C(n_137),
.Y(n_2538)
);

AOI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2487),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2484),
.B(n_140),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2485),
.Y(n_2541)
);

CKINVDCx20_ASAP7_75t_R g2542 ( 
.A(n_2446),
.Y(n_2542)
);

NOR4xp25_ASAP7_75t_SL g2543 ( 
.A(n_2453),
.B(n_145),
.C(n_143),
.D(n_144),
.Y(n_2543)
);

OAI221xp5_ASAP7_75t_L g2544 ( 
.A1(n_2450),
.A2(n_146),
.B1(n_143),
.B2(n_144),
.C(n_147),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2501),
.B(n_149),
.Y(n_2545)
);

OR2x6_ASAP7_75t_L g2546 ( 
.A(n_2443),
.B(n_149),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2502),
.B(n_150),
.Y(n_2547)
);

AOI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2492),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2507),
.B(n_153),
.Y(n_2549)
);

NAND2xp33_ASAP7_75t_SL g2550 ( 
.A(n_2500),
.B(n_154),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2471),
.B(n_154),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2474),
.B(n_2451),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2509),
.B(n_155),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2473),
.Y(n_2554)
);

NAND2xp33_ASAP7_75t_R g2555 ( 
.A(n_2510),
.B(n_155),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2518),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2499),
.Y(n_2557)
);

AO221x2_ASAP7_75t_L g2558 ( 
.A1(n_2472),
.A2(n_160),
.B1(n_163),
.B2(n_159),
.C(n_162),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2511),
.B(n_158),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_R g2560 ( 
.A(n_2505),
.B(n_159),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2486),
.B(n_160),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_SL g2562 ( 
.A(n_2454),
.B(n_2464),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2512),
.Y(n_2563)
);

AO221x2_ASAP7_75t_L g2564 ( 
.A1(n_2467),
.A2(n_165),
.B1(n_168),
.B2(n_164),
.C(n_166),
.Y(n_2564)
);

AO221x2_ASAP7_75t_L g2565 ( 
.A1(n_2514),
.A2(n_168),
.B1(n_170),
.B2(n_166),
.C(n_169),
.Y(n_2565)
);

INVxp67_ASAP7_75t_L g2566 ( 
.A(n_2442),
.Y(n_2566)
);

AO221x2_ASAP7_75t_L g2567 ( 
.A1(n_2517),
.A2(n_170),
.B1(n_165),
.B2(n_169),
.C(n_171),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2452),
.B(n_172),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_2516),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2462),
.B(n_173),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2465),
.B(n_174),
.Y(n_2571)
);

OAI22xp33_ASAP7_75t_L g2572 ( 
.A1(n_2488),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2504),
.B(n_176),
.Y(n_2573)
);

AOI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2479),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2574)
);

AND2x4_ASAP7_75t_SL g2575 ( 
.A(n_2510),
.B(n_180),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2481),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2449),
.B(n_184),
.Y(n_2577)
);

OAI221xp5_ASAP7_75t_L g2578 ( 
.A1(n_2515),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_2578)
);

BUFx2_ASAP7_75t_L g2579 ( 
.A(n_2459),
.Y(n_2579)
);

AO221x2_ASAP7_75t_L g2580 ( 
.A1(n_2491),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_2580)
);

INVx4_ASAP7_75t_L g2581 ( 
.A(n_2478),
.Y(n_2581)
);

INVxp67_ASAP7_75t_L g2582 ( 
.A(n_2441),
.Y(n_2582)
);

OAI221xp5_ASAP7_75t_L g2583 ( 
.A1(n_2447),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.C(n_195),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2463),
.B(n_192),
.Y(n_2584)
);

OAI221xp5_ASAP7_75t_L g2585 ( 
.A1(n_2489),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.C(n_196),
.Y(n_2585)
);

AOI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2482),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2466),
.B(n_197),
.Y(n_2587)
);

NOR2x1_ASAP7_75t_L g2588 ( 
.A(n_2445),
.B(n_199),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2468),
.B(n_201),
.Y(n_2589)
);

A2O1A1Ixp33_ASAP7_75t_L g2590 ( 
.A1(n_2470),
.A2(n_207),
.B(n_215),
.C(n_201),
.Y(n_2590)
);

NAND2xp33_ASAP7_75t_SL g2591 ( 
.A(n_2461),
.B(n_203),
.Y(n_2591)
);

INVxp67_ASAP7_75t_L g2592 ( 
.A(n_2469),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2503),
.B(n_204),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2457),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2503),
.B(n_204),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2506),
.Y(n_2596)
);

CKINVDCx20_ASAP7_75t_R g2597 ( 
.A(n_2460),
.Y(n_2597)
);

CKINVDCx14_ASAP7_75t_R g2598 ( 
.A(n_2486),
.Y(n_2598)
);

INVxp67_ASAP7_75t_SL g2599 ( 
.A(n_2506),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2457),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2503),
.B(n_206),
.Y(n_2601)
);

OAI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2476),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.C(n_210),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2503),
.B(n_208),
.Y(n_2603)
);

OAI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2476),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.C(n_214),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_R g2605 ( 
.A(n_2440),
.B(n_213),
.Y(n_2605)
);

INVxp67_ASAP7_75t_L g2606 ( 
.A(n_2469),
.Y(n_2606)
);

AO221x2_ASAP7_75t_L g2607 ( 
.A1(n_2493),
.A2(n_217),
.B1(n_214),
.B2(n_216),
.C(n_218),
.Y(n_2607)
);

INVx1_ASAP7_75t_SL g2608 ( 
.A(n_2456),
.Y(n_2608)
);

NAND2xp33_ASAP7_75t_SL g2609 ( 
.A(n_2461),
.B(n_218),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2503),
.B(n_219),
.Y(n_2610)
);

AOI22xp5_ASAP7_75t_L g2611 ( 
.A1(n_2496),
.A2(n_223),
.B1(n_219),
.B2(n_220),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2503),
.B(n_220),
.Y(n_2612)
);

OAI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2495),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2613)
);

OAI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2495),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2503),
.B(n_227),
.Y(n_2615)
);

NOR2x1_ASAP7_75t_L g2616 ( 
.A(n_2513),
.B(n_228),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2503),
.B(n_229),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2457),
.Y(n_2618)
);

INVx1_ASAP7_75t_SL g2619 ( 
.A(n_2605),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2524),
.Y(n_2620)
);

INVx1_ASAP7_75t_SL g2621 ( 
.A(n_2542),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2608),
.B(n_230),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2534),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2527),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2554),
.B(n_230),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2579),
.B(n_2598),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2592),
.B(n_232),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2606),
.B(n_2566),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2582),
.B(n_2536),
.Y(n_2629)
);

OR2x2_ASAP7_75t_L g2630 ( 
.A(n_2596),
.B(n_2599),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2618),
.Y(n_2631)
);

INVxp67_ASAP7_75t_L g2632 ( 
.A(n_2521),
.Y(n_2632)
);

INVx1_ASAP7_75t_SL g2633 ( 
.A(n_2530),
.Y(n_2633)
);

CKINVDCx16_ASAP7_75t_R g2634 ( 
.A(n_2555),
.Y(n_2634)
);

HB1xp67_ASAP7_75t_L g2635 ( 
.A(n_2563),
.Y(n_2635)
);

INVx1_ASAP7_75t_SL g2636 ( 
.A(n_2597),
.Y(n_2636)
);

AND3x1_ASAP7_75t_L g2637 ( 
.A(n_2588),
.B(n_233),
.C(n_234),
.Y(n_2637)
);

INVxp67_ASAP7_75t_L g2638 ( 
.A(n_2616),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2532),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2556),
.B(n_2594),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2600),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2584),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2587),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2562),
.B(n_236),
.Y(n_2644)
);

BUFx3_ASAP7_75t_L g2645 ( 
.A(n_2541),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2560),
.Y(n_2646)
);

NAND2x1p5_ASAP7_75t_L g2647 ( 
.A(n_2581),
.B(n_237),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2568),
.Y(n_2648)
);

AND3x1_ASAP7_75t_L g2649 ( 
.A(n_2522),
.B(n_237),
.C(n_238),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2570),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2552),
.B(n_242),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2577),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2571),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2535),
.Y(n_2654)
);

BUFx3_ASAP7_75t_L g2655 ( 
.A(n_2557),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2525),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2551),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2569),
.Y(n_2658)
);

INVx2_ASAP7_75t_SL g2659 ( 
.A(n_2575),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2545),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2547),
.Y(n_2661)
);

CKINVDCx16_ASAP7_75t_R g2662 ( 
.A(n_2591),
.Y(n_2662)
);

AOI22xp33_ASAP7_75t_L g2663 ( 
.A1(n_2607),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2529),
.B(n_248),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2561),
.B(n_249),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2549),
.Y(n_2666)
);

AO22x1_ASAP7_75t_L g2667 ( 
.A1(n_2593),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2607),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2540),
.B(n_254),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2553),
.Y(n_2670)
);

OR2x2_ASAP7_75t_L g2671 ( 
.A(n_2595),
.B(n_254),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2559),
.Y(n_2672)
);

INVx1_ASAP7_75t_SL g2673 ( 
.A(n_2550),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2601),
.Y(n_2674)
);

HB1xp67_ASAP7_75t_L g2675 ( 
.A(n_2617),
.Y(n_2675)
);

OAI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2533),
.A2(n_258),
.B1(n_255),
.B2(n_257),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2546),
.Y(n_2677)
);

OAI221xp5_ASAP7_75t_L g2678 ( 
.A1(n_2611),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.C(n_260),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2603),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2610),
.Y(n_2680)
);

INVx4_ASAP7_75t_L g2681 ( 
.A(n_2546),
.Y(n_2681)
);

NOR2x1_ASAP7_75t_L g2682 ( 
.A(n_2612),
.B(n_261),
.Y(n_2682)
);

INVxp67_ASAP7_75t_L g2683 ( 
.A(n_2528),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2573),
.B(n_262),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2615),
.Y(n_2685)
);

INVx1_ASAP7_75t_SL g2686 ( 
.A(n_2609),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2537),
.B(n_262),
.Y(n_2687)
);

AOI211x1_ASAP7_75t_SL g2688 ( 
.A1(n_2590),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2589),
.Y(n_2689)
);

OR2x2_ASAP7_75t_L g2690 ( 
.A(n_2538),
.B(n_2558),
.Y(n_2690)
);

NAND2x1p5_ASAP7_75t_L g2691 ( 
.A(n_2586),
.B(n_268),
.Y(n_2691)
);

INVx1_ASAP7_75t_SL g2692 ( 
.A(n_2548),
.Y(n_2692)
);

INVx2_ASAP7_75t_SL g2693 ( 
.A(n_2580),
.Y(n_2693)
);

OAI21xp33_ASAP7_75t_L g2694 ( 
.A1(n_2539),
.A2(n_268),
.B(n_269),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2572),
.B(n_270),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2538),
.Y(n_2696)
);

NOR2x1_ASAP7_75t_L g2697 ( 
.A(n_2585),
.B(n_271),
.Y(n_2697)
);

INVx1_ASAP7_75t_SL g2698 ( 
.A(n_2574),
.Y(n_2698)
);

AOI221xp5_ASAP7_75t_L g2699 ( 
.A1(n_2602),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.C(n_275),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2567),
.B(n_278),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2564),
.Y(n_2701)
);

CKINVDCx16_ASAP7_75t_R g2702 ( 
.A(n_2543),
.Y(n_2702)
);

INVx2_ASAP7_75t_SL g2703 ( 
.A(n_2565),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2576),
.Y(n_2704)
);

INVx2_ASAP7_75t_SL g2705 ( 
.A(n_2523),
.Y(n_2705)
);

INVxp67_ASAP7_75t_L g2706 ( 
.A(n_2578),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2614),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2583),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2613),
.B(n_282),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2604),
.Y(n_2710)
);

HB1xp67_ASAP7_75t_L g2711 ( 
.A(n_2544),
.Y(n_2711)
);

INVx1_ASAP7_75t_SL g2712 ( 
.A(n_2605),
.Y(n_2712)
);

OR2x2_ASAP7_75t_L g2713 ( 
.A(n_2592),
.B(n_283),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2526),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2519),
.B(n_285),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2526),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2526),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2519),
.B(n_286),
.Y(n_2718)
);

OR2x2_ASAP7_75t_L g2719 ( 
.A(n_2592),
.B(n_287),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2526),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2519),
.B(n_288),
.Y(n_2721)
);

INVx1_ASAP7_75t_SL g2722 ( 
.A(n_2605),
.Y(n_2722)
);

OR2x2_ASAP7_75t_L g2723 ( 
.A(n_2592),
.B(n_289),
.Y(n_2723)
);

OAI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2598),
.A2(n_292),
.B1(n_289),
.B2(n_290),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2527),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2519),
.B(n_294),
.Y(n_2726)
);

NAND3x1_ASAP7_75t_SL g2727 ( 
.A(n_2521),
.B(n_293),
.C(n_294),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2526),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2519),
.B(n_293),
.Y(n_2729)
);

AND2x4_ASAP7_75t_L g2730 ( 
.A(n_2519),
.B(n_296),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2527),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2527),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2519),
.B(n_297),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2519),
.B(n_298),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2592),
.B(n_299),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2526),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2526),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2552),
.B(n_300),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2519),
.B(n_300),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2526),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2520),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_R g2742 ( 
.A(n_2555),
.B(n_302),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2526),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2525),
.A2(n_305),
.B1(n_301),
.B2(n_303),
.Y(n_2744)
);

NOR2xp33_ASAP7_75t_L g2745 ( 
.A(n_2552),
.B(n_305),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2526),
.Y(n_2746)
);

BUFx3_ASAP7_75t_L g2747 ( 
.A(n_2531),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2526),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2519),
.B(n_307),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2526),
.Y(n_2750)
);

INVxp67_ASAP7_75t_L g2751 ( 
.A(n_2521),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2526),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2592),
.B(n_308),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2519),
.B(n_308),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2526),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2526),
.Y(n_2756)
);

AND2x4_ASAP7_75t_L g2757 ( 
.A(n_2519),
.B(n_310),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2592),
.B(n_309),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2634),
.A2(n_312),
.B1(n_309),
.B2(n_311),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2635),
.Y(n_2760)
);

OAI211xp5_ASAP7_75t_L g2761 ( 
.A1(n_2742),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2693),
.B(n_313),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2632),
.B(n_2751),
.Y(n_2763)
);

XNOR2xp5_ASAP7_75t_L g2764 ( 
.A(n_2637),
.B(n_314),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2711),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2765)
);

AOI211xp5_ASAP7_75t_L g2766 ( 
.A1(n_2676),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_SL g2767 ( 
.A(n_2662),
.B(n_319),
.Y(n_2767)
);

OAI22xp33_ASAP7_75t_L g2768 ( 
.A1(n_2690),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2626),
.B(n_320),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2702),
.A2(n_324),
.B1(n_321),
.B2(n_323),
.Y(n_2770)
);

AOI222xp33_ASAP7_75t_L g2771 ( 
.A1(n_2706),
.A2(n_326),
.B1(n_328),
.B2(n_324),
.C1(n_325),
.C2(n_327),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2623),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2630),
.B(n_330),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2638),
.B(n_331),
.Y(n_2774)
);

OAI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2668),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2775)
);

AOI21xp33_ASAP7_75t_R g2776 ( 
.A1(n_2701),
.A2(n_333),
.B(n_334),
.Y(n_2776)
);

OAI22xp33_ASAP7_75t_L g2777 ( 
.A1(n_2696),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_2777)
);

OAI221xp5_ASAP7_75t_L g2778 ( 
.A1(n_2710),
.A2(n_338),
.B1(n_335),
.B2(n_337),
.C(n_339),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2675),
.B(n_338),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_2619),
.Y(n_2780)
);

INVx1_ASAP7_75t_SL g2781 ( 
.A(n_2712),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2681),
.B(n_339),
.Y(n_2782)
);

OAI21xp33_ASAP7_75t_L g2783 ( 
.A1(n_2697),
.A2(n_340),
.B(n_341),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2707),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2784)
);

OAI21xp33_ASAP7_75t_L g2785 ( 
.A1(n_2663),
.A2(n_342),
.B(n_343),
.Y(n_2785)
);

AOI31xp33_ASAP7_75t_L g2786 ( 
.A1(n_2673),
.A2(n_346),
.A3(n_344),
.B(n_345),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2714),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2716),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2624),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2717),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2720),
.Y(n_2791)
);

AOI221xp5_ASAP7_75t_L g2792 ( 
.A1(n_2708),
.A2(n_2667),
.B1(n_2703),
.B2(n_2649),
.C(n_2698),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2725),
.Y(n_2793)
);

AOI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2699),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2728),
.Y(n_2795)
);

AOI21xp33_ASAP7_75t_L g2796 ( 
.A1(n_2705),
.A2(n_349),
.B(n_351),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2731),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2732),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2736),
.Y(n_2799)
);

AOI22xp33_ASAP7_75t_L g2800 ( 
.A1(n_2704),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_2800)
);

OAI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2644),
.A2(n_355),
.B(n_356),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2695),
.A2(n_357),
.B(n_358),
.Y(n_2802)
);

OAI221xp5_ASAP7_75t_L g2803 ( 
.A1(n_2694),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.C(n_360),
.Y(n_2803)
);

INVxp67_ASAP7_75t_L g2804 ( 
.A(n_2686),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2652),
.B(n_360),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2737),
.Y(n_2806)
);

AOI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2692),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2677),
.B(n_362),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2674),
.B(n_363),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2689),
.B(n_364),
.Y(n_2810)
);

HB1xp67_ASAP7_75t_L g2811 ( 
.A(n_2629),
.Y(n_2811)
);

INVxp67_ASAP7_75t_SL g2812 ( 
.A(n_2645),
.Y(n_2812)
);

AOI322xp5_ASAP7_75t_L g2813 ( 
.A1(n_2700),
.A2(n_370),
.A3(n_369),
.B1(n_367),
.B2(n_365),
.C1(n_366),
.C2(n_368),
.Y(n_2813)
);

OAI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2744),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2679),
.B(n_369),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2740),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2743),
.Y(n_2817)
);

INVxp67_ASAP7_75t_L g2818 ( 
.A(n_2682),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2746),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_R g2820 ( 
.A(n_2658),
.B(n_371),
.Y(n_2820)
);

AOI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2741),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_2821)
);

INVx2_ASAP7_75t_SL g2822 ( 
.A(n_2655),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2748),
.Y(n_2823)
);

AOI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2678),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2750),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2752),
.Y(n_2826)
);

OAI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2656),
.A2(n_378),
.B1(n_375),
.B2(n_377),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2680),
.B(n_378),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2755),
.Y(n_2829)
);

OAI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2651),
.A2(n_379),
.B(n_380),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2685),
.B(n_380),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2756),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2628),
.Y(n_2833)
);

AOI221xp5_ASAP7_75t_L g2834 ( 
.A1(n_2738),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.C(n_384),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2640),
.Y(n_2835)
);

NAND2xp33_ASAP7_75t_L g2836 ( 
.A(n_2646),
.B(n_383),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2745),
.B(n_384),
.C(n_385),
.Y(n_2837)
);

OAI211xp5_ASAP7_75t_L g2838 ( 
.A1(n_2709),
.A2(n_388),
.B(n_385),
.C(n_386),
.Y(n_2838)
);

INVx2_ASAP7_75t_SL g2839 ( 
.A(n_2747),
.Y(n_2839)
);

INVx2_ASAP7_75t_SL g2840 ( 
.A(n_2726),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_SL g2841 ( 
.A1(n_2722),
.A2(n_389),
.B1(n_386),
.B2(n_388),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2691),
.A2(n_392),
.B1(n_389),
.B2(n_390),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2654),
.B(n_393),
.Y(n_2843)
);

OAI21xp33_ASAP7_75t_L g2844 ( 
.A1(n_2642),
.A2(n_393),
.B(n_394),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2631),
.Y(n_2845)
);

NAND2xp33_ASAP7_75t_L g2846 ( 
.A(n_2636),
.B(n_397),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2726),
.Y(n_2847)
);

INVxp67_ASAP7_75t_SL g2848 ( 
.A(n_2647),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2639),
.Y(n_2849)
);

AOI21xp33_ASAP7_75t_L g2850 ( 
.A1(n_2643),
.A2(n_397),
.B(n_398),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2641),
.Y(n_2851)
);

OAI322xp33_ASAP7_75t_L g2852 ( 
.A1(n_2724),
.A2(n_406),
.A3(n_403),
.B1(n_401),
.B2(n_399),
.C1(n_400),
.C2(n_402),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2648),
.Y(n_2853)
);

O2A1O1Ixp33_ASAP7_75t_L g2854 ( 
.A1(n_2683),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_2854)
);

AOI21xp33_ASAP7_75t_SL g2855 ( 
.A1(n_2659),
.A2(n_406),
.B(n_407),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2650),
.Y(n_2856)
);

INVxp67_ASAP7_75t_L g2857 ( 
.A(n_2660),
.Y(n_2857)
);

NAND2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2730),
.B(n_407),
.Y(n_2858)
);

OAI21xp33_ASAP7_75t_L g2859 ( 
.A1(n_2661),
.A2(n_408),
.B(n_409),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2653),
.Y(n_2860)
);

INVx1_ASAP7_75t_SL g2861 ( 
.A(n_2633),
.Y(n_2861)
);

OAI211xp5_ASAP7_75t_L g2862 ( 
.A1(n_2666),
.A2(n_2670),
.B(n_2672),
.C(n_2664),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2657),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2757),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2621),
.B(n_2620),
.Y(n_2865)
);

NOR2xp33_ASAP7_75t_L g2866 ( 
.A(n_2713),
.B(n_411),
.Y(n_2866)
);

OR2x2_ASAP7_75t_L g2867 ( 
.A(n_2719),
.B(n_411),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_SL g2868 ( 
.A1(n_2792),
.A2(n_2688),
.B(n_2684),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2772),
.Y(n_2869)
);

OR2x2_ASAP7_75t_L g2870 ( 
.A(n_2763),
.B(n_2723),
.Y(n_2870)
);

OR2x2_ASAP7_75t_L g2871 ( 
.A(n_2804),
.B(n_2735),
.Y(n_2871)
);

INVx8_ASAP7_75t_L g2872 ( 
.A(n_2808),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2812),
.B(n_2757),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2818),
.B(n_2780),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2781),
.B(n_2622),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_L g2876 ( 
.A(n_2861),
.B(n_2671),
.Y(n_2876)
);

INVx1_ASAP7_75t_SL g2877 ( 
.A(n_2858),
.Y(n_2877)
);

NAND2x1p5_ASAP7_75t_L g2878 ( 
.A(n_2839),
.B(n_2625),
.Y(n_2878)
);

AOI221xp5_ASAP7_75t_L g2879 ( 
.A1(n_2770),
.A2(n_2753),
.B1(n_2758),
.B2(n_2687),
.C(n_2669),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2840),
.B(n_2627),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2822),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2787),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2847),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2788),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_R g2885 ( 
.A(n_2836),
.B(n_2715),
.Y(n_2885)
);

INVx1_ASAP7_75t_SL g2886 ( 
.A(n_2767),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2864),
.Y(n_2887)
);

INVx5_ASAP7_75t_L g2888 ( 
.A(n_2805),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2790),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2865),
.B(n_2665),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2833),
.A2(n_2718),
.B1(n_2729),
.B2(n_2721),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2811),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2848),
.B(n_2733),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2789),
.B(n_2734),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2793),
.B(n_2739),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2797),
.B(n_2798),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2835),
.B(n_2749),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2760),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2791),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2773),
.B(n_2754),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2795),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2769),
.B(n_2727),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2799),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2782),
.B(n_412),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2806),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2765),
.B(n_2843),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2841),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2862),
.B(n_412),
.Y(n_2908)
);

INVxp33_ASAP7_75t_L g2909 ( 
.A(n_2774),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2809),
.B(n_413),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2815),
.B(n_414),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2816),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2831),
.B(n_414),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2817),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2783),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2819),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2823),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2825),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2826),
.Y(n_2919)
);

INVx1_ASAP7_75t_SL g2920 ( 
.A(n_2846),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2829),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_2857),
.B(n_418),
.Y(n_2922)
);

AND2x4_ASAP7_75t_L g2923 ( 
.A(n_2853),
.B(n_418),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2845),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2776),
.B(n_419),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2832),
.Y(n_2926)
);

OAI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2794),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2856),
.B(n_421),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2860),
.B(n_422),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2866),
.B(n_423),
.Y(n_2930)
);

NOR2xp67_ASAP7_75t_SL g2931 ( 
.A(n_2761),
.B(n_426),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2849),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2762),
.Y(n_2933)
);

NAND2x1_ASAP7_75t_L g2934 ( 
.A(n_2851),
.B(n_426),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2779),
.B(n_427),
.Y(n_2935)
);

INVx2_ASAP7_75t_SL g2936 ( 
.A(n_2872),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_2885),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2873),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2892),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2898),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2932),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2869),
.Y(n_2942)
);

HB1xp67_ASAP7_75t_L g2943 ( 
.A(n_2888),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2907),
.B(n_2786),
.Y(n_2944)
);

INVx1_ASAP7_75t_SL g2945 ( 
.A(n_2877),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2882),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2884),
.Y(n_2947)
);

INVx2_ASAP7_75t_SL g2948 ( 
.A(n_2872),
.Y(n_2948)
);

CKINVDCx5p33_ASAP7_75t_R g2949 ( 
.A(n_2874),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2888),
.B(n_2768),
.Y(n_2950)
);

HB1xp67_ASAP7_75t_L g2951 ( 
.A(n_2888),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2889),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2899),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2901),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2903),
.Y(n_2955)
);

INVx3_ASAP7_75t_L g2956 ( 
.A(n_2878),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_2904),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2881),
.Y(n_2958)
);

INVx1_ASAP7_75t_SL g2959 ( 
.A(n_2920),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2905),
.Y(n_2960)
);

INVx8_ASAP7_75t_L g2961 ( 
.A(n_2922),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2909),
.B(n_2828),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2912),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2914),
.Y(n_2964)
);

HB1xp67_ASAP7_75t_L g2965 ( 
.A(n_2934),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2893),
.Y(n_2966)
);

HB1xp67_ASAP7_75t_L g2967 ( 
.A(n_2875),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2916),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2917),
.Y(n_2969)
);

INVx1_ASAP7_75t_SL g2970 ( 
.A(n_2886),
.Y(n_2970)
);

NOR2x1_ASAP7_75t_L g2971 ( 
.A(n_2908),
.B(n_2837),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2918),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2919),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2921),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2926),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2871),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2883),
.Y(n_2977)
);

INVx2_ASAP7_75t_SL g2978 ( 
.A(n_2923),
.Y(n_2978)
);

INVxp33_ASAP7_75t_SL g2979 ( 
.A(n_2876),
.Y(n_2979)
);

INVxp33_ASAP7_75t_L g2980 ( 
.A(n_2890),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2887),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2880),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2902),
.B(n_2764),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2900),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2924),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2928),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2929),
.Y(n_2987)
);

INVxp33_ASAP7_75t_SL g2988 ( 
.A(n_2931),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2896),
.Y(n_2989)
);

INVx2_ASAP7_75t_SL g2990 ( 
.A(n_2897),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2915),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_2933),
.B(n_2810),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2894),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2895),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2870),
.Y(n_2995)
);

CKINVDCx5p33_ASAP7_75t_R g2996 ( 
.A(n_2910),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2935),
.Y(n_2997)
);

CKINVDCx5p33_ASAP7_75t_R g2998 ( 
.A(n_2911),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2913),
.Y(n_2999)
);

NOR2x1_ASAP7_75t_L g3000 ( 
.A(n_2868),
.B(n_2759),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2930),
.Y(n_3001)
);

INVxp33_ASAP7_75t_SL g3002 ( 
.A(n_2925),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2906),
.Y(n_3003)
);

INVx2_ASAP7_75t_SL g3004 ( 
.A(n_2927),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2891),
.Y(n_3005)
);

BUFx4f_ASAP7_75t_SL g3006 ( 
.A(n_2879),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2892),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2945),
.B(n_2855),
.Y(n_3008)
);

NOR3xp33_ASAP7_75t_L g3009 ( 
.A(n_3000),
.B(n_2778),
.C(n_2796),
.Y(n_3009)
);

AOI21xp5_ASAP7_75t_L g3010 ( 
.A1(n_2988),
.A2(n_2830),
.B(n_2802),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2966),
.B(n_2784),
.Y(n_3011)
);

NOR3x1_ASAP7_75t_L g3012 ( 
.A(n_2944),
.B(n_2838),
.C(n_2801),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_3006),
.A2(n_2775),
.B1(n_2785),
.B2(n_2824),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2991),
.A2(n_2766),
.B1(n_2807),
.B2(n_2821),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2959),
.B(n_2813),
.Y(n_3015)
);

NAND4xp25_ASAP7_75t_L g3016 ( 
.A(n_2970),
.B(n_2771),
.C(n_2834),
.D(n_2854),
.Y(n_3016)
);

OAI221xp5_ASAP7_75t_L g3017 ( 
.A1(n_2971),
.A2(n_2859),
.B1(n_2844),
.B2(n_2803),
.C(n_2800),
.Y(n_3017)
);

NAND3xp33_ASAP7_75t_L g3018 ( 
.A(n_2950),
.B(n_2951),
.C(n_2943),
.Y(n_3018)
);

AO22x2_ASAP7_75t_L g3019 ( 
.A1(n_3003),
.A2(n_2867),
.B1(n_2842),
.B2(n_2827),
.Y(n_3019)
);

NAND3xp33_ASAP7_75t_L g3020 ( 
.A(n_2965),
.B(n_2850),
.C(n_2863),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2979),
.B(n_2814),
.Y(n_3021)
);

OAI21xp33_ASAP7_75t_L g3022 ( 
.A1(n_2980),
.A2(n_2820),
.B(n_2777),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2939),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_SL g3024 ( 
.A(n_2949),
.B(n_2852),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2956),
.B(n_427),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_3007),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2940),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_SL g3028 ( 
.A1(n_2937),
.A2(n_428),
.B(n_430),
.Y(n_3028)
);

NOR3xp33_ASAP7_75t_SL g3029 ( 
.A(n_2957),
.B(n_432),
.C(n_433),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2983),
.A2(n_432),
.B(n_433),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2996),
.B(n_434),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2936),
.B(n_2948),
.Y(n_3032)
);

NOR4xp25_ASAP7_75t_L g3033 ( 
.A(n_3004),
.B(n_437),
.C(n_434),
.D(n_436),
.Y(n_3033)
);

NAND5xp2_ASAP7_75t_L g3034 ( 
.A(n_2995),
.B(n_438),
.C(n_436),
.D(n_437),
.E(n_439),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2984),
.Y(n_3035)
);

NAND4xp75_ASAP7_75t_L g3036 ( 
.A(n_2976),
.B(n_440),
.C(n_438),
.D(n_439),
.Y(n_3036)
);

AOI311xp33_ASAP7_75t_L g3037 ( 
.A1(n_2982),
.A2(n_442),
.A3(n_440),
.B(n_441),
.C(n_443),
.Y(n_3037)
);

NAND4xp25_ASAP7_75t_L g3038 ( 
.A(n_2938),
.B(n_446),
.C(n_444),
.D(n_445),
.Y(n_3038)
);

NAND3xp33_ASAP7_75t_L g3039 ( 
.A(n_2967),
.B(n_446),
.C(n_447),
.Y(n_3039)
);

NOR2xp33_ASAP7_75t_L g3040 ( 
.A(n_3002),
.B(n_447),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2962),
.A2(n_448),
.B(n_449),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2998),
.B(n_448),
.Y(n_3042)
);

OAI221xp5_ASAP7_75t_L g3043 ( 
.A1(n_3005),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.C(n_452),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2978),
.B(n_452),
.Y(n_3044)
);

NAND4xp75_ASAP7_75t_L g3045 ( 
.A(n_2977),
.B(n_455),
.C(n_453),
.D(n_454),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2961),
.B(n_3001),
.Y(n_3046)
);

NOR2xp33_ASAP7_75t_L g3047 ( 
.A(n_2961),
.B(n_453),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2990),
.B(n_457),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2997),
.B(n_2999),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2958),
.B(n_457),
.Y(n_3050)
);

AOI211xp5_ASAP7_75t_L g3051 ( 
.A1(n_2992),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_3051)
);

NOR3xp33_ASAP7_75t_L g3052 ( 
.A(n_2986),
.B(n_461),
.C(n_462),
.Y(n_3052)
);

AND4x1_ASAP7_75t_L g3053 ( 
.A(n_2987),
.B(n_464),
.C(n_461),
.D(n_463),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2989),
.B(n_465),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2993),
.A2(n_465),
.B(n_466),
.Y(n_3055)
);

NOR3x1_ASAP7_75t_L g3056 ( 
.A(n_2994),
.B(n_467),
.C(n_468),
.Y(n_3056)
);

NAND3xp33_ASAP7_75t_L g3057 ( 
.A(n_2981),
.B(n_2985),
.C(n_2941),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2942),
.A2(n_470),
.B(n_472),
.Y(n_3058)
);

AOI221xp5_ASAP7_75t_L g3059 ( 
.A1(n_3018),
.A2(n_2952),
.B1(n_2953),
.B2(n_2947),
.C(n_2946),
.Y(n_3059)
);

AOI21xp33_ASAP7_75t_L g3060 ( 
.A1(n_3046),
.A2(n_2955),
.B(n_2954),
.Y(n_3060)
);

OAI221xp5_ASAP7_75t_SL g3061 ( 
.A1(n_3013),
.A2(n_2964),
.B1(n_2968),
.B2(n_2963),
.C(n_2960),
.Y(n_3061)
);

NOR2xp33_ASAP7_75t_L g3062 ( 
.A(n_3022),
.B(n_2969),
.Y(n_3062)
);

AOI221xp5_ASAP7_75t_L g3063 ( 
.A1(n_3019),
.A2(n_2974),
.B1(n_2975),
.B2(n_2973),
.C(n_2972),
.Y(n_3063)
);

OAI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_3020),
.A2(n_3010),
.B(n_3024),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_3030),
.A2(n_3017),
.B(n_3014),
.Y(n_3065)
);

NAND4xp25_ASAP7_75t_SL g3066 ( 
.A(n_3015),
.B(n_475),
.C(n_473),
.D(n_474),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_3032),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_3033),
.B(n_475),
.Y(n_3068)
);

NAND4xp25_ASAP7_75t_SL g3069 ( 
.A(n_3028),
.B(n_478),
.C(n_476),
.D(n_477),
.Y(n_3069)
);

AOI31xp33_ASAP7_75t_L g3070 ( 
.A1(n_3008),
.A2(n_479),
.A3(n_476),
.B(n_477),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_3047),
.B(n_480),
.Y(n_3071)
);

AOI221xp5_ASAP7_75t_L g3072 ( 
.A1(n_3019),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.C(n_483),
.Y(n_3072)
);

BUFx6f_ASAP7_75t_L g3073 ( 
.A(n_3025),
.Y(n_3073)
);

AOI221x1_ASAP7_75t_L g3074 ( 
.A1(n_3052),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.C(n_484),
.Y(n_3074)
);

AO22x2_ASAP7_75t_L g3075 ( 
.A1(n_3057),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_3075)
);

NAND4xp75_ASAP7_75t_L g3076 ( 
.A(n_3012),
.B(n_3056),
.C(n_3026),
.D(n_3023),
.Y(n_3076)
);

AOI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_3016),
.A2(n_3021),
.B1(n_3035),
.B2(n_3011),
.Y(n_3077)
);

AO22x2_ASAP7_75t_L g3078 ( 
.A1(n_3027),
.A2(n_488),
.B1(n_486),
.B2(n_487),
.Y(n_3078)
);

OAI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_3029),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_3079)
);

NAND5xp2_ASAP7_75t_SL g3080 ( 
.A(n_3043),
.B(n_492),
.C(n_490),
.D(n_491),
.E(n_493),
.Y(n_3080)
);

BUFx6f_ASAP7_75t_L g3081 ( 
.A(n_3050),
.Y(n_3081)
);

NAND3xp33_ASAP7_75t_SL g3082 ( 
.A(n_3051),
.B(n_494),
.C(n_496),
.Y(n_3082)
);

AOI211xp5_ASAP7_75t_SL g3083 ( 
.A1(n_3049),
.A2(n_500),
.B(n_497),
.C(n_499),
.Y(n_3083)
);

AOI221xp5_ASAP7_75t_L g3084 ( 
.A1(n_3039),
.A2(n_501),
.B1(n_497),
.B2(n_500),
.C(n_502),
.Y(n_3084)
);

A2O1A1Ixp33_ASAP7_75t_L g3085 ( 
.A1(n_3041),
.A2(n_503),
.B(n_501),
.C(n_502),
.Y(n_3085)
);

AOI22xp5_ASAP7_75t_L g3086 ( 
.A1(n_3040),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_3086)
);

AOI22xp33_ASAP7_75t_SL g3087 ( 
.A1(n_3058),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3087)
);

A2O1A1Ixp33_ASAP7_75t_L g3088 ( 
.A1(n_3055),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_3036),
.A2(n_510),
.B(n_511),
.Y(n_3089)
);

NOR4xp25_ASAP7_75t_SL g3090 ( 
.A(n_3048),
.B(n_515),
.C(n_512),
.D(n_514),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_SL g3091 ( 
.A(n_3045),
.B(n_514),
.Y(n_3091)
);

NAND4xp25_ASAP7_75t_SL g3092 ( 
.A(n_3054),
.B(n_521),
.C(n_516),
.D(n_520),
.Y(n_3092)
);

CKINVDCx5p33_ASAP7_75t_R g3093 ( 
.A(n_3042),
.Y(n_3093)
);

NOR2x1_ASAP7_75t_L g3094 ( 
.A(n_3038),
.B(n_520),
.Y(n_3094)
);

OAI22xp5_ASAP7_75t_L g3095 ( 
.A1(n_3031),
.A2(n_525),
.B1(n_522),
.B2(n_523),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3053),
.B(n_527),
.Y(n_3096)
);

AND2x4_ASAP7_75t_L g3097 ( 
.A(n_3044),
.B(n_527),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_3037),
.A2(n_531),
.B1(n_528),
.B2(n_530),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_3034),
.A2(n_531),
.B(n_532),
.Y(n_3099)
);

AOI211xp5_ASAP7_75t_L g3100 ( 
.A1(n_3009),
.A2(n_535),
.B(n_533),
.C(n_534),
.Y(n_3100)
);

AOI22xp5_ASAP7_75t_L g3101 ( 
.A1(n_3009),
.A2(n_537),
.B1(n_534),
.B2(n_536),
.Y(n_3101)
);

AOI221xp5_ASAP7_75t_L g3102 ( 
.A1(n_3009),
.A2(n_539),
.B1(n_536),
.B2(n_538),
.C(n_541),
.Y(n_3102)
);

AO22x1_ASAP7_75t_L g3103 ( 
.A1(n_3009),
.A2(n_541),
.B1(n_538),
.B2(n_539),
.Y(n_3103)
);

AOI221xp5_ASAP7_75t_L g3104 ( 
.A1(n_3009),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.C(n_545),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_3073),
.Y(n_3105)
);

NOR4xp75_ASAP7_75t_L g3106 ( 
.A(n_3076),
.B(n_546),
.C(n_543),
.D(n_545),
.Y(n_3106)
);

XNOR2xp5_ASAP7_75t_L g3107 ( 
.A(n_3077),
.B(n_547),
.Y(n_3107)
);

AO211x2_ASAP7_75t_L g3108 ( 
.A1(n_3064),
.A2(n_550),
.B(n_548),
.C(n_549),
.Y(n_3108)
);

NOR2x1_ASAP7_75t_L g3109 ( 
.A(n_3069),
.B(n_548),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_3067),
.B(n_549),
.Y(n_3110)
);

NOR2x1_ASAP7_75t_L g3111 ( 
.A(n_3066),
.B(n_3092),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3073),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_3103),
.B(n_554),
.Y(n_3113)
);

NAND2xp33_ASAP7_75t_L g3114 ( 
.A(n_3093),
.B(n_556),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_3081),
.Y(n_3115)
);

OAI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_3098),
.A2(n_3101),
.B1(n_3065),
.B2(n_3068),
.Y(n_3116)
);

AOI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_3091),
.A2(n_3062),
.B1(n_3094),
.B2(n_3072),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_3081),
.B(n_558),
.Y(n_3118)
);

AND2x4_ASAP7_75t_L g3119 ( 
.A(n_3089),
.B(n_558),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_3078),
.Y(n_3120)
);

AOI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_3082),
.A2(n_562),
.B1(n_559),
.B2(n_561),
.Y(n_3121)
);

INVx1_ASAP7_75t_SL g3122 ( 
.A(n_3096),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_3097),
.Y(n_3123)
);

NAND2xp33_ASAP7_75t_L g3124 ( 
.A(n_3085),
.B(n_562),
.Y(n_3124)
);

INVxp33_ASAP7_75t_L g3125 ( 
.A(n_3079),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_3075),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3083),
.B(n_563),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_R g3128 ( 
.A(n_3114),
.B(n_3080),
.Y(n_3128)
);

NAND2xp33_ASAP7_75t_R g3129 ( 
.A(n_3119),
.B(n_3090),
.Y(n_3129)
);

NAND2xp33_ASAP7_75t_SL g3130 ( 
.A(n_3113),
.B(n_3071),
.Y(n_3130)
);

NOR2xp33_ASAP7_75t_R g3131 ( 
.A(n_3124),
.B(n_3070),
.Y(n_3131)
);

NAND2xp33_ASAP7_75t_SL g3132 ( 
.A(n_3120),
.B(n_3095),
.Y(n_3132)
);

NAND3xp33_ASAP7_75t_SL g3133 ( 
.A(n_3106),
.B(n_3100),
.C(n_3102),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_R g3134 ( 
.A(n_3107),
.B(n_3074),
.Y(n_3134)
);

NAND2xp33_ASAP7_75t_SL g3135 ( 
.A(n_3126),
.B(n_3061),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_R g3136 ( 
.A(n_3127),
.B(n_3087),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_3109),
.B(n_3063),
.Y(n_3137)
);

NOR3xp33_ASAP7_75t_SL g3138 ( 
.A(n_3116),
.B(n_3060),
.C(n_3059),
.Y(n_3138)
);

AOI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_3135),
.A2(n_3111),
.B1(n_3117),
.B2(n_3112),
.Y(n_3139)
);

CKINVDCx20_ASAP7_75t_R g3140 ( 
.A(n_3132),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3137),
.Y(n_3141)
);

OAI22xp5_ASAP7_75t_SL g3142 ( 
.A1(n_3140),
.A2(n_3122),
.B1(n_3115),
.B2(n_3105),
.Y(n_3142)
);

AOI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_3141),
.A2(n_3129),
.B1(n_3133),
.B2(n_3130),
.Y(n_3143)
);

INVxp67_ASAP7_75t_L g3144 ( 
.A(n_3142),
.Y(n_3144)
);

OAI21x1_ASAP7_75t_L g3145 ( 
.A1(n_3143),
.A2(n_3139),
.B(n_3123),
.Y(n_3145)
);

AOI31xp33_ASAP7_75t_L g3146 ( 
.A1(n_3144),
.A2(n_3125),
.A3(n_3118),
.B(n_3110),
.Y(n_3146)
);

AOI31xp33_ASAP7_75t_L g3147 ( 
.A1(n_3145),
.A2(n_3104),
.A3(n_3121),
.B(n_3084),
.Y(n_3147)
);

XOR2xp5_ASAP7_75t_L g3148 ( 
.A(n_3146),
.B(n_3086),
.Y(n_3148)
);

OAI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_3147),
.A2(n_3138),
.B(n_3088),
.Y(n_3149)
);

A2O1A1Ixp33_ASAP7_75t_SL g3150 ( 
.A1(n_3149),
.A2(n_3099),
.B(n_3134),
.C(n_3136),
.Y(n_3150)
);

AOI222xp33_ASAP7_75t_SL g3151 ( 
.A1(n_3148),
.A2(n_3131),
.B1(n_3128),
.B2(n_3108),
.C1(n_568),
.C2(n_569),
.Y(n_3151)
);

INVxp67_ASAP7_75t_SL g3152 ( 
.A(n_3150),
.Y(n_3152)
);

OAI221xp5_ASAP7_75t_R g3153 ( 
.A1(n_3152),
.A2(n_3151),
.B1(n_567),
.B2(n_565),
.C(n_566),
.Y(n_3153)
);

AOI211xp5_ASAP7_75t_L g3154 ( 
.A1(n_3153),
.A2(n_575),
.B(n_573),
.C(n_574),
.Y(n_3154)
);


endmodule