module fake_jpeg_17474_n_355 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_355);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_22),
.Y(n_61)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_31),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_61),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_25),
.B(n_30),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_30),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_36),
.B1(n_40),
.B2(n_34),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_30),
.B1(n_34),
.B2(n_40),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_66),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_36),
.B1(n_34),
.B2(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_70),
.B1(n_62),
.B2(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_104),
.Y(n_126)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_32),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_52),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_25),
.B(n_24),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_73),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_70),
.B1(n_85),
.B2(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_33),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_35),
.B(n_32),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_34),
.B1(n_29),
.B2(n_36),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_107),
.B1(n_92),
.B2(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_123),
.B1(n_128),
.B2(n_134),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_135),
.B(n_81),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_82),
.B1(n_71),
.B2(n_62),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_40),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_148),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_68),
.B1(n_67),
.B2(n_51),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_84),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_52),
.C(n_50),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_69),
.B1(n_44),
.B2(n_41),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_31),
.B1(n_37),
.B2(n_29),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_29),
.B1(n_37),
.B2(n_22),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_145),
.B1(n_147),
.B2(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_139),
.Y(n_168)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_125),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_47),
.B1(n_79),
.B2(n_37),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_89),
.A2(n_39),
.A3(n_27),
.B1(n_23),
.B2(n_78),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_158),
.Y(n_187)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_170),
.B1(n_89),
.B2(n_142),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_138),
.B(n_133),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_121),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_147),
.B(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_177),
.B(n_191),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_119),
.B1(n_123),
.B2(n_146),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_179),
.B1(n_164),
.B2(n_115),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_118),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_166),
.B1(n_161),
.B2(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_156),
.B1(n_167),
.B2(n_168),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_146),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_194),
.C(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_129),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_147),
.B(n_88),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_134),
.C(n_128),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_145),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_156),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_173),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_214),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_208),
.B1(n_220),
.B2(n_178),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_158),
.B(n_155),
.C(n_147),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_207),
.B(n_176),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_216),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_157),
.B1(n_154),
.B2(n_152),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_101),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_213),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_98),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_150),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_98),
.B1(n_171),
.B2(n_150),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_180),
.B1(n_178),
.B2(n_195),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_140),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_175),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_227),
.B(n_237),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_180),
.B1(n_193),
.B2(n_192),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_238),
.B1(n_245),
.B2(n_81),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_242),
.B1(n_249),
.B2(n_245),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_240),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_191),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_207),
.A2(n_180),
.B1(n_193),
.B2(n_192),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_188),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_177),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_244),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_194),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_246),
.B(n_248),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_178),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_201),
.A2(n_207),
.B(n_206),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_176),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_163),
.B(n_106),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_266),
.B1(n_271),
.B2(n_241),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_210),
.B1(n_218),
.B2(n_200),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_253),
.A2(n_258),
.B1(n_262),
.B2(n_39),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_218),
.B1(n_208),
.B2(n_217),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_215),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_270),
.C(n_227),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_215),
.B(n_213),
.C(n_163),
.D(n_24),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_225),
.C(n_248),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_171),
.B1(n_163),
.B2(n_87),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_27),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_231),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_258),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_27),
.B1(n_39),
.B2(n_14),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_237),
.B(n_23),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_23),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_106),
.C(n_108),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_13),
.B(n_17),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_274),
.B1(n_275),
.B2(n_281),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_279),
.C(n_282),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_239),
.B1(n_230),
.B2(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_230),
.B1(n_247),
.B2(n_225),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_243),
.C(n_109),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_25),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_289),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_264),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_39),
.B1(n_27),
.B2(n_10),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_25),
.C(n_26),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_250),
.C(n_253),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_6),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_257),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_306),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_280),
.B1(n_285),
.B2(n_287),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_7),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_26),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_250),
.B(n_254),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_10),
.B1(n_16),
.B2(n_14),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_261),
.B(n_269),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_9),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_307),
.A2(n_309),
.B1(n_4),
.B2(n_5),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_310),
.B(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_25),
.C(n_1),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_7),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_306),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_25),
.C(n_1),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_320),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_6),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_4),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_291),
.B(n_293),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_331),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_318),
.Y(n_335)
);

XOR2x1_ASAP7_75t_SL g328 ( 
.A(n_308),
.B(n_298),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_304),
.B(n_295),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_333),
.A2(n_325),
.B1(n_323),
.B2(n_328),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_318),
.C(n_5),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_337),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_339),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_4),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_340),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_326),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_5),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_338),
.Y(n_349)
);

AOI322xp5_ASAP7_75t_L g344 ( 
.A1(n_336),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_11),
.C1(n_26),
.C2(n_332),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_342),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_332),
.A2(n_11),
.B(n_26),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_348),
.A2(n_349),
.B(n_341),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_347),
.B(n_346),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_344),
.B(n_11),
.C(n_26),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_0),
.B(n_3),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_353),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);


endmodule