module fake_jpeg_12104_n_582 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_582);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_582;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_64),
.B(n_98),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_74),
.B1(n_30),
.B2(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_28),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g126 ( 
.A(n_81),
.Y(n_126)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_33),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_103),
.B(n_104),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_21),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_107),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_52),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_53),
.B1(n_24),
.B2(n_25),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_131),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_112),
.A2(n_165),
.B1(n_172),
.B2(n_84),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_37),
.B1(n_25),
.B2(n_21),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_115),
.B(n_0),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_53),
.B1(n_24),
.B2(n_37),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_73),
.B1(n_69),
.B2(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_36),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_0),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_56),
.A2(n_37),
.B1(n_21),
.B2(n_31),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_141),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_54),
.A2(n_53),
.B1(n_29),
.B2(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_166),
.B1(n_79),
.B2(n_78),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_83),
.A2(n_51),
.B(n_23),
.C(n_107),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_159),
.Y(n_207)
);

OR2x2_ASAP7_75t_SL g159 ( 
.A(n_63),
.B(n_49),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_92),
.A2(n_31),
.B1(n_29),
.B2(n_49),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_163),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_57),
.A2(n_29),
.B1(n_36),
.B2(n_26),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_66),
.A2(n_51),
.B1(n_23),
.B2(n_30),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_70),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_172)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_113),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_175),
.B(n_184),
.Y(n_289)
);

AO22x1_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_81),
.B1(n_76),
.B2(n_103),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_215),
.Y(n_243)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_181),
.Y(n_265)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_130),
.B(n_102),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_185),
.B(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_188),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_75),
.B1(n_99),
.B2(n_91),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_193),
.Y(n_287)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_135),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_195),
.B(n_211),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_196),
.Y(n_275)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_197),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_132),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g271 ( 
.A(n_198),
.Y(n_271)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_141),
.A2(n_101),
.B1(n_90),
.B2(n_86),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_201),
.A2(n_213),
.B1(n_171),
.B2(n_167),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_202),
.A2(n_168),
.B1(n_155),
.B2(n_146),
.Y(n_259)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_13),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_209),
.A2(n_218),
.B1(n_221),
.B2(n_223),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_77),
.B1(n_62),
.B2(n_61),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_145),
.B1(n_111),
.B2(n_117),
.Y(n_246)
);

AOI32xp33_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_60),
.A3(n_8),
.B1(n_11),
.B2(n_19),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_163),
.A2(n_18),
.B1(n_16),
.B2(n_14),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_125),
.B(n_18),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_120),
.B(n_16),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_147),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_216),
.Y(n_258)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_132),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_219),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_220),
.B(n_222),
.Y(n_283)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_252)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_227),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_234),
.Y(n_273)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_138),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_157),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_235),
.B(n_236),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_166),
.B(n_148),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_237),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_246),
.A2(n_259),
.B1(n_267),
.B2(n_268),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_248),
.A2(n_257),
.B1(n_269),
.B2(n_279),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_168),
.B(n_126),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_251),
.A2(n_264),
.B(n_266),
.C(n_231),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_146),
.B1(n_129),
.B2(n_139),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_189),
.A2(n_126),
.B(n_152),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_202),
.B(n_201),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_177),
.A2(n_139),
.B1(n_129),
.B2(n_151),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_177),
.A2(n_170),
.B1(n_152),
.B2(n_151),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_226),
.A2(n_170),
.B1(n_127),
.B2(n_126),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_226),
.A2(n_127),
.B1(n_176),
.B2(n_193),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_286),
.B1(n_191),
.B2(n_236),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_203),
.B(n_0),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_285),
.C(n_218),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_208),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_182),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_280),
.A2(n_292),
.B1(n_1),
.B2(n_3),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_216),
.B(n_14),
.C(n_12),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_178),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_187),
.A2(n_12),
.B1(n_11),
.B2(n_8),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_293),
.B(n_323),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_294),
.B(n_301),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_230),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_295),
.Y(n_378)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_219),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_297),
.B(n_303),
.C(n_315),
.Y(n_374)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_229),
.C(n_221),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_300),
.B(n_320),
.C(n_326),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_192),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_243),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_304),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_237),
.B(n_194),
.C(n_174),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_217),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_307),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_240),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_309),
.B(n_316),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_241),
.A2(n_205),
.B1(n_225),
.B2(n_188),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_312),
.A2(n_319),
.B(n_247),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_232),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_313),
.B(n_342),
.Y(n_379)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_291),
.C(n_244),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_258),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_317),
.A2(n_300),
.B(n_308),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_327),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_241),
.A2(n_183),
.B1(n_197),
.B2(n_179),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_SL g320 ( 
.A(n_283),
.B(n_12),
.C(n_198),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_321),
.A2(n_336),
.B1(n_338),
.B2(n_292),
.Y(n_368)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_284),
.B(n_209),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_325),
.A2(n_278),
.B1(n_262),
.B2(n_287),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_1),
.C(n_3),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_284),
.B(n_3),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_245),
.Y(n_329)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_4),
.C(n_5),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_285),
.Y(n_352)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_334),
.Y(n_364)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_343),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_250),
.A2(n_259),
.B1(n_267),
.B2(n_268),
.Y(n_336)
);

INVx13_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_337),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_250),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_266),
.A2(n_4),
.B(n_5),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_320),
.B(n_306),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_265),
.B(n_4),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_340),
.B(n_341),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_275),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_247),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_308),
.A2(n_248),
.B1(n_257),
.B2(n_246),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_368),
.B1(n_384),
.B2(n_286),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_346),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_352),
.B(n_253),
.Y(n_420)
);

AO22x1_ASAP7_75t_SL g353 ( 
.A1(n_296),
.A2(n_255),
.B1(n_274),
.B2(n_272),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_383),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_313),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_372),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_306),
.A2(n_273),
.B(n_238),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_359),
.A2(n_366),
.B(n_279),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_297),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_382),
.C(n_317),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_304),
.B1(n_298),
.B2(n_303),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_362),
.A2(n_371),
.B1(n_318),
.B2(n_326),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_272),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_365),
.B(n_367),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_294),
.B(n_293),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_337),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_299),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_239),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_301),
.B(n_275),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_263),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_336),
.A2(n_321),
.B1(n_317),
.B2(n_338),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_389),
.A2(n_396),
.B1(n_406),
.B2(n_368),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_305),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_394),
.C(n_399),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_391),
.B(n_388),
.Y(n_442)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_317),
.C(n_263),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_395),
.B(n_409),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_362),
.A2(n_317),
.B1(n_330),
.B2(n_325),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_384),
.A2(n_331),
.B1(n_334),
.B2(n_342),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_398),
.A2(n_411),
.B1(n_359),
.B2(n_349),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_261),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_261),
.C(n_262),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_403),
.C(n_404),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_274),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_255),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_358),
.A2(n_322),
.B1(n_311),
.B2(n_280),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_407),
.Y(n_444)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_379),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_379),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_410),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_373),
.Y(n_438)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_258),
.C(n_239),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_418),
.C(n_422),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

AOI21xp33_ASAP7_75t_L g416 ( 
.A1(n_370),
.A2(n_310),
.B(n_271),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_416),
.A2(n_372),
.B1(n_347),
.B2(n_364),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_351),
.B(n_254),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_424),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_254),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_425),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_383),
.B(n_271),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_427),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_355),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_429),
.A2(n_440),
.B1(n_450),
.B2(n_452),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_455),
.B1(n_419),
.B2(n_405),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_382),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_433),
.B(n_442),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_436),
.A2(n_443),
.B1(n_456),
.B2(n_406),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_397),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_392),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_396),
.A2(n_344),
.B1(n_355),
.B2(n_378),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_411),
.A2(n_346),
.B1(n_345),
.B2(n_388),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_390),
.B(n_352),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_449),
.C(n_459),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_345),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_426),
.A2(n_376),
.B1(n_387),
.B2(n_380),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_389),
.A2(n_387),
.B1(n_381),
.B2(n_380),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_350),
.B1(n_347),
.B2(n_369),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_412),
.A2(n_423),
.B1(n_398),
.B2(n_401),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_400),
.B(n_401),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_457),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_381),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_458),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_385),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_422),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_464),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_465),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_418),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_466),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_394),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_467),
.B(n_475),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_468),
.B(n_479),
.Y(n_514)
);

XNOR2x1_ASAP7_75t_SL g469 ( 
.A(n_428),
.B(n_391),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_433),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_402),
.C(n_414),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_472),
.C(n_484),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_404),
.C(n_403),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_408),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_477),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_474),
.A2(n_479),
.B1(n_486),
.B2(n_487),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_424),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_445),
.B(n_356),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_478),
.B(n_490),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_436),
.A2(n_417),
.B1(n_407),
.B2(n_350),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_429),
.A2(n_417),
.B1(n_385),
.B2(n_375),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_480),
.A2(n_438),
.B1(n_430),
.B2(n_451),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_457),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_483),
.B(n_481),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_369),
.C(n_363),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_457),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_485),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_456),
.A2(n_363),
.B1(n_353),
.B2(n_307),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_443),
.A2(n_438),
.B1(n_435),
.B2(n_461),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_353),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_428),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_287),
.C(n_249),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_249),
.C(n_242),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_441),
.B(n_377),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_496),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_440),
.B1(n_452),
.B2(n_432),
.Y(n_495)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_449),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_487),
.A2(n_435),
.B1(n_450),
.B2(n_430),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_497),
.A2(n_512),
.B1(n_514),
.B2(n_310),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_454),
.Y(n_498)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_499),
.A2(n_485),
.B1(n_484),
.B2(n_466),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

AOI21xp33_ASAP7_75t_L g502 ( 
.A1(n_462),
.A2(n_455),
.B(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_488),
.Y(n_521)
);

XOR2x2_ASAP7_75t_L g507 ( 
.A(n_475),
.B(n_447),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_509),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_463),
.B(n_472),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_469),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_486),
.A2(n_444),
.B1(n_453),
.B2(n_377),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_489),
.C(n_470),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_516),
.B(n_525),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_521),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_505),
.B(n_463),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_510),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_SL g520 ( 
.A1(n_491),
.A2(n_462),
.B(n_471),
.C(n_473),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g537 ( 
.A1(n_520),
.A2(n_514),
.B(n_498),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_523),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_476),
.C(n_471),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_533),
.C(n_501),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_480),
.Y(n_526)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_526),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_499),
.A2(n_464),
.B1(n_310),
.B2(n_242),
.Y(n_528)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_528),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_530),
.A2(n_512),
.B(n_492),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_253),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_513),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_282),
.C(n_6),
.Y(n_533)
);

AOI31xp33_ASAP7_75t_L g550 ( 
.A1(n_535),
.A2(n_541),
.A3(n_546),
.B(n_529),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_500),
.Y(n_536)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_536),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_539),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_497),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_538),
.A2(n_520),
.B1(n_528),
.B2(n_492),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_503),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_548),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_530),
.A2(n_514),
.B(n_491),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_549),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_508),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_516),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_550),
.A2(n_557),
.B1(n_520),
.B2(n_507),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_543),
.B(n_518),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_553),
.B(n_556),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_527),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_554),
.B(n_555),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_536),
.B(n_511),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_515),
.Y(n_556)
);

FAx1_ASAP7_75t_SL g557 ( 
.A(n_547),
.B(n_520),
.CI(n_524),
.CON(n_557),
.SN(n_557)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_560),
.A2(n_544),
.B(n_548),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_534),
.C(n_543),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_523),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_562),
.A2(n_557),
.B(n_552),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_567),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_551),
.A2(n_538),
.B(n_545),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_565),
.A2(n_566),
.B(n_552),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_561),
.A2(n_537),
.B(n_517),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_559),
.A2(n_501),
.B(n_517),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_SL g572 ( 
.A1(n_568),
.A2(n_557),
.B(n_553),
.Y(n_572)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_571),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_572),
.A2(n_569),
.B(n_558),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_573),
.B(n_570),
.C(n_558),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_575),
.A2(n_569),
.B(n_563),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_576),
.A2(n_521),
.B(n_494),
.Y(n_578)
);

AOI321xp33_ASAP7_75t_SL g579 ( 
.A1(n_577),
.A2(n_578),
.A3(n_574),
.B1(n_532),
.B2(n_539),
.C(n_504),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_579),
.A2(n_511),
.B1(n_282),
.B2(n_7),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_282),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_582)
);


endmodule