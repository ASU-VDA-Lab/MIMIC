module fake_aes_12465_n_726 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_726);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_726;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_59), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_1), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_18), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_49), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_3), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g117 ( .A(n_62), .B(n_91), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_104), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_3), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_69), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_16), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_33), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_8), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_43), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_13), .Y(n_126) );
XOR2xp5_ASAP7_75t_L g127 ( .A(n_78), .B(n_16), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_18), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_105), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_6), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_4), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_28), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_44), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_5), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_92), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_46), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_17), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_102), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_50), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_58), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_37), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_64), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
INVxp67_ASAP7_75t_SL g151 ( .A(n_103), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_124), .B(n_1), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_124), .B(n_2), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_122), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_114), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_109), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_120), .B(n_2), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_135), .B(n_5), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_114), .B(n_22), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_168), .Y(n_173) );
NAND3xp33_ASAP7_75t_L g174 ( .A(n_165), .B(n_130), .C(n_110), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_168), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_164), .B(n_129), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_168), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_168), .Y(n_178) );
AND2x6_ASAP7_75t_L g179 ( .A(n_153), .B(n_136), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_160), .B(n_136), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_160), .B(n_119), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_168), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_153), .A2(n_121), .B1(n_112), .B2(n_126), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_165), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_172), .B(n_138), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
NOR2x1p5_ASAP7_75t_L g194 ( .A(n_167), .B(n_123), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_153), .B(n_138), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_186), .B(n_153), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_192), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_192), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_192), .B(n_153), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_193), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_185), .B(n_169), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_193), .B(n_162), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_193), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_179), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
OAI221xp5_ASAP7_75t_L g209 ( .A1(n_182), .A2(n_167), .B1(n_155), .B2(n_172), .C(n_171), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_194), .B(n_169), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_179), .B(n_162), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_195), .A2(n_169), .B(n_162), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_179), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_187), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_179), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_179), .B(n_171), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_179), .B(n_171), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_174), .B(n_171), .Y(n_218) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_197), .B(n_115), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_176), .A2(n_155), .B1(n_111), .B2(n_131), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_197), .B(n_118), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_197), .B(n_132), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_170), .B(n_166), .C(n_163), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_197), .A2(n_142), .B1(n_113), .B2(n_116), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_188), .A2(n_170), .B(n_166), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_189), .B(n_140), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_197), .B(n_188), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_197), .B(n_163), .Y(n_228) );
NAND2xp33_ASAP7_75t_L g229 ( .A(n_196), .B(n_141), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_196), .B(n_146), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_175), .B(n_147), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_175), .B(n_148), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_190), .A2(n_163), .B(n_166), .C(n_170), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_207), .B(n_175), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_210), .B(n_128), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_227), .A2(n_183), .B(n_177), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_205), .Y(n_237) );
OAI21xp33_ASAP7_75t_SL g238 ( .A1(n_204), .A2(n_127), .B(n_113), .Y(n_238) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_225), .A2(n_180), .B(n_177), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_199), .A2(n_127), .B1(n_116), .B2(n_121), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_207), .B(n_175), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_199), .B(n_112), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_227), .A2(n_202), .B(n_216), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_210), .A2(n_125), .B1(n_137), .B2(n_126), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_218), .B(n_133), .Y(n_245) );
AOI33xp33_ASAP7_75t_L g246 ( .A1(n_220), .A2(n_133), .A3(n_137), .B1(n_143), .B2(n_142), .B3(n_139), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_205), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_207), .B(n_175), .Y(n_248) );
BUFx8_ASAP7_75t_L g249 ( .A(n_207), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_202), .A2(n_178), .B(n_173), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_224), .B(n_143), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_212), .A2(n_139), .B(n_145), .C(n_150), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_178), .B(n_173), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_208), .A2(n_180), .B(n_183), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_209), .A2(n_145), .B1(n_150), .B2(n_152), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_226), .B(n_151), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_152), .B(n_191), .C(n_190), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_208), .A2(n_184), .B(n_198), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_211), .A2(n_184), .B(n_198), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_207), .A2(n_117), .B1(n_159), .B2(n_191), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
AOI22x1_ASAP7_75t_L g262 ( .A1(n_203), .A2(n_159), .B1(n_161), .B2(n_156), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_213), .A2(n_159), .B1(n_161), .B2(n_156), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_200), .A2(n_161), .B(n_156), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_250), .A2(n_219), .B(n_200), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_237), .B(n_225), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_235), .B(n_214), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_239), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_214), .B(n_228), .Y(n_269) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_252), .A2(n_228), .A3(n_201), .B(n_206), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_264), .A2(n_233), .B(n_201), .Y(n_271) );
AOI31xp67_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_203), .A3(n_206), .B(n_230), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_247), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_261), .B(n_213), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_262), .A2(n_231), .B(n_221), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_235), .B(n_229), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_252), .A2(n_215), .B(n_222), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_251), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_240), .A2(n_215), .B1(n_232), .B2(n_161), .Y(n_279) );
NAND2xp33_ASAP7_75t_SL g280 ( .A(n_246), .B(n_6), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_249), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_236), .A2(n_161), .B(n_156), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_253), .A2(n_161), .B(n_156), .Y(n_283) );
O2A1O1Ixp5_ASAP7_75t_SL g284 ( .A1(n_260), .A2(n_161), .B(n_156), .C(n_154), .Y(n_284) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_258), .A2(n_156), .B(n_154), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_238), .B(n_7), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_254), .A2(n_154), .B(n_54), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_249), .Y(n_288) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_268), .A2(n_255), .B(n_259), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_284), .A2(n_257), .B(n_263), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_273), .B(n_244), .Y(n_291) );
CKINVDCx11_ASAP7_75t_R g292 ( .A(n_288), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_282), .A2(n_256), .B(n_245), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_284), .A2(n_248), .B(n_241), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g295 ( .A(n_286), .B(n_280), .C(n_279), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_281), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_275), .A2(n_248), .B(n_241), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_283), .A2(n_255), .B(n_234), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_273), .B(n_234), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_266), .B(n_7), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_275), .A2(n_154), .B(n_55), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_285), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_278), .A2(n_154), .B(n_9), .C(n_10), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_278), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_300), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_307), .B(n_270), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_309), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_291), .B(n_276), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_307), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_309), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_304), .A2(n_287), .B(n_265), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_302), .B(n_270), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_292), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_302), .B(n_270), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_291), .B(n_281), .Y(n_320) );
AOI21x1_ASAP7_75t_L g321 ( .A1(n_304), .A2(n_271), .B(n_269), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_308), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_308), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_301), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
OR2x6_ASAP7_75t_SL g329 ( .A(n_295), .B(n_267), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_300), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_297), .A2(n_277), .B1(n_269), .B2(n_274), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_303), .B(n_270), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_322), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_319), .B(n_305), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_331), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_333), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_314), .B(n_270), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_319), .B(n_305), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_331), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_331), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_334), .B(n_305), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_334), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_334), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_335), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_311), .A2(n_293), .A3(n_299), .B(n_306), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_313), .A2(n_295), .B1(n_274), .B2(n_289), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_335), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_324), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_327), .B(n_289), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_310), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_327), .B(n_289), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_310), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_328), .B(n_289), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_326), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_326), .B(n_289), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_330), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_328), .B(n_298), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_325), .B(n_298), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_315), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_317), .B(n_298), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_310), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_311), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_317), .B(n_293), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_336), .B(n_294), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_336), .B(n_294), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_338), .B(n_310), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_338), .B(n_310), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_340), .B(n_312), .Y(n_384) );
OR2x6_ASAP7_75t_L g385 ( .A(n_371), .B(n_321), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_351), .B(n_320), .C(n_299), .D(n_329), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_340), .B(n_332), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_371), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_349), .B(n_316), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_370), .B(n_321), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_373), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_337), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_371), .B(n_318), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_373), .B(n_8), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_349), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_366), .B(n_329), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_343), .B(n_316), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_343), .B(n_316), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_339), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_339), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_294), .Y(n_403) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_355), .B(n_274), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_370), .B(n_304), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_358), .B(n_154), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_361), .B(n_154), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_339), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_361), .B(n_9), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_344), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_357), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_344), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_366), .B(n_360), .Y(n_415) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_355), .B(n_274), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_363), .B(n_10), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_360), .B(n_377), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_345), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_367), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_370), .B(n_290), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_377), .B(n_11), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_367), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_363), .B(n_11), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_375), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_375), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_370), .B(n_290), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_345), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_374), .B(n_12), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_372), .B(n_290), .Y(n_430) );
AND2x4_ASAP7_75t_SL g431 ( .A(n_346), .B(n_272), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_345), .Y(n_432) );
INVx5_ASAP7_75t_SL g433 ( .A(n_342), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_347), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_347), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_346), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_347), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_374), .B(n_14), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_378), .B(n_14), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_372), .B(n_65), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_342), .Y(n_441) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_346), .B(n_272), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_341), .B(n_15), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_348), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_379), .B(n_15), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_348), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_379), .B(n_17), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_381), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_388), .B(n_348), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_409), .B(n_341), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_401), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_388), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_399), .B(n_380), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_409), .B(n_380), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_378), .Y(n_456) );
AND2x4_ASAP7_75t_SL g457 ( .A(n_388), .B(n_352), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_436), .B(n_352), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_384), .B(n_352), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_385), .B(n_359), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_381), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_445), .B(n_365), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_417), .B(n_365), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_445), .B(n_365), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_392), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_392), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_393), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_384), .B(n_354), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_393), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_397), .B(n_354), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_396), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_401), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_406), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_447), .B(n_354), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_417), .B(n_351), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_402), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_408), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_447), .B(n_356), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_400), .B(n_376), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_400), .B(n_376), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_429), .B(n_356), .Y(n_482) );
OR2x6_ASAP7_75t_L g483 ( .A(n_385), .B(n_356), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_406), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_396), .Y(n_485) );
NAND2xp67_ASAP7_75t_L g486 ( .A(n_398), .B(n_364), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_413), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_424), .B(n_364), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_382), .B(n_359), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_382), .B(n_364), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_413), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_408), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_410), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_410), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_429), .B(n_368), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_383), .B(n_359), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_407), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_407), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_424), .B(n_368), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_412), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_438), .B(n_368), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_385), .B(n_362), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_415), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_383), .B(n_362), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_418), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_420), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_411), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_403), .B(n_369), .Y(n_508) );
OAI21xp33_ASAP7_75t_SL g509 ( .A1(n_416), .A2(n_369), .B(n_362), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_403), .B(n_369), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_394), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_420), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_385), .B(n_362), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_390), .B(n_421), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_411), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_414), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_438), .B(n_350), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_425), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_439), .B(n_350), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_430), .B(n_350), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_387), .B(n_350), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_430), .B(n_350), .Y(n_522) );
NOR2x1p5_ASAP7_75t_L g523 ( .A(n_386), .B(n_342), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_430), .B(n_350), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_421), .B(n_350), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_422), .B(n_19), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_414), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_425), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_421), .B(n_342), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_426), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_404), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_448), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_456), .B(n_426), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_457), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_526), .A2(n_395), .B(n_439), .C(n_443), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_511), .B(n_387), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_500), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_456), .B(n_423), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_503), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_389), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_523), .B(n_440), .Y(n_542) );
OAI21xp33_ASAP7_75t_SL g543 ( .A1(n_453), .A2(n_416), .B(n_389), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_473), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_484), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_484), .B(n_428), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_505), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_449), .Y(n_548) );
NOR2x1p5_ASAP7_75t_SL g549 ( .A(n_521), .B(n_419), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_461), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_465), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_466), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_457), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_526), .B(n_440), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_467), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_454), .B(n_427), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_454), .B(n_427), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_469), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_470), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_471), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_485), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_462), .B(n_427), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_531), .B(n_440), .Y(n_563) );
AND2x4_ASAP7_75t_SL g564 ( .A(n_531), .B(n_419), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_455), .B(n_404), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_450), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_464), .B(n_390), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_487), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_491), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_489), .B(n_390), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_475), .B(n_428), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_496), .B(n_405), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_519), .B(n_432), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_504), .B(n_405), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_506), .B(n_432), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_512), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_480), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_479), .B(n_437), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_480), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_518), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_528), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_481), .B(n_405), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_481), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_530), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_497), .B(n_433), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_486), .Y(n_586) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_483), .B(n_437), .Y(n_587) );
NAND2x2_ASAP7_75t_L g588 ( .A(n_453), .B(n_19), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_514), .B(n_431), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_459), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_468), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_497), .B(n_433), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_498), .B(n_433), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_458), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_482), .B(n_444), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_495), .B(n_444), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_508), .B(n_434), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_508), .B(n_434), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_498), .B(n_433), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_452), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_509), .A2(n_446), .B(n_435), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_490), .B(n_442), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_510), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_488), .B(n_446), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_514), .B(n_442), .Y(n_605) );
OAI22xp33_ASAP7_75t_SL g606 ( .A1(n_483), .A2(n_435), .B1(n_441), .B2(n_431), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_510), .B(n_441), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_490), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_514), .B(n_441), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_533), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_588), .A2(n_483), .B1(n_517), .B2(n_451), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_543), .A2(n_501), .B(n_499), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_536), .A2(n_522), .B1(n_524), .B2(n_520), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_535), .A2(n_476), .B(n_460), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_533), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_544), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g617 ( .A1(n_534), .A2(n_507), .B(n_472), .C(n_527), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_540), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_535), .A2(n_525), .B(n_520), .C(n_524), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_534), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_554), .A2(n_522), .B1(n_525), .B2(n_529), .Y(n_621) );
OAI21xp33_ASAP7_75t_SL g622 ( .A1(n_566), .A2(n_529), .B(n_527), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_556), .B(n_502), .Y(n_623) );
AOI21xp33_ASAP7_75t_SL g624 ( .A1(n_544), .A2(n_460), .B(n_513), .Y(n_624) );
OA21x2_ASAP7_75t_L g625 ( .A1(n_601), .A2(n_502), .B(n_513), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_547), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_537), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_573), .B(n_452), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_539), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_549), .A2(n_460), .B(n_502), .C(n_513), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_557), .B(n_472), .Y(n_631) );
AOI322xp5_ASAP7_75t_L g632 ( .A1(n_579), .A2(n_516), .A3(n_515), .B1(n_507), .B2(n_494), .C1(n_493), .C2(n_492), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_579), .B(n_474), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_539), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_573), .B(n_474), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_586), .A2(n_516), .B(n_515), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_553), .A2(n_494), .B1(n_493), .B2(n_492), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_567), .B(n_478), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_553), .A2(n_478), .B(n_477), .C(n_342), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_583), .B(n_562), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_566), .A2(n_477), .B1(n_342), .B2(n_277), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_532), .Y(n_642) );
AOI222xp33_ASAP7_75t_L g643 ( .A1(n_601), .A2(n_20), .B1(n_21), .B2(n_342), .C1(n_271), .C2(n_25), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_542), .B(n_20), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_591), .B(n_594), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_564), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_546), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_591), .B(n_21), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_587), .A2(n_23), .B(n_24), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_606), .A2(n_26), .B(n_27), .C(n_29), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_590), .B(n_538), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_565), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_548), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_603), .B(n_34), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_550), .A2(n_35), .B1(n_36), .B2(n_38), .C(n_39), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_551), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_563), .A2(n_41), .B(n_42), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_545), .B(n_107), .Y(n_658) );
AO21x1_ASAP7_75t_L g659 ( .A1(n_589), .A2(n_45), .B(n_47), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_608), .B(n_48), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_617), .A2(n_605), .B(n_589), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_619), .A2(n_605), .B(n_609), .C(n_570), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_646), .A2(n_541), .B1(n_609), .B2(n_577), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_614), .B(n_580), .C(n_555), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_614), .A2(n_602), .B1(n_582), .B2(n_607), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_622), .B(n_559), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_644), .A2(n_607), .B(n_585), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_610), .B(n_552), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_620), .A2(n_592), .B(n_593), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_611), .A2(n_572), .B1(n_599), .B2(n_574), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_646), .A2(n_598), .B1(n_597), .B2(n_578), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_624), .A2(n_659), .B(n_620), .C(n_630), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_645), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_643), .B(n_576), .C(n_560), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_628), .B(n_597), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_643), .B(n_581), .C(n_561), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_648), .A2(n_598), .B(n_558), .Y(n_677) );
XOR2xp5_ASAP7_75t_L g678 ( .A(n_621), .B(n_571), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_635), .B(n_604), .Y(n_679) );
XOR2xp5_ASAP7_75t_L g680 ( .A(n_613), .B(n_596), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_642), .B(n_584), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_616), .A2(n_569), .B(n_568), .C(n_575), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_612), .A2(n_595), .B(n_575), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_647), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_625), .A2(n_600), .B(n_52), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_615), .B(n_51), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_653), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_629), .A2(n_53), .B1(n_56), .B2(n_57), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g689 ( .A1(n_640), .A2(n_60), .A3(n_63), .B1(n_66), .B2(n_67), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_634), .B(n_68), .Y(n_690) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_618), .A2(n_70), .A3(n_71), .B1(n_73), .B2(n_75), .C1(n_77), .C2(n_79), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_626), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_625), .A2(n_80), .B(n_82), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_641), .B(n_83), .C(n_84), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g695 ( .A1(n_650), .A2(n_86), .B(n_87), .C(n_88), .Y(n_695) );
AOI211xp5_ASAP7_75t_SL g696 ( .A1(n_657), .A2(n_90), .B(n_94), .C(n_95), .Y(n_696) );
AND3x1_ASAP7_75t_L g697 ( .A(n_639), .B(n_96), .C(n_97), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_627), .B(n_98), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_656), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_632), .B(n_99), .C(n_100), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_637), .A2(n_101), .B1(n_106), .B2(n_636), .C(n_651), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_649), .B(n_654), .C(n_652), .D(n_655), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_664), .A2(n_683), .B1(n_672), .B2(n_671), .Y(n_703) );
AOI211xp5_ASAP7_75t_SL g704 ( .A1(n_693), .A2(n_695), .B(n_701), .C(n_685), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_700), .B(n_702), .C(n_694), .Y(n_705) );
NAND4xp75_ASAP7_75t_L g706 ( .A(n_667), .B(n_666), .C(n_697), .D(n_661), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_692), .B(n_680), .Y(n_707) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_689), .B(n_662), .C(n_649), .Y(n_708) );
NOR3x1_ASAP7_75t_L g709 ( .A(n_676), .B(n_674), .C(n_669), .Y(n_709) );
NAND4xp25_ASAP7_75t_SL g710 ( .A(n_703), .B(n_670), .C(n_665), .D(n_682), .Y(n_710) );
NOR2x1_ASAP7_75t_L g711 ( .A(n_706), .B(n_663), .Y(n_711) );
NAND4xp75_ASAP7_75t_L g712 ( .A(n_709), .B(n_677), .C(n_690), .D(n_686), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_708), .B(n_658), .C(n_660), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_710), .B(n_705), .C(n_707), .Y(n_714) );
NAND4xp75_ASAP7_75t_L g715 ( .A(n_711), .B(n_677), .C(n_688), .D(n_704), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_712), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_716), .B(n_713), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_715), .Y(n_718) );
AOI22x1_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_714), .B1(n_678), .B2(n_673), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_717), .B(n_681), .Y(n_720) );
OAI22x1_ASAP7_75t_L g721 ( .A1(n_719), .A2(n_717), .B1(n_684), .B2(n_687), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_720), .A2(n_699), .B1(n_675), .B2(n_668), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_722), .B(n_679), .Y(n_723) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_721), .B(n_698), .Y(n_724) );
AO21x2_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_623), .B(n_691), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_633), .B1(n_638), .B2(n_631), .C(n_696), .Y(n_726) );
endmodule