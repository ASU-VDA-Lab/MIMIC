module fake_jpeg_3661_n_349 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_46),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_15),
.B(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_56),
.Y(n_107)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_17),
.A2(n_11),
.B(n_13),
.Y(n_50)
);

OR2x4_ASAP7_75t_L g146 ( 
.A(n_50),
.B(n_13),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_25),
.B(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g152 ( 
.A(n_63),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_9),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_64),
.B(n_82),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_21),
.B(n_9),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_9),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_84),
.Y(n_126)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_87),
.Y(n_108)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_88),
.B(n_97),
.Y(n_149)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_95),
.Y(n_123)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_94),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_93),
.Y(n_153)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_98),
.Y(n_130)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_44),
.Y(n_135)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_34),
.B1(n_40),
.B2(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_150),
.B1(n_49),
.B2(n_70),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_64),
.A2(n_82),
.B1(n_77),
.B2(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_118),
.B1(n_139),
.B2(n_144),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_47),
.A2(n_34),
.B1(n_40),
.B2(n_38),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_29),
.B1(n_28),
.B2(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_44),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_148),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_60),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_42),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_51),
.A2(n_39),
.B1(n_28),
.B2(n_29),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_96),
.B1(n_52),
.B2(n_80),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_162),
.B1(n_180),
.B2(n_190),
.Y(n_204)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_71),
.B1(n_67),
.B2(n_31),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_187),
.B(n_188),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_79),
.B1(n_72),
.B2(n_68),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_57),
.B1(n_95),
.B2(n_73),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_154),
.B1(n_110),
.B2(n_140),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_78),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_178),
.Y(n_203)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_78),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_63),
.B1(n_85),
.B2(n_87),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_184),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_112),
.B(n_0),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_1),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_14),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_141),
.B1(n_109),
.B2(n_111),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_136),
.B1(n_154),
.B2(n_104),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_149),
.B(n_119),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_213),
.B(n_217),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_134),
.B(n_145),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_136),
.B1(n_120),
.B2(n_103),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_216),
.B1(n_163),
.B2(n_174),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_109),
.B(n_140),
.C(n_111),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_182),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_235),
.B(n_221),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_230),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_157),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_227),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_161),
.B(n_171),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_202),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_229),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_157),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_157),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_166),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_160),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_204),
.B1(n_215),
.B2(n_197),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_165),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_189),
.B(n_133),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_133),
.B(n_113),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_247),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_231),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_242),
.B1(n_253),
.B2(n_254),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_206),
.B1(n_210),
.B2(n_204),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_225),
.B(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_216),
.B1(n_127),
.B2(n_120),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_236),
.B1(n_234),
.B2(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_202),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_222),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_211),
.B1(n_177),
.B2(n_127),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_222),
.B1(n_218),
.B2(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_261),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_266),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_268),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_256),
.B1(n_250),
.B2(n_244),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_285),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_231),
.C(n_246),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_280),
.C(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_246),
.C(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_223),
.B1(n_240),
.B2(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_245),
.C(n_242),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_245),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_224),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_240),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_243),
.B(n_250),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_208),
.B(n_198),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_299),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_270),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_300),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_264),
.B1(n_263),
.B2(n_265),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_272),
.B1(n_273),
.B2(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_241),
.B1(n_236),
.B2(n_234),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_279),
.B1(n_275),
.B2(n_228),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_212),
.B(n_191),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_303),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_277),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_294),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_288),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.C(n_312),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_274),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_276),
.C(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_297),
.C(n_295),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.C(n_310),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_285),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_301),
.C(n_209),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_205),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_205),
.C(n_200),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_322),
.B(n_184),
.Y(n_330)
);

AO221x1_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.C(n_198),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_323),
.B(n_327),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_326),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_313),
.B1(n_311),
.B2(n_176),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_328),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_196),
.C(n_200),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_196),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_168),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_319),
.C(n_110),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_333),
.B(n_334),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_113),
.C(n_151),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_151),
.B(n_159),
.Y(n_337)
);

AOI221xp5_ASAP7_75t_L g342 ( 
.A1(n_337),
.A2(n_129),
.B1(n_115),
.B2(n_1),
.C(n_14),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_179),
.C(n_129),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_339),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_179),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_179),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_129),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_342),
.Y(n_346)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_340),
.B(n_338),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_345),
.B(n_343),
.C(n_115),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_346),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_115),
.Y(n_349)
);


endmodule