module real_jpeg_21626_n_5 (n_4, n_0, n_1, n_26, n_2, n_27, n_28, n_29, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_26;
input n_2;
input n_27;
input n_28;
input n_29;
input n_3;

output n_5;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_23;
wire n_11;
wire n_14;
wire n_7;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

BUFx16f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_1),
.B(n_15),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_13),
.C(n_23),
.Y(n_12)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g6 ( 
.A1(n_4),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

XOR2xp5_ASAP7_75t_L g5 ( 
.A(n_6),
.B(n_12),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_19),
.C(n_20),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_26),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_27),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_28),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_29),
.Y(n_24)
);


endmodule