module real_jpeg_24666_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_47),
.B1(n_54),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_47),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_2),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_2),
.A2(n_40),
.B1(n_42),
.B2(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_146),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_146),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_32),
.B1(n_40),
.B2(n_42),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_32),
.B1(n_54),
.B2(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_4),
.A2(n_57),
.B(n_147),
.C(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_4),
.B(n_55),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_36),
.B(n_42),
.C(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_4),
.B(n_24),
.C(n_27),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_4),
.B(n_95),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_4),
.B(n_11),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_4),
.B(n_26),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_7),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_52),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_11),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_90),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_88),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_74),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_15),
.B(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_65),
.B2(n_73),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_33),
.C(n_48),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_18),
.A2(n_33),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_18),
.A2(n_78),
.B1(n_84),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_18),
.A2(n_78),
.B1(n_190),
.B2(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_29),
.B(n_30),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_19),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_20),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_20),
.B(n_31),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_22),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_25),
.A2(n_32),
.B(n_37),
.Y(n_232)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_26),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_26),
.B(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_27),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_27),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_29),
.B(n_30),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_29),
.A2(n_99),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_32),
.A2(n_42),
.B(n_56),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_43),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_34),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_38),
.B(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_35),
.B(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_39),
.B(n_85),
.Y(n_139)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_43),
.A2(n_86),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_43),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_44),
.B(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_55),
.B(n_58),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_61)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_51),
.Y(n_145)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_62),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_55),
.B(n_81),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_55),
.B(n_144),
.Y(n_176)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_60),
.B(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_66),
.B(n_165),
.C(n_175),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_66),
.A2(n_71),
.B1(n_175),
.B2(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_68),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_70),
.B(n_143),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_83),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_75),
.A2(n_79),
.B1(n_104),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.C(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_78),
.B(n_188),
.C(n_190),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_80),
.B(n_176),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_87),
.B(n_199),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI211xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_148),
.B(n_154),
.C(n_318),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_122),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_122),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_92),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_101),
.CI(n_106),
.CON(n_92),
.SN(n_92)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_94),
.B(n_96),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_101),
.C(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_95),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_97),
.B(n_234),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_99),
.B(n_246),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_114),
.B(n_118),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_118),
.B1(n_119),
.B2(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_115),
.B1(n_126),
.B2(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_107),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_107),
.A2(n_126),
.B1(n_231),
.B2(n_290),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_113),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_108),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_108),
.B(n_113),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_108),
.B(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_112),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_117),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_117),
.B(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_127),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.C(n_140),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_130),
.B(n_136),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_131),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_134),
.A2(n_168),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_134),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_139),
.B(n_192),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_155),
.C(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_150),
.B(n_151),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_180),
.B(n_317),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_177),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_158),
.B(n_177),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_159),
.B(n_162),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_164),
.B(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_165),
.A2(n_166),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_173),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_170),
.B(n_259),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_174),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_312),
.B(n_316),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_224),
.B(n_299),
.C(n_311),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_212),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_183),
.B(n_212),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_196),
.B2(n_211),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_194),
.B2(n_195),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_186),
.B(n_195),
.C(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_189),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_193),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_198),
.B(n_203),
.C(n_204),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.C(n_219),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_214),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_222),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_298),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_240),
.B(n_297),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_227),
.B(n_237),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_230),
.B(n_233),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_231),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_292),
.B(n_296),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_283),
.B(n_291),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_263),
.B(n_282),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_244),
.B(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_270),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_245),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_262),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_256),
.C(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_271),
.B(n_281),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_269),
.Y(n_281)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_277),
.B(n_280),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_279),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_285),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_310),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_308),
.B2(n_309),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_309),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_314),
.Y(n_316)
);


endmodule