module fake_jpeg_19680_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_24),
.B1(n_30),
.B2(n_16),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_53),
.B1(n_40),
.B2(n_34),
.Y(n_81)
);

NAND2x1p5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_15),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_38),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_24),
.B1(n_16),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_37),
.B1(n_36),
.B2(n_16),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_24),
.B1(n_36),
.B2(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_62),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_76),
.B(n_78),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_39),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_41),
.B(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_24),
.A3(n_40),
.B1(n_34),
.B2(n_54),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

AOI22x1_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_110),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_39),
.C(n_33),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_57),
.C(n_60),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_99),
.B1(n_113),
.B2(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_112),
.B1(n_84),
.B2(n_68),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_106),
.B(n_19),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_59),
.B(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_22),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_28),
.B1(n_26),
.B2(n_21),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_120),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_93),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_64),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_125),
.C(n_108),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_129),
.B1(n_107),
.B2(n_103),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_65),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_119),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_131),
.B1(n_136),
.B2(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_17),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_124),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_67),
.C(n_63),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_67),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_77),
.B1(n_21),
.B2(n_28),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_27),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_66),
.B1(n_26),
.B2(n_22),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_139),
.Y(n_160)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_19),
.B1(n_23),
.B2(n_9),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_25),
.B1(n_9),
.B2(n_14),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_27),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_137),
.B(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_138),
.A2(n_100),
.B1(n_97),
.B2(n_91),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_94),
.B(n_20),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_27),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_94),
.B1(n_108),
.B2(n_98),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_158),
.C(n_163),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_151),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_112),
.B(n_92),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_160),
.B(n_143),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

AO21x2_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_92),
.B(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_172),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_6),
.C(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_95),
.B(n_92),
.C(n_19),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_19),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_87),
.B1(n_109),
.B2(n_95),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_118),
.B1(n_124),
.B2(n_151),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_173),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_19),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_0),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_87),
.B1(n_109),
.B2(n_23),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_23),
.B1(n_25),
.B2(n_20),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_20),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_189),
.B1(n_167),
.B2(n_149),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_178),
.B(n_180),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_139),
.B(n_119),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_202),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_123),
.B(n_131),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_186),
.B(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_115),
.B1(n_136),
.B2(n_123),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_194),
.B1(n_150),
.B2(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_200),
.C(n_8),
.Y(n_227)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_7),
.C(n_13),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_0),
.B(n_1),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_1),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_145),
.A2(n_153),
.B(n_160),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_150),
.B(n_165),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_153),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_211),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_217),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_179),
.B1(n_203),
.B2(n_181),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_172),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_227),
.Y(n_239)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_176),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_148),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_174),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_202),
.B(n_181),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_190),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_243),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_241),
.B(n_244),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_186),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_223),
.C(n_220),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_193),
.B(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_196),
.C(n_188),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_214),
.C(n_215),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_214),
.B1(n_208),
.B2(n_216),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_246),
.A2(n_220),
.B1(n_212),
.B2(n_222),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_207),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_251),
.B1(n_262),
.B2(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_255),
.C(n_258),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_191),
.B1(n_177),
.B2(n_212),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_257),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_235),
.B1(n_229),
.B2(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_234),
.C(n_230),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_187),
.B1(n_218),
.B2(n_175),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_195),
.C(n_192),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_201),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_200),
.C(n_185),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_240),
.C(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_183),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_274),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_183),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_269),
.A2(n_272),
.B1(n_249),
.B2(n_256),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_244),
.B1(n_182),
.B2(n_194),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_227),
.C(n_241),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_258),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_275),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_14),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_284),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_271),
.B(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_8),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_8),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_272),
.Y(n_293)
);

NOR2x1p5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_282),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_267),
.B(n_273),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_297),
.B(n_298),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_276),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_288),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_265),
.B(n_266),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_11),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_304),
.B(n_296),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_294),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_303),
.B(n_299),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_308),
.A2(n_306),
.B(n_307),
.C(n_11),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_11),
.C(n_12),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_12),
.B(n_4),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_3),
.C(n_4),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_5),
.C(n_306),
.Y(n_313)
);


endmodule