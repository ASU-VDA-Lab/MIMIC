module fake_jpeg_2426_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_14),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_42),
.Y(n_65)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_65),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_43),
.B1(n_52),
.B2(n_50),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_57),
.B1(n_59),
.B2(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_51),
.B1(n_53),
.B2(n_41),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_56),
.B1(n_41),
.B2(n_47),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_56),
.B(n_54),
.C(n_51),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_63),
.B(n_62),
.C(n_44),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_85),
.B1(n_75),
.B2(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_23),
.B1(n_37),
.B2(n_33),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_85),
.A2(n_64),
.B1(n_62),
.B2(n_44),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_90),
.B1(n_100),
.B2(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_50),
.B1(n_40),
.B2(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_99),
.Y(n_102)
);

BUFx2_ASAP7_75t_SL g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_49),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_16),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_92),
.C(n_87),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_112),
.B(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_4),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_5),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_6),
.Y(n_116)
);

NOR4xp25_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_7),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_124),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_105),
.C(n_108),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_8),
.B(n_9),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_22),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_24),
.C(n_28),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_106),
.B1(n_11),
.B2(n_12),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_134),
.Y(n_138)
);

OAI322xp33_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_115),
.A3(n_106),
.B1(n_25),
.B2(n_27),
.C1(n_17),
.C2(n_19),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_126),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_143),
.B(n_128),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_127),
.C(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_121),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_139),
.B1(n_133),
.B2(n_125),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_141),
.B(n_124),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_148),
.A2(n_134),
.B1(n_122),
.B2(n_38),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_30),
.Y(n_150)
);


endmodule