module fake_jpeg_11513_n_11 (n_0, n_3, n_2, n_1, n_11);

input n_0;
input n_3;
input n_2;
input n_1;

output n_11;

wire n_10;
wire n_4;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx3_ASAP7_75t_L g4 ( 
.A(n_1),
.Y(n_4)
);

AOI22xp33_ASAP7_75t_L g5 ( 
.A1(n_0),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

AOI22xp5_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_7)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_7),
.B(n_8),
.Y(n_9)
);

AOI322xp5_ASAP7_75t_L g8 ( 
.A1(n_5),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_6),
.C1(n_4),
.C2(n_1),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_5),
.Y(n_10)
);

OAI211xp5_ASAP7_75t_L g11 ( 
.A1(n_10),
.A2(n_7),
.B(n_4),
.C(n_0),
.Y(n_11)
);


endmodule