module real_aes_8251_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_729, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_729;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g462 ( .A1(n_0), .A2(n_200), .B(n_463), .C(n_466), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_1), .B(n_457), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_1), .A2(n_713), .B1(n_714), .B2(n_722), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_1), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g122 ( .A(n_2), .Y(n_122) );
INVx1_ASAP7_75t_L g235 ( .A(n_3), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_4), .B(n_152), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_5), .A2(n_452), .B(n_540), .Y(n_539) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_6), .A2(n_175), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_7), .A2(n_38), .B1(n_145), .B2(n_169), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_8), .B(n_175), .Y(n_247) );
AND2x6_ASAP7_75t_L g160 ( .A(n_9), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_10), .A2(n_160), .B(n_443), .C(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_11), .B(n_39), .Y(n_114) );
INVx1_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_13), .B(n_150), .Y(n_183) );
INVx1_ASAP7_75t_L g227 ( .A(n_14), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_15), .A2(n_76), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_15), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_16), .B(n_152), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_17), .B(n_176), .Y(n_214) );
AO32x2_ASAP7_75t_L g197 ( .A1(n_18), .A2(n_174), .A3(n_175), .B1(n_198), .B2(n_202), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_19), .B(n_145), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_20), .B(n_176), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_21), .A2(n_56), .B1(n_145), .B2(n_169), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g172 ( .A1(n_22), .A2(n_82), .B1(n_145), .B2(n_150), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_23), .B(n_145), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_24), .A2(n_174), .B(n_443), .C(n_490), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_25), .A2(n_174), .B(n_443), .C(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_26), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_27), .B(n_137), .Y(n_256) );
OAI22xp5_ASAP7_75t_SL g699 ( .A1(n_28), .A2(n_94), .B1(n_700), .B2(n_701), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_28), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_29), .A2(n_698), .B1(n_699), .B2(n_702), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_29), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_30), .A2(n_452), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_31), .B(n_137), .Y(n_162) );
INVx2_ASAP7_75t_L g147 ( .A(n_32), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_33), .A2(n_449), .B(n_475), .C(n_476), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_34), .B(n_145), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_35), .B(n_137), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_36), .A2(n_43), .B1(n_433), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_36), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_37), .B(n_185), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_40), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_41), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_42), .B(n_152), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_43), .A2(n_128), .B1(n_433), .B2(n_434), .Y(n_127) );
INVx1_ASAP7_75t_L g433 ( .A(n_43), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_44), .B(n_452), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_45), .B(n_117), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_46), .A2(n_449), .B(n_475), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_47), .B(n_145), .Y(n_242) );
INVx1_ASAP7_75t_L g464 ( .A(n_48), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_49), .A2(n_92), .B1(n_169), .B2(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g527 ( .A(n_50), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_51), .B(n_145), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_52), .B(n_145), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_53), .A2(n_696), .B1(n_697), .B2(n_703), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_53), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_54), .B(n_452), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_55), .B(n_233), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g218 ( .A1(n_57), .A2(n_61), .B1(n_145), .B2(n_150), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_58), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_59), .B(n_145), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_60), .B(n_145), .Y(n_255) );
INVx1_ASAP7_75t_L g161 ( .A(n_62), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_63), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_64), .B(n_457), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_65), .A2(n_230), .B(n_233), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_66), .B(n_145), .Y(n_236) );
INVx1_ASAP7_75t_L g140 ( .A(n_67), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_68), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_69), .B(n_152), .Y(n_480) );
AO32x2_ASAP7_75t_L g166 ( .A1(n_70), .A2(n_167), .A3(n_173), .B1(n_174), .B2(n_175), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_71), .B(n_153), .Y(n_517) );
INVx1_ASAP7_75t_L g254 ( .A(n_72), .Y(n_254) );
INVx1_ASAP7_75t_L g148 ( .A(n_73), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_74), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_75), .B(n_479), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_76), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_77), .A2(n_443), .B(n_445), .C(n_449), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_78), .B(n_150), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_79), .Y(n_541) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_81), .B(n_478), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_83), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_84), .B(n_169), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_85), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_86), .B(n_150), .Y(n_157) );
INVx2_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_88), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_89), .B(n_171), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_90), .B(n_150), .Y(n_243) );
INVx2_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
OR2x2_ASAP7_75t_L g119 ( .A(n_91), .B(n_120), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_93), .A2(n_104), .B1(n_150), .B2(n_151), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_94), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_95), .B(n_452), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_96), .A2(n_106), .B1(n_115), .B2(n_726), .Y(n_105) );
INVx1_ASAP7_75t_L g477 ( .A(n_97), .Y(n_477) );
INVxp67_ASAP7_75t_L g544 ( .A(n_98), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_99), .B(n_150), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g446 ( .A(n_101), .Y(n_446) );
INVx1_ASAP7_75t_L g513 ( .A(n_102), .Y(n_513) );
AND2x2_ASAP7_75t_L g529 ( .A(n_103), .B(n_137), .Y(n_529) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_107), .Y(n_727) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
AO22x2_ASAP7_75t_SL g126 ( .A1(n_109), .A2(n_127), .B1(n_435), .B2(n_694), .Y(n_126) );
INVx1_ASAP7_75t_L g694 ( .A(n_109), .Y(n_694) );
NOR2x2_ASAP7_75t_L g708 ( .A(n_109), .B(n_120), .Y(n_708) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g121 ( .A(n_114), .B(n_122), .Y(n_121) );
NAND2x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_123), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g725 ( .A(n_119), .Y(n_725) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_121), .A2(n_125), .B1(n_126), .B2(n_695), .C(n_704), .Y(n_124) );
OAI321xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_705), .A3(n_709), .B1(n_712), .B2(n_723), .C(n_724), .Y(n_123) );
INVx1_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g434 ( .A(n_128), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_128), .A2(n_434), .B1(n_719), .B2(n_720), .Y(n_718) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_354), .Y(n_128) );
NAND3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_303), .C(n_345), .Y(n_129) );
AOI211xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_208), .B(n_257), .C(n_279), .Y(n_130) );
OAI211xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_163), .B(n_191), .C(n_203), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_133), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g366 ( .A(n_133), .B(n_283), .Y(n_366) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g268 ( .A(n_134), .B(n_194), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_134), .B(n_179), .Y(n_385) );
INVx1_ASAP7_75t_L g403 ( .A(n_134), .Y(n_403) );
AND2x2_ASAP7_75t_L g412 ( .A(n_134), .B(n_300), .Y(n_412) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g295 ( .A(n_135), .B(n_179), .Y(n_295) );
AND2x2_ASAP7_75t_L g353 ( .A(n_135), .B(n_300), .Y(n_353) );
INVx1_ASAP7_75t_L g397 ( .A(n_135), .Y(n_397) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g274 ( .A(n_136), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g282 ( .A(n_136), .Y(n_282) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_136), .Y(n_322) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_142), .B(n_162), .Y(n_136) );
INVx2_ASAP7_75t_L g173 ( .A(n_137), .Y(n_173) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_137), .A2(n_180), .B(n_190), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_137), .A2(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g496 ( .A(n_137), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_137), .A2(n_524), .B(n_525), .Y(n_523) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_L g176 ( .A(n_138), .B(n_139), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_155), .B(n_160), .Y(n_142) );
O2A1O1Ixp5_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_148), .B(n_149), .C(n_152), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_145), .Y(n_448) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
AND2x6_ASAP7_75t_L g443 ( .A(n_146), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g151 ( .A(n_147), .Y(n_151) );
INVx1_ASAP7_75t_L g234 ( .A(n_147), .Y(n_234) );
INVx2_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_152), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_152), .A2(n_251), .B(n_252), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_152), .B(n_544), .Y(n_543) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_153), .A2(n_168), .B1(n_171), .B2(n_172), .Y(n_167) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_154), .Y(n_159) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
INVx1_ASAP7_75t_L g444 ( .A(n_154), .Y(n_444) );
AND2x2_ASAP7_75t_L g453 ( .A(n_154), .B(n_234), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_158), .Y(n_155) );
INVx1_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g479 ( .A(n_159), .Y(n_479) );
BUFx3_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_160), .A2(n_181), .B(n_186), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_160), .A2(n_226), .B(n_231), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_160), .A2(n_241), .B(n_244), .Y(n_240) );
INVx4_ASAP7_75t_SL g450 ( .A(n_160), .Y(n_450) );
AND2x4_ASAP7_75t_L g452 ( .A(n_160), .B(n_453), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_160), .B(n_453), .Y(n_514) );
INVxp67_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_177), .Y(n_164) );
AND2x2_ASAP7_75t_L g261 ( .A(n_165), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g294 ( .A(n_165), .Y(n_294) );
OR2x2_ASAP7_75t_L g420 ( .A(n_165), .B(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_165), .B(n_179), .Y(n_424) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g194 ( .A(n_166), .Y(n_194) );
INVx1_ASAP7_75t_L g206 ( .A(n_166), .Y(n_206) );
AND2x2_ASAP7_75t_L g283 ( .A(n_166), .B(n_196), .Y(n_283) );
AND2x2_ASAP7_75t_L g323 ( .A(n_166), .B(n_197), .Y(n_323) );
INVx2_ASAP7_75t_L g466 ( .A(n_170), .Y(n_466) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_170), .Y(n_481) );
INVx2_ASAP7_75t_L g189 ( .A(n_171), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_171), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_171), .A2(n_200), .B1(n_217), .B2(n_218), .Y(n_216) );
INVx4_ASAP7_75t_L g465 ( .A(n_171), .Y(n_465) );
INVx1_ASAP7_75t_L g493 ( .A(n_173), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_174), .B(n_216), .C(n_219), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_174), .A2(n_250), .B(n_253), .Y(n_249) );
INVx4_ASAP7_75t_L g219 ( .A(n_175), .Y(n_219) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_175), .A2(n_240), .B(n_247), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_175), .A2(n_503), .B(n_504), .Y(n_502) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_175), .Y(n_538) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g202 ( .A(n_176), .Y(n_202) );
INVxp67_ASAP7_75t_L g365 ( .A(n_177), .Y(n_365) );
AND2x4_ASAP7_75t_L g390 ( .A(n_177), .B(n_283), .Y(n_390) );
BUFx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_178), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g195 ( .A(n_179), .B(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g269 ( .A(n_179), .B(n_197), .Y(n_269) );
INVx1_ASAP7_75t_L g275 ( .A(n_179), .Y(n_275) );
INVx2_ASAP7_75t_L g301 ( .A(n_179), .Y(n_301) );
AND2x2_ASAP7_75t_L g317 ( .A(n_179), .B(n_318), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
O2A1O1Ixp5_ASAP7_75t_L g253 ( .A1(n_189), .A2(n_232), .B(n_254), .C(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_192), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
BUFx2_ASAP7_75t_L g272 ( .A(n_194), .Y(n_272) );
AND2x2_ASAP7_75t_L g380 ( .A(n_194), .B(n_196), .Y(n_380) );
AND2x2_ASAP7_75t_L g297 ( .A(n_195), .B(n_282), .Y(n_297) );
AND2x2_ASAP7_75t_L g396 ( .A(n_195), .B(n_397), .Y(n_396) );
NOR2xp67_ASAP7_75t_L g318 ( .A(n_196), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g421 ( .A(n_196), .B(n_282), .Y(n_421) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g207 ( .A(n_197), .Y(n_207) );
AND2x2_ASAP7_75t_L g300 ( .A(n_197), .B(n_301), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_200), .A2(n_232), .B(n_235), .C(n_236), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_200), .A2(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g224 ( .A(n_202), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_202), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
AND2x2_ASAP7_75t_L g346 ( .A(n_205), .B(n_281), .Y(n_346) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_206), .B(n_282), .Y(n_331) );
INVx2_ASAP7_75t_L g330 ( .A(n_207), .Y(n_330) );
OAI222xp33_ASAP7_75t_L g334 ( .A1(n_207), .A2(n_274), .B1(n_335), .B2(n_337), .C1(n_338), .C2(n_341), .Y(n_334) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g259 ( .A(n_212), .Y(n_259) );
OR2x2_ASAP7_75t_L g370 ( .A(n_212), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
NOR2x1_ASAP7_75t_L g343 ( .A(n_213), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g349 ( .A(n_213), .B(n_263), .Y(n_349) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g310 ( .A(n_214), .Y(n_310) );
AO21x1_ASAP7_75t_L g309 ( .A1(n_216), .A2(n_219), .B(n_310), .Y(n_309) );
AO21x2_ASAP7_75t_L g440 ( .A1(n_219), .A2(n_441), .B(n_454), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_219), .B(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g457 ( .A(n_219), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_219), .B(n_483), .Y(n_482) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_219), .A2(n_512), .B(n_519), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_220), .A2(n_313), .B1(n_352), .B2(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_238), .Y(n_220) );
INVx3_ASAP7_75t_L g285 ( .A(n_221), .Y(n_285) );
OR2x2_ASAP7_75t_L g418 ( .A(n_221), .B(n_294), .Y(n_418) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g291 ( .A(n_222), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g307 ( .A(n_222), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g315 ( .A(n_222), .B(n_263), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_222), .B(n_239), .Y(n_371) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g262 ( .A(n_223), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g266 ( .A(n_223), .B(n_239), .Y(n_266) );
AND2x2_ASAP7_75t_L g342 ( .A(n_223), .B(n_289), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_223), .B(n_248), .Y(n_382) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_237), .Y(n_223) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_224), .A2(n_249), .B(n_256), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .C(n_230), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_228), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_228), .A2(n_517), .B(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_230), .A2(n_446), .B(n_447), .C(n_448), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_232), .A2(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_238), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_238), .B(n_259), .Y(n_298) );
AND2x2_ASAP7_75t_L g302 ( .A(n_238), .B(n_292), .Y(n_302) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
INVx3_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
AND2x2_ASAP7_75t_L g288 ( .A(n_239), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g423 ( .A(n_239), .B(n_406), .Y(n_423) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_248), .Y(n_277) );
INVx2_ASAP7_75t_L g289 ( .A(n_248), .Y(n_289) );
AND2x2_ASAP7_75t_L g333 ( .A(n_248), .B(n_309), .Y(n_333) );
INVx1_ASAP7_75t_L g376 ( .A(n_248), .Y(n_376) );
OR2x2_ASAP7_75t_L g407 ( .A(n_248), .B(n_309), .Y(n_407) );
AND2x2_ASAP7_75t_L g427 ( .A(n_248), .B(n_263), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_264), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g265 ( .A(n_259), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_259), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g384 ( .A(n_261), .Y(n_384) );
INVx2_ASAP7_75t_SL g278 ( .A(n_262), .Y(n_278) );
AND2x2_ASAP7_75t_L g398 ( .A(n_262), .B(n_292), .Y(n_398) );
INVx2_ASAP7_75t_L g344 ( .A(n_263), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_263), .B(n_376), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B1(n_270), .B2(n_276), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_266), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g432 ( .A(n_266), .Y(n_432) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g357 ( .A(n_268), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_268), .B(n_300), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_269), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g373 ( .A(n_269), .B(n_322), .Y(n_373) );
INVx2_ASAP7_75t_L g429 ( .A(n_269), .Y(n_429) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x2_ASAP7_75t_L g299 ( .A(n_272), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_272), .B(n_317), .Y(n_350) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_274), .B(n_294), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g411 ( .A(n_277), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_SL g361 ( .A1(n_278), .A2(n_362), .B(n_364), .C(n_367), .Y(n_361) );
OR2x2_ASAP7_75t_L g388 ( .A(n_278), .B(n_292), .Y(n_388) );
OAI221xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_284), .B1(n_286), .B2(n_293), .C(n_296), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_281), .B(n_330), .Y(n_337) );
AND2x2_ASAP7_75t_L g379 ( .A(n_281), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g415 ( .A(n_281), .Y(n_415) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_282), .Y(n_306) );
INVx1_ASAP7_75t_L g319 ( .A(n_282), .Y(n_319) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_285), .B(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g393 ( .A(n_285), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_285), .B(n_333), .Y(n_409) );
INVx2_ASAP7_75t_L g395 ( .A(n_286), .Y(n_395) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g336 ( .A(n_288), .B(n_307), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_288), .A2(n_304), .B(n_346), .C(n_347), .Y(n_345) );
AND2x2_ASAP7_75t_L g314 ( .A(n_289), .B(n_309), .Y(n_314) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_293), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
OR2x2_ASAP7_75t_L g362 ( .A(n_294), .B(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_299), .B2(n_302), .Y(n_296) );
INVx1_ASAP7_75t_L g416 ( .A(n_298), .Y(n_416) );
INVx1_ASAP7_75t_L g363 ( .A(n_300), .Y(n_363) );
INVx1_ASAP7_75t_L g414 ( .A(n_302), .Y(n_414) );
AOI211xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_307), .B(n_311), .C(n_334), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g326 ( .A(n_306), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g377 ( .A(n_307), .Y(n_377) );
AND2x2_ASAP7_75t_L g426 ( .A(n_307), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B(n_324), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_314), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g332 ( .A(n_315), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g408 ( .A(n_315), .Y(n_408) );
OAI32xp33_ASAP7_75t_L g419 ( .A1(n_315), .A2(n_367), .A3(n_374), .B1(n_415), .B2(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_320), .Y(n_316) );
INVx1_ASAP7_75t_SL g387 ( .A(n_317), .Y(n_387) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g327 ( .A(n_323), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B(n_332), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_326), .A2(n_374), .B1(n_400), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_330), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_353), .A2(n_395), .B1(n_396), .B2(n_398), .C(n_399), .Y(n_394) );
NAND5xp2_ASAP7_75t_L g354 ( .A(n_355), .B(n_378), .C(n_394), .D(n_404), .E(n_422), .Y(n_354) );
AOI211xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_361), .C(n_368), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g425 ( .A(n_362), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_372), .B2(n_374), .Y(n_368) );
INVx1_ASAP7_75t_SL g401 ( .A(n_371), .Y(n_401) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI322xp33_ASAP7_75t_L g383 ( .A1(n_374), .A2(n_384), .A3(n_385), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_389), .Y(n_383) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g386 ( .A(n_376), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_376), .B(n_401), .Y(n_400) );
AOI211xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_381), .B(n_383), .C(n_391), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_387), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_413) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g430 ( .A(n_397), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_412), .B1(n_413), .B2(n_417), .C(n_419), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_408), .B(n_409), .C(n_410), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g431 ( .A(n_407), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_425), .B2(n_426), .C(n_428), .Y(n_422) );
AOI21xp33_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_430), .B(n_431), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_436), .B(n_637), .Y(n_435) );
AND4x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_577), .C(n_592), .D(n_617), .Y(n_436) );
NOR2xp33_ASAP7_75t_SL g437 ( .A(n_438), .B(n_550), .Y(n_437) );
OAI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_468), .B(n_530), .Y(n_438) );
AND2x2_ASAP7_75t_L g580 ( .A(n_439), .B(n_485), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_439), .B(n_484), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_439), .B(n_469), .Y(n_643) );
INVx1_ASAP7_75t_L g647 ( .A(n_439), .Y(n_647) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_456), .Y(n_439) );
INVx2_ASAP7_75t_L g564 ( .A(n_440), .Y(n_564) );
BUFx2_ASAP7_75t_L g591 ( .A(n_440), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_451), .Y(n_441) );
INVx5_ASAP7_75t_L g461 ( .A(n_443), .Y(n_461) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_SL g459 ( .A1(n_450), .A2(n_460), .B(n_461), .C(n_462), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_450), .A2(n_461), .B(n_541), .C(n_542), .Y(n_540) );
BUFx2_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
AND2x2_ASAP7_75t_L g531 ( .A(n_456), .B(n_485), .Y(n_531) );
INVx2_ASAP7_75t_L g547 ( .A(n_456), .Y(n_547) );
AND2x2_ASAP7_75t_L g556 ( .A(n_456), .B(n_484), .Y(n_556) );
AND2x2_ASAP7_75t_L g635 ( .A(n_456), .B(n_564), .Y(n_635) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_467), .Y(n_456) );
INVx2_ASAP7_75t_L g475 ( .A(n_461), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_497), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_469), .B(n_562), .Y(n_600) );
INVx1_ASAP7_75t_L g688 ( .A(n_469), .Y(n_688) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_484), .Y(n_469) );
AND2x2_ASAP7_75t_L g546 ( .A(n_470), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g560 ( .A(n_470), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_470), .Y(n_589) );
OR2x2_ASAP7_75t_L g621 ( .A(n_470), .B(n_563), .Y(n_621) );
AND2x2_ASAP7_75t_L g629 ( .A(n_470), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g662 ( .A(n_470), .B(n_631), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_470), .B(n_531), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_470), .B(n_591), .Y(n_687) );
AND2x2_ASAP7_75t_L g693 ( .A(n_470), .B(n_580), .Y(n_693) );
INVx5_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g553 ( .A(n_471), .Y(n_553) );
AND2x2_ASAP7_75t_L g583 ( .A(n_471), .B(n_563), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_471), .B(n_576), .Y(n_616) );
AND2x2_ASAP7_75t_L g636 ( .A(n_471), .B(n_485), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_471), .B(n_536), .Y(n_670) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_480), .C(n_481), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_478), .A2(n_481), .B(n_527), .C(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g576 ( .A(n_484), .B(n_547), .Y(n_576) );
AND2x2_ASAP7_75t_L g587 ( .A(n_484), .B(n_583), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_484), .B(n_563), .Y(n_626) );
INVx2_ASAP7_75t_L g641 ( .A(n_484), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_484), .B(n_575), .Y(n_664) );
AND2x2_ASAP7_75t_L g683 ( .A(n_484), .B(n_635), .Y(n_683) );
INVx5_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_485), .Y(n_582) );
AND2x2_ASAP7_75t_L g590 ( .A(n_485), .B(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g631 ( .A(n_485), .B(n_547), .Y(n_631) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_489), .B(n_493), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
AND2x2_ASAP7_75t_L g554 ( .A(n_499), .B(n_537), .Y(n_554) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_500), .B(n_511), .Y(n_534) );
OR2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_537), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_500), .B(n_537), .Y(n_572) );
AND2x2_ASAP7_75t_L g599 ( .A(n_500), .B(n_536), .Y(n_599) );
AND2x2_ASAP7_75t_L g651 ( .A(n_500), .B(n_510), .Y(n_651) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_501), .B(n_521), .Y(n_559) );
AND2x2_ASAP7_75t_L g595 ( .A(n_501), .B(n_511), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_508), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g585 ( .A(n_509), .B(n_567), .Y(n_585) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
OAI322xp33_ASAP7_75t_L g550 ( .A1(n_510), .A2(n_551), .A3(n_555), .B1(n_557), .B2(n_560), .C1(n_565), .C2(n_573), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_510), .B(n_536), .Y(n_558) );
OR2x2_ASAP7_75t_L g568 ( .A(n_510), .B(n_522), .Y(n_568) );
AND2x2_ASAP7_75t_L g570 ( .A(n_510), .B(n_522), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_510), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_510), .B(n_537), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_510), .B(n_666), .Y(n_665) );
INVx5_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_511), .B(n_554), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_521), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g548 ( .A(n_521), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_521), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g610 ( .A(n_521), .B(n_537), .Y(n_610) );
AOI211xp5_ASAP7_75t_SL g638 ( .A1(n_521), .A2(n_639), .B(n_642), .C(n_654), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_521), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g676 ( .A(n_521), .B(n_651), .Y(n_676) );
INVx5_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g604 ( .A(n_522), .B(n_537), .Y(n_604) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
AND2x2_ASAP7_75t_L g653 ( .A(n_522), .B(n_651), .Y(n_653) );
AND2x2_ASAP7_75t_SL g684 ( .A(n_522), .B(n_554), .Y(n_684) );
AND2x2_ASAP7_75t_L g691 ( .A(n_522), .B(n_650), .Y(n_691) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_529), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B1(n_546), .B2(n_548), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_531), .B(n_553), .Y(n_601) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g549 ( .A(n_534), .Y(n_549) );
OR2x2_ASAP7_75t_L g609 ( .A(n_534), .B(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_534), .A2(n_658), .B1(n_660), .B2(n_661), .C(n_663), .Y(n_657) );
INVx2_ASAP7_75t_L g596 ( .A(n_535), .Y(n_596) );
AND2x2_ASAP7_75t_L g569 ( .A(n_536), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g659 ( .A(n_536), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_536), .B(n_651), .Y(n_672) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_L g614 ( .A(n_537), .Y(n_614) );
AND2x2_ASAP7_75t_L g650 ( .A(n_537), .B(n_651), .Y(n_650) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B(n_545), .Y(n_537) );
AND2x2_ASAP7_75t_L g652 ( .A(n_546), .B(n_591), .Y(n_652) );
AND2x2_ASAP7_75t_L g562 ( .A(n_547), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_547), .B(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_SL g633 ( .A(n_549), .B(n_596), .Y(n_633) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g639 ( .A(n_552), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OR2x2_ASAP7_75t_L g625 ( .A(n_553), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g690 ( .A(n_553), .B(n_635), .Y(n_690) );
INVx2_ASAP7_75t_L g623 ( .A(n_554), .Y(n_623) );
NAND4xp25_ASAP7_75t_SL g686 ( .A(n_555), .B(n_687), .C(n_688), .D(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_556), .B(n_620), .Y(n_655) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_SL g692 ( .A(n_559), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_SL g654 ( .A1(n_560), .A2(n_623), .B(n_627), .C(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g649 ( .A(n_562), .B(n_641), .Y(n_649) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_563), .Y(n_575) );
INVx1_ASAP7_75t_L g630 ( .A(n_563), .Y(n_630) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_564), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B(n_569), .C(n_571), .Y(n_565) );
AND2x2_ASAP7_75t_L g586 ( .A(n_566), .B(n_570), .Y(n_586) );
OAI322xp33_ASAP7_75t_SL g624 ( .A1(n_566), .A2(n_625), .A3(n_627), .B1(n_628), .B2(n_632), .C1(n_633), .C2(n_634), .Y(n_624) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g646 ( .A(n_568), .B(n_572), .Y(n_646) );
INVx1_ASAP7_75t_L g627 ( .A(n_570), .Y(n_627) );
INVx1_ASAP7_75t_SL g645 ( .A(n_572), .Y(n_645) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AOI222xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_584), .B1(n_586), .B2(n_587), .C1(n_588), .C2(n_729), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
OAI322xp33_ASAP7_75t_L g667 ( .A1(n_579), .A2(n_641), .A3(n_646), .B1(n_668), .B2(n_669), .C1(n_671), .C2(n_672), .Y(n_667) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_580), .A2(n_594), .B1(n_618), .B2(n_622), .C(n_624), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OAI222xp33_ASAP7_75t_L g597 ( .A1(n_585), .A2(n_598), .B1(n_600), .B2(n_601), .C1(n_602), .C2(n_605), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_587), .A2(n_594), .B1(n_664), .B2(n_665), .Y(n_663) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AOI211xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_597), .C(n_608), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_594), .A2(n_631), .B(n_674), .C(n_677), .Y(n_673) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g603 ( .A(n_595), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g666 ( .A(n_599), .Y(n_666) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_606), .B(n_631), .Y(n_660) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B(n_615), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g677 ( .A1(n_609), .A2(n_678), .B1(n_679), .B2(n_680), .C(n_681), .Y(n_677) );
INVxp33_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_613), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_620), .B(n_631), .Y(n_671) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g682 ( .A(n_635), .B(n_641), .Y(n_682) );
AND4x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_656), .C(n_673), .D(n_685), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_644), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g678 ( .A(n_649), .Y(n_678) );
INVx1_ASAP7_75t_SL g668 ( .A(n_653), .Y(n_668) );
NOR2xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_667), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_669), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_676), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g704 ( .A(n_695), .Y(n_704) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx3_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g723 ( .A(n_711), .Y(n_723) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
XNOR2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
endmodule