module fake_jpeg_25162_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_65),
.B(n_69),
.Y(n_122)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_73),
.B(n_82),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_90),
.C(n_42),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_40),
.B1(n_44),
.B2(n_24),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_81),
.B1(n_83),
.B2(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_25),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_24),
.B1(n_36),
.B2(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_23),
.B1(n_28),
.B2(n_25),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_96),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_32),
.B1(n_45),
.B2(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_16),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_35),
.Y(n_116)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_109),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_32),
.B1(n_17),
.B2(n_34),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_107),
.B1(n_27),
.B2(n_31),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_20),
.B1(n_17),
.B2(n_34),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_94),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_87),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_72),
.A2(n_90),
.B1(n_82),
.B2(n_71),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_76),
.B1(n_66),
.B2(n_92),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_77),
.B(n_68),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_93),
.B(n_85),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_35),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_78),
.B1(n_81),
.B2(n_74),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_129),
.B(n_133),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_103),
.B1(n_98),
.B2(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_91),
.B1(n_89),
.B2(n_86),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_127),
.B1(n_99),
.B2(n_101),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_144),
.B(n_135),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_152),
.C(n_140),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_84),
.B1(n_17),
.B2(n_18),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_33),
.B1(n_21),
.B2(n_27),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_16),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_34),
.B1(n_20),
.B2(n_104),
.Y(n_187)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_85),
.B(n_35),
.C(n_30),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_34),
.B(n_18),
.C(n_20),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_121),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_21),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_33),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_30),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_112),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_174),
.B1(n_180),
.B2(n_114),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_103),
.B(n_120),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_161),
.A2(n_162),
.B(n_182),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_164),
.B1(n_169),
.B2(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_120),
.B1(n_99),
.B2(n_101),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_119),
.B1(n_102),
.B2(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_168),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_33),
.B1(n_21),
.B2(n_112),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_141),
.B1(n_149),
.B2(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_148),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_112),
.C(n_105),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_152),
.C(n_155),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_31),
.B1(n_18),
.B2(n_20),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_152),
.B(n_142),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_31),
.B(n_26),
.Y(n_182)
);

AOI31xp33_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_16),
.A3(n_26),
.B(n_18),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_181),
.C(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_139),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_191),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_199),
.C(n_164),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_194),
.B1(n_207),
.B2(n_221),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_156),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_183),
.B(n_137),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_152),
.C(n_154),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_202),
.B(n_208),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_148),
.B(n_132),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_209),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_218),
.B(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_112),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_9),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_175),
.B(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_185),
.B1(n_176),
.B2(n_172),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_185),
.B(n_161),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_241),
.C(n_212),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_182),
.C(n_168),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_199),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_215),
.B(n_218),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_189),
.C(n_181),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_168),
.B1(n_189),
.B2(n_181),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_168),
.B(n_158),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_207),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_195),
.A2(n_114),
.B1(n_42),
.B2(n_26),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_250),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_191),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_259),
.Y(n_275)
);

AOI22x1_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_201),
.B1(n_200),
.B2(n_213),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_252),
.A2(n_248),
.B1(n_229),
.B2(n_245),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_220),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_231),
.B(n_205),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_203),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_264),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_208),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_203),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_269),
.B1(n_227),
.B2(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_267),
.B(n_246),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_197),
.Y(n_268)
);

INVx13_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_270),
.B(n_271),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_233),
.B1(n_247),
.B2(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_248),
.C(n_224),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_283),
.C(n_287),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_247),
.B1(n_227),
.B2(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_224),
.C(n_197),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_286),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_244),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_258),
.CI(n_263),
.CON(n_289),
.SN(n_289)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_256),
.C(n_254),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_298),
.C(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_256),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_254),
.C(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_204),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_274),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_7),
.C(n_13),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_0),
.B(n_2),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_283),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_303),
.B(n_278),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_306),
.B(n_307),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_287),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_281),
.B(n_274),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_285),
.B1(n_278),
.B2(n_3),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_313),
.B1(n_296),
.B2(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_309),
.B(n_312),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_285),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_315),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_291),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_289),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_288),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_291),
.C(n_294),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_295),
.C(n_296),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_295),
.B1(n_289),
.B2(n_301),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_310),
.B(n_299),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_306),
.B(n_308),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_324),
.B(n_321),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_311),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.C(n_318),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_313),
.C(n_10),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_326),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_325),
.C(n_10),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_10),
.Y(n_336)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_8),
.A3(n_13),
.B1(n_5),
.B2(n_6),
.C1(n_14),
.C2(n_11),
.Y(n_337)
);

AOI31xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_5),
.A3(n_11),
.B(n_12),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_12),
.Y(n_341)
);


endmodule