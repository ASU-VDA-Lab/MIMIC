module fake_jpeg_14662_n_96 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_26),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_0),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_36),
.Y(n_40)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_45),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_25),
.B1(n_12),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_47),
.B1(n_41),
.B2(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_13),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_38),
.Y(n_63)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_48),
.C(n_51),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_30),
.B(n_27),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_49),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_58),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_51),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_50),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.C(n_59),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_56),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.C(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_52),
.B1(n_60),
.B2(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_83),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_68),
.C(n_64),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_23),
.B(n_27),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_87),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_28),
.C(n_30),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_92),
.C(n_30),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_93),
.Y(n_96)
);


endmodule