module fake_jpeg_8496_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_5),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_4),
.B(n_3),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_14),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_0),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_17),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_18),
.B1(n_12),
.B2(n_11),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

OA21x2_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_8),
.B(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_23),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_8),
.B1(n_12),
.B2(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_19),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_11),
.C(n_14),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_32),
.C(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

AOI21x1_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_30),
.B(n_15),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_12),
.C(n_37),
.Y(n_38)
);

BUFx24_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);


endmodule