module fake_jpeg_31940_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_42),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_61),
.Y(n_74)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_0),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_0),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_35),
.B1(n_15),
.B2(n_36),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_80),
.B1(n_102),
.B2(n_5),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_19),
.C(n_37),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_68),
.B(n_78),
.C(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_15),
.B1(n_35),
.B2(n_39),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_79),
.A2(n_94),
.B1(n_100),
.B2(n_101),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_21),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_82),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_4),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_103),
.B1(n_106),
.B2(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_39),
.B1(n_32),
.B2(n_29),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_2),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_9),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_113),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_60),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_41),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_96),
.B1(n_94),
.B2(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_141),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_118),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_6),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_130),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_66),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_134),
.Y(n_155)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_120),
.B1(n_117),
.B2(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_6),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_91),
.B(n_112),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_6),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_122),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_69),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_135),
.A2(n_107),
.B1(n_76),
.B2(n_78),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_67),
.B(n_69),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_64),
.B(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_99),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_123),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_65),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_89),
.A2(n_86),
.B(n_87),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_99),
.B1(n_95),
.B2(n_75),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_71),
.B1(n_81),
.B2(n_111),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_71),
.B1(n_81),
.B2(n_97),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_177),
.B1(n_180),
.B2(n_138),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_165),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_76),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_152),
.B(n_172),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_104),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_161),
.B1(n_170),
.B2(n_121),
.Y(n_187)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_163),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_99),
.B1(n_75),
.B2(n_111),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_129),
.B2(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_70),
.B1(n_85),
.B2(n_92),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_164),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_70),
.B1(n_99),
.B2(n_97),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_134),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_142),
.B1(n_125),
.B2(n_119),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_124),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_114),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_122),
.B(n_131),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_138),
.Y(n_191)
);

INVx11_ASAP7_75t_SL g175 ( 
.A(n_141),
.Y(n_175)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_125),
.B1(n_119),
.B2(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_140),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_181),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_121),
.A2(n_126),
.B1(n_144),
.B2(n_128),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_134),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_144),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_184),
.B(n_200),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_161),
.B1(n_153),
.B2(n_169),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_190),
.A2(n_157),
.B1(n_174),
.B2(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_191),
.B(n_210),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_127),
.B(n_138),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_193),
.A2(n_212),
.B(n_174),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_197),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_164),
.B1(n_153),
.B2(n_146),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_190),
.B1(n_193),
.B2(n_176),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_149),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_178),
.B(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_202),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_173),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_151),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_148),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_180),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_218),
.B1(n_206),
.B2(n_195),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_155),
.B1(n_153),
.B2(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_156),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_183),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_159),
.B(n_155),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_230),
.B(n_231),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_238),
.B1(n_184),
.B2(n_200),
.Y(n_250)
);

XOR2x2_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_153),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_198),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_184),
.A2(n_174),
.B(n_196),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_206),
.B(n_200),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_236),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_185),
.C(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_194),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_215),
.B1(n_187),
.B2(n_191),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_212),
.B(n_183),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_232),
.B(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_219),
.B1(n_228),
.B2(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_185),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_216),
.B1(n_206),
.B2(n_233),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_199),
.C(n_201),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_250),
.C(n_225),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_219),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_199),
.Y(n_257)
);

NOR4xp25_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_246),
.C(n_256),
.D(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_195),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_198),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_234),
.B1(n_229),
.B2(n_220),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_244),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_225),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_265),
.C(n_270),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_267),
.B1(n_252),
.B2(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_182),
.B1(n_230),
.B2(n_238),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_241),
.B1(n_255),
.B2(n_259),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_231),
.C(n_239),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_252),
.C(n_248),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_284),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_285),
.C(n_274),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_281),
.B1(n_286),
.B2(n_186),
.Y(n_297)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_242),
.C(n_247),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_249),
.B1(n_258),
.B2(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_241),
.C(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_262),
.B(n_264),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_296),
.B(n_214),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_265),
.B(n_240),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_261),
.C(n_240),
.Y(n_298)
);

OAI221xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_282),
.B1(n_285),
.B2(n_278),
.C(n_204),
.Y(n_301)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_237),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_306),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_186),
.B(n_188),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_188),
.B(n_203),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_295),
.B1(n_293),
.B2(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_311),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_292),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_290),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_315),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_303),
.B1(n_296),
.B2(n_298),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_314),
.A2(n_312),
.B(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_315),
.C(n_302),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_311),
.Y(n_320)
);


endmodule