module real_jpeg_3974_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_1),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_1),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_126),
.B1(n_161),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_1),
.A2(n_56),
.B1(n_126),
.B2(n_277),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_1),
.A2(n_126),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_59),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_59),
.B1(n_113),
.B2(n_130),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_3),
.A2(n_59),
.B1(n_358),
.B2(n_360),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_4),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_4),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_4),
.A2(n_89),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_5),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_162),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_5),
.A2(n_88),
.B1(n_162),
.B2(n_286),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_5),
.A2(n_162),
.B1(n_344),
.B2(n_346),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_6),
.A2(n_74),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_7),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_7),
.A2(n_57),
.B1(n_209),
.B2(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_7),
.B(n_51),
.C(n_217),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_7),
.B(n_114),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_7),
.B(n_292),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_7),
.B(n_61),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_7),
.B(n_353),
.Y(n_352)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_9),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_9),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_9),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_9),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_10),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_10),
.A2(n_68),
.B1(n_138),
.B2(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_10),
.A2(n_138),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_10),
.A2(n_138),
.B1(n_228),
.B2(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_11),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_13),
.A2(n_72),
.B1(n_76),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_13),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_14),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_14),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_14),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_14),
.Y(n_163)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_16),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_16),
.A2(n_67),
.B1(n_71),
.B2(n_216),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_16),
.A2(n_67),
.B1(n_124),
.B2(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_261),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_260),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_234),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_21),
.B(n_234),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_168),
.C(n_185),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_22),
.A2(n_23),
.B1(n_168),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_96),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_24),
.B(n_97),
.C(n_167),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_69),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_25),
.B(n_69),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_52),
.B1(n_60),
.B2(n_62),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_26),
.A2(n_270),
.B(n_275),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_26),
.A2(n_60),
.B1(n_300),
.B2(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_26),
.A2(n_275),
.B(n_343),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_61),
.B1(n_63),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_27),
.A2(n_61),
.B1(n_170),
.B2(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_27),
.B(n_276),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_32),
.Y(n_172)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_32),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_41),
.A2(n_300),
.B(n_302),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_44),
.Y(n_296)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_48),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_52),
.A2(n_60),
.B(n_302),
.Y(n_409)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_58),
.Y(n_176)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_58),
.Y(n_274)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_58),
.Y(n_278)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_61),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_68),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_79),
.B1(n_86),
.B2(n_93),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_73),
.Y(n_295)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_77),
.Y(n_359)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_78),
.Y(n_311)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_79),
.B(n_293),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_79),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_79),
.A2(n_215),
.B1(n_357),
.B2(n_389),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_85),
.Y(n_289)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_87),
.A2(n_178),
.B1(n_179),
.B2(n_183),
.Y(n_177)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_95),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_134),
.B1(n_166),
.B2(n_167),
.Y(n_96)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_114),
.B1(n_122),
.B2(n_128),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_98),
.A2(n_224),
.B(n_232),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_98),
.A2(n_232),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_98),
.B(n_122),
.Y(n_385)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_99),
.A2(n_129),
.B1(n_233),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_99),
.A2(n_225),
.B1(n_233),
.B2(n_381),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_110),
.B2(n_112),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g363 ( 
.A(n_108),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_108),
.Y(n_384)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_109),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_109),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_110),
.B(n_242),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_114),
.Y(n_233)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_116),
.Y(n_301)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_121),
.Y(n_369)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_123),
.B(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_141),
.B1(n_159),
.B2(n_164),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_164),
.B(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g405 ( 
.A1(n_139),
.A2(n_208),
.B(n_209),
.Y(n_405)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_141),
.A2(n_159),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_142),
.A2(n_405),
.B(n_406),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_153),
.B1(n_155),
.B2(n_157),
.Y(n_152)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_164),
.B(n_209),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_165),
.B(n_189),
.Y(n_259)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_168),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_169),
.B(n_177),
.Y(n_252)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_214),
.B1(n_219),
.B2(n_222),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_178),
.A2(n_183),
.B(n_247),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_178),
.A2(n_285),
.B(n_290),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_178),
.A2(n_209),
.B(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_182),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_185),
.B(n_424),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.C(n_223),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_186),
.A2(n_187),
.B1(n_223),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_192),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_212),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_193),
.A2(n_212),
.B1(n_213),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_193),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_198),
.A3(n_201),
.B1(n_204),
.B2(n_208),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_197),
.Y(n_350)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_209),
.A2(n_350),
.B(n_351),
.Y(n_349)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_223),
.Y(n_419)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_233),
.A2(n_381),
.B(n_385),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g434 ( 
.A(n_234),
.Y(n_434)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.CI(n_251),
.CON(n_234),
.SN(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_246),
.B2(n_250),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_SL g281 ( 
.A(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_259),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_412),
.B(n_431),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_393),
.B(n_411),
.Y(n_263)
);

AO21x1_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_372),
.B(n_392),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_337),
.B(n_371),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_305),
.B(n_336),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_283),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_268),
.B(n_283),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_279),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_269),
.A2(n_279),
.B1(n_280),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_274),
.Y(n_366)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_297),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_298),
.C(n_304),
.Y(n_338)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_288),
.Y(n_360)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_303),
.B2(n_304),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_327),
.B(n_335),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_314),
.B(n_326),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_325),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_322),
.B(n_324),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_324),
.A2(n_356),
.B(n_361),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_333),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_333),
.Y(n_335)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_339),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_354),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_347),
.B2(n_348),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_347),
.C(n_354),
.Y(n_373)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI32xp33_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_363),
.A3(n_364),
.B1(n_367),
.B2(n_370),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_362),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_362),
.Y(n_378)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_373),
.B(n_374),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_379),
.B2(n_391),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_378),
.C(n_391),
.Y(n_394)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_379),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_386),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_387),
.C(n_388),
.Y(n_399)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx12f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_394),
.B(n_395),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_402),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_396)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_400),
.C(n_402),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_407),
.B2(n_410),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_408),
.C(n_409),
.Y(n_422)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_407),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_426),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_415),
.A2(n_432),
.B(n_433),
.Y(n_431)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_423),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_423),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_422),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_420),
.A2(n_421),
.B1(n_422),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_428),
.Y(n_432)
);


endmodule