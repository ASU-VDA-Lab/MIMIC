module real_jpeg_32804_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_1),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_1),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_1),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_1),
.B(n_211),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_1),
.B(n_345),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_3),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_3),
.B(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_4),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_5),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_5),
.B(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_6),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_6),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_167),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_8),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_8),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_8),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_8),
.B(n_379),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_8),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_9),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_9),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_9),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_96),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_9),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_9),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_9),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_9),
.B(n_172),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_12),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_12),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_12),
.B(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_37),
.Y(n_45)
);

AND2x4_ASAP7_75t_SL g59 ( 
.A(n_15),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_15),
.B(n_102),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_15),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_15),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_15),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_16),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_16),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_16),
.B(n_223),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_327),
.B(n_432),
.C(n_443),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_226),
.B(n_279),
.C(n_326),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_179),
.B(n_225),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_134),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_73),
.C(n_109),
.Y(n_28)
);

XOR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_57),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_31),
.B(n_57),
.C(n_178),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_38),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_36),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_34),
.Y(n_307)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_38),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_38),
.B(n_163),
.C(n_165),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_39),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_53),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_41),
.A2(n_221),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_42),
.B(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_42),
.A2(n_107),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_42),
.B(n_45),
.Y(n_268)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_44),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_45),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_45),
.A2(n_258),
.B(n_265),
.Y(n_257)
);

OAI221xp5_ASAP7_75t_L g265 ( 
.A1(n_45),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.C(n_264),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_45),
.B(n_259),
.C(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_52),
.Y(n_144)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_55),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_56),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_67),
.C(n_71),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_58),
.A2(n_59),
.B1(n_82),
.B2(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_58),
.A2(n_59),
.B1(n_155),
.B2(n_156),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_58),
.B(n_82),
.C(n_358),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_58),
.B(n_156),
.C(n_387),
.Y(n_411)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_62)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_63),
.A2(n_71),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_70),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_71),
.B(n_313),
.C(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_89),
.C(n_103),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_82),
.C(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_80),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_80),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_82),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_82),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_82),
.B(n_261),
.C(n_305),
.Y(n_364)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_99),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_128),
.B2(n_133),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_129),
.C(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_118),
.C(n_122),
.Y(n_163)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_115),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_126),
.Y(n_359)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_161),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_135),
.B(n_162),
.C(n_177),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_138),
.C(n_150),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_150),
.Y(n_137)
);

XNOR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_145),
.Y(n_188)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_151),
.A2(n_152),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_152),
.B(n_311),
.C(n_322),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g412 ( 
.A1(n_155),
.A2(n_156),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_155),
.B(n_196),
.C(n_311),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_177),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_171),
.C(n_174),
.Y(n_199)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_224),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_224),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_202),
.B2(n_203),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_201),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_199),
.B2(n_200),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_192),
.Y(n_198)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_196),
.A2(n_197),
.B1(n_310),
.B2(n_311),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_196),
.A2(n_197),
.B1(n_259),
.B2(n_264),
.Y(n_429)
);

NOR3xp33_ASAP7_75t_L g444 ( 
.A(n_196),
.B(n_264),
.C(n_344),
.Y(n_444)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_216),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_241),
.C(n_242),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_210),
.C(n_214),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_214),
.B2(n_215),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_208),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_208),
.A2(n_214),
.B1(n_338),
.B2(n_343),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_208),
.B(n_343),
.C(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_217),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_218),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_233),
.B1(n_280),
.B2(n_323),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_234),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_256),
.Y(n_238)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_255),
.C(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_250),
.C(n_252),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_247),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_247),
.A2(n_250),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_247),
.A2(n_250),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_247),
.B(n_377),
.C(n_382),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_250),
.B(n_291),
.C(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_253),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_324),
.C(n_325),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_267),
.C(n_269),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_258)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_262),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2x1_ASAP7_75t_SL g326 ( 
.A(n_280),
.B(n_323),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_281),
.Y(n_394)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_300),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_285),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_286),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_299),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_289),
.Y(n_367)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_299),
.B(n_366),
.C(n_367),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_300),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_354),
.C(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_315),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_310),
.A2(n_311),
.B1(n_316),
.B2(n_317),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_312),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_398),
.C(n_423),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_390),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OA21x2_ASAP7_75t_SL g435 ( 
.A1(n_330),
.A2(n_436),
.B(n_437),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_368),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_332),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_356),
.C(n_365),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_353),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_349),
.B1(n_351),
.B2(n_352),
.Y(n_335)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_344),
.Y(n_336)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_338),
.Y(n_343)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_344),
.B(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_348),
.Y(n_410)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_349),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_350),
.B(n_441),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_350),
.B(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_352),
.C(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_363),
.C(n_364),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_396),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_368),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_421),
.C(n_422),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVxp33_ASAP7_75t_SL g421 ( 
.A(n_372),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_373),
.Y(n_422)
);

XOR2x2_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_374),
.B(n_384),
.C(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_380),
.B2(n_382),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_380),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_389),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_388),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_395),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.C(n_394),
.Y(n_391)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_L g439 ( 
.A1(n_399),
.A2(n_424),
.B(n_434),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_420),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_420),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_417),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_415),
.B2(n_416),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_415),
.C(n_418),
.Y(n_431)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_412),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_411),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_411),
.C(n_412),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_413),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_415),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_431),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_431),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_427),
.B(n_442),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_435),
.B(n_439),
.C(n_440),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);


endmodule