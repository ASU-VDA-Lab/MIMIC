module real_aes_8565_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g499 ( .A1(n_0), .A2(n_142), .B(n_500), .C(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_1), .B(n_161), .Y(n_503) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_3), .A2(n_128), .B(n_133), .C(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_4), .A2(n_123), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_5), .B(n_198), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_6), .A2(n_123), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_7), .B(n_161), .Y(n_227) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_8), .A2(n_146), .B(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_L g128 ( .A(n_9), .B(n_129), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_10), .A2(n_128), .B(n_133), .C(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g140 ( .A(n_11), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_12), .B(n_40), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_13), .B(n_138), .Y(n_175) );
INVx1_ASAP7_75t_L g121 ( .A(n_14), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_15), .B(n_198), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_16), .A2(n_141), .B(n_155), .C(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_17), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_18), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_19), .B(n_267), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_20), .A2(n_185), .B(n_186), .C(n_188), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_21), .A2(n_133), .B(n_202), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_22), .B(n_138), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_23), .B(n_138), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_24), .Y(n_209) );
INVx1_ASAP7_75t_L g197 ( .A(n_25), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_26), .A2(n_133), .B(n_202), .C(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_27), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_28), .Y(n_168) );
INVx1_ASAP7_75t_L g263 ( .A(n_29), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_30), .A2(n_123), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g126 ( .A(n_31), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_32), .A2(n_214), .B(n_435), .C(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_33), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_34), .A2(n_185), .B(n_223), .C(n_225), .Y(n_222) );
INVxp67_ASAP7_75t_L g264 ( .A(n_35), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_36), .B(n_459), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_37), .A2(n_133), .B(n_196), .C(n_202), .Y(n_195) );
CKINVDCx14_ASAP7_75t_R g221 ( .A(n_38), .Y(n_221) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_39), .A2(n_97), .B1(n_101), .B2(n_712), .C1(n_713), .C2(n_717), .Y(n_100) );
INVx1_ASAP7_75t_L g712 ( .A(n_39), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_41), .A2(n_137), .B(n_139), .C(n_142), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_42), .B(n_258), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_43), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_44), .A2(n_99), .B1(n_721), .B2(n_730), .C1(n_738), .C2(n_744), .Y(n_98) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_44), .A2(n_427), .B1(n_720), .B2(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_44), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_45), .B(n_198), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_46), .B(n_123), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_47), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_48), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_49), .A2(n_214), .B(n_435), .C(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g502 ( .A(n_50), .Y(n_502) );
INVx1_ASAP7_75t_L g437 ( .A(n_51), .Y(n_437) );
INVx1_ASAP7_75t_L g183 ( .A(n_52), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_53), .B(n_123), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_54), .Y(n_483) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_55), .Y(n_131) );
INVx1_ASAP7_75t_L g129 ( .A(n_56), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_57), .B(n_123), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_58), .B(n_161), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_59), .A2(n_201), .B(n_448), .C(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g120 ( .A(n_60), .Y(n_120) );
INVx1_ASAP7_75t_SL g224 ( .A(n_61), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_62), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_63), .B(n_198), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_64), .B(n_161), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_65), .B(n_141), .Y(n_512) );
INVx1_ASAP7_75t_L g212 ( .A(n_66), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_67), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_68), .B(n_174), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_69), .A2(n_133), .B(n_214), .C(n_488), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_70), .Y(n_446) );
INVx1_ASAP7_75t_L g725 ( .A(n_71), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_72), .A2(n_123), .B(n_130), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_73), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_74), .A2(n_123), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_75), .A2(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g153 ( .A(n_76), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_77), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_78), .B(n_173), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_79), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_80), .A2(n_123), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g156 ( .A(n_81), .Y(n_156) );
INVx2_ASAP7_75t_L g118 ( .A(n_82), .Y(n_118) );
INVx1_ASAP7_75t_L g172 ( .A(n_83), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_84), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_85), .B(n_138), .Y(n_513) );
INVx2_ASAP7_75t_L g107 ( .A(n_86), .Y(n_107) );
OR2x2_ASAP7_75t_L g426 ( .A(n_86), .B(n_108), .Y(n_426) );
OR2x2_ASAP7_75t_L g729 ( .A(n_86), .B(n_716), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_87), .A2(n_133), .B(n_211), .C(n_214), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_88), .B(n_123), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_89), .Y(n_470) );
INVxp67_ASAP7_75t_L g450 ( .A(n_90), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_91), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g187 ( .A(n_92), .Y(n_187) );
INVx1_ASAP7_75t_L g489 ( .A(n_93), .Y(n_489) );
INVx1_ASAP7_75t_L g509 ( .A(n_94), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_95), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g440 ( .A(n_96), .B(n_117), .Y(n_440) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_111), .B1(n_423), .B2(n_427), .Y(n_102) );
AOI22x1_ASAP7_75t_SL g718 ( .A1(n_103), .A2(n_423), .B1(n_719), .B2(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_107), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_108), .Y(n_716) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx2_ASAP7_75t_L g719 ( .A(n_111), .Y(n_719) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_353), .Y(n_111) );
NAND5xp2_ASAP7_75t_L g112 ( .A(n_113), .B(n_268), .C(n_300), .D(n_317), .E(n_340), .Y(n_112) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_191), .B1(n_228), .B2(n_232), .C(n_236), .Y(n_113) );
INVx1_ASAP7_75t_L g380 ( .A(n_114), .Y(n_380) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_163), .Y(n_114) );
AND3x2_ASAP7_75t_L g355 ( .A(n_115), .B(n_165), .C(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_148), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_116), .B(n_234), .Y(n_233) );
BUFx3_ASAP7_75t_L g243 ( .A(n_116), .Y(n_243) );
AND2x2_ASAP7_75t_L g247 ( .A(n_116), .B(n_179), .Y(n_247) );
INVx2_ASAP7_75t_L g277 ( .A(n_116), .Y(n_277) );
OR2x2_ASAP7_75t_L g288 ( .A(n_116), .B(n_180), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_116), .B(n_164), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_116), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g367 ( .A(n_116), .B(n_180), .Y(n_367) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_145), .Y(n_116) );
INVx1_ASAP7_75t_L g166 ( .A(n_117), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_117), .A2(n_169), .B(n_194), .C(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g217 ( .A(n_117), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_117), .A2(n_433), .B(n_434), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_117), .A2(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x2_ASAP7_75t_L g147 ( .A(n_118), .B(n_119), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
BUFx2_ASAP7_75t_L g258 ( .A(n_123), .Y(n_258) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_128), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_124), .B(n_128), .Y(n_169) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
INVx1_ASAP7_75t_L g201 ( .A(n_125), .Y(n_201) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
INVx1_ASAP7_75t_L g189 ( .A(n_126), .Y(n_189) );
INVx1_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_127), .Y(n_138) );
INVx3_ASAP7_75t_L g141 ( .A(n_127), .Y(n_141) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_127), .Y(n_158) );
INVx1_ASAP7_75t_L g459 ( .A(n_127), .Y(n_459) );
INVx4_ASAP7_75t_SL g144 ( .A(n_128), .Y(n_144) );
BUFx3_ASAP7_75t_L g202 ( .A(n_128), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_132), .B(n_136), .C(n_144), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_SL g152 ( .A1(n_132), .A2(n_144), .B(n_153), .C(n_154), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_SL g182 ( .A1(n_132), .A2(n_144), .B(n_183), .C(n_184), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_132), .A2(n_144), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_132), .A2(n_144), .B(n_260), .C(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g435 ( .A(n_132), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_132), .A2(n_144), .B(n_446), .C(n_447), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_132), .A2(n_144), .B(n_498), .C(n_499), .Y(n_497) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx3_ASAP7_75t_L g143 ( .A(n_134), .Y(n_143) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_134), .Y(n_226) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx5_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
INVx2_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g159 ( .A(n_143), .Y(n_159) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_143), .Y(n_439) );
INVx1_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_146), .Y(n_150) );
INVx4_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_146), .A2(n_455), .B(n_456), .Y(n_454) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g255 ( .A(n_147), .Y(n_255) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_148), .Y(n_246) );
AND2x2_ASAP7_75t_L g308 ( .A(n_148), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_148), .B(n_164), .Y(n_327) );
INVx1_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g235 ( .A(n_149), .B(n_164), .Y(n_235) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_149), .Y(n_242) );
AND2x2_ASAP7_75t_L g294 ( .A(n_149), .B(n_180), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_149), .B(n_163), .C(n_277), .Y(n_319) );
AND2x2_ASAP7_75t_L g384 ( .A(n_149), .B(n_165), .Y(n_384) );
AND2x2_ASAP7_75t_L g418 ( .A(n_149), .B(n_164), .Y(n_418) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_160), .Y(n_149) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_150), .A2(n_181), .B(n_190), .Y(n_180) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_150), .A2(n_219), .B(n_227), .Y(n_218) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_150), .A2(n_444), .B(n_451), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_157), .B(n_187), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_157), .A2(n_198), .B1(n_263), .B2(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g448 ( .A(n_157), .Y(n_448) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_161), .A2(n_496), .B(n_503), .Y(n_495) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_162), .B(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_162), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_162), .A2(n_208), .B(n_215), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_162), .B(n_473), .Y(n_472) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_162), .A2(n_486), .B(n_493), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_162), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_162), .A2(n_508), .B(n_514), .Y(n_507) );
INVxp67_ASAP7_75t_L g244 ( .A(n_163), .Y(n_244) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_179), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_164), .B(n_277), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_164), .B(n_308), .Y(n_316) );
AND2x2_ASAP7_75t_L g366 ( .A(n_164), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_164), .Y(n_394) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g301 ( .A(n_165), .B(n_294), .Y(n_301) );
BUFx3_ASAP7_75t_L g333 ( .A(n_165), .Y(n_333) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_177), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_166), .B(n_483), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_169), .A2(n_209), .B(n_210), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_169), .A2(n_509), .B(n_510), .Y(n_508) );
O2A1O1Ixp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_175), .C(n_176), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_173), .A2(n_176), .B(n_212), .C(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g436 ( .A1(n_173), .A2(n_437), .B(n_438), .C(n_439), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_173), .A2(n_439), .B(n_470), .C(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g309 ( .A(n_179), .Y(n_309) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_185), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_185), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g461 ( .A(n_188), .Y(n_461) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_191), .A2(n_369), .B1(n_371), .B2(n_372), .Y(n_368) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_205), .Y(n_191) );
AND2x2_ASAP7_75t_L g228 ( .A(n_192), .B(n_229), .Y(n_228) );
INVx3_ASAP7_75t_SL g239 ( .A(n_192), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_192), .B(n_272), .Y(n_304) );
OR2x2_ASAP7_75t_L g323 ( .A(n_192), .B(n_206), .Y(n_323) );
AND2x2_ASAP7_75t_L g328 ( .A(n_192), .B(n_280), .Y(n_328) );
AND2x2_ASAP7_75t_L g331 ( .A(n_192), .B(n_273), .Y(n_331) );
AND2x2_ASAP7_75t_L g343 ( .A(n_192), .B(n_218), .Y(n_343) );
AND2x2_ASAP7_75t_L g359 ( .A(n_192), .B(n_207), .Y(n_359) );
AND2x4_ASAP7_75t_L g362 ( .A(n_192), .B(n_230), .Y(n_362) );
OR2x2_ASAP7_75t_L g379 ( .A(n_192), .B(n_315), .Y(n_379) );
OR2x2_ASAP7_75t_L g410 ( .A(n_192), .B(n_252), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_192), .B(n_338), .Y(n_412) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_203), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .C(n_200), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_198), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g500 ( .A(n_198), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_200), .A2(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_201), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g286 ( .A(n_205), .B(n_250), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_205), .B(n_273), .Y(n_405) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_218), .Y(n_205) );
AND2x2_ASAP7_75t_L g238 ( .A(n_206), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g272 ( .A(n_206), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g280 ( .A(n_206), .B(n_252), .Y(n_280) );
AND2x2_ASAP7_75t_L g298 ( .A(n_206), .B(n_230), .Y(n_298) );
OR2x2_ASAP7_75t_L g315 ( .A(n_206), .B(n_273), .Y(n_315) );
INVx2_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g231 ( .A(n_207), .Y(n_231) );
AND2x2_ASAP7_75t_L g338 ( .A(n_207), .B(n_218), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
INVx1_ASAP7_75t_L g267 ( .A(n_217), .Y(n_267) );
INVx2_ASAP7_75t_L g230 ( .A(n_218), .Y(n_230) );
INVx1_ASAP7_75t_L g350 ( .A(n_218), .Y(n_350) );
AND2x2_ASAP7_75t_L g400 ( .A(n_218), .B(n_239), .Y(n_400) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_226), .Y(n_491) );
AND2x2_ASAP7_75t_L g249 ( .A(n_229), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g284 ( .A(n_229), .B(n_239), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_229), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x2_ASAP7_75t_L g271 ( .A(n_230), .B(n_239), .Y(n_271) );
OR2x2_ASAP7_75t_L g387 ( .A(n_231), .B(n_361), .Y(n_387) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_234), .B(n_367), .Y(n_373) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OAI32xp33_ASAP7_75t_L g329 ( .A1(n_235), .A2(n_330), .A3(n_332), .B1(n_334), .B2(n_335), .Y(n_329) );
OR2x2_ASAP7_75t_L g346 ( .A(n_235), .B(n_288), .Y(n_346) );
OAI21xp33_ASAP7_75t_SL g371 ( .A1(n_235), .A2(n_245), .B(n_276), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_240), .B1(n_245), .B2(n_248), .Y(n_236) );
INVxp33_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_238), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_239), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g297 ( .A(n_239), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g397 ( .A(n_239), .B(n_338), .Y(n_397) );
OR2x2_ASAP7_75t_L g421 ( .A(n_239), .B(n_315), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_240), .A2(n_303), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_244), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g281 ( .A(n_242), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_242), .B(n_247), .Y(n_299) );
AND2x2_ASAP7_75t_L g321 ( .A(n_243), .B(n_294), .Y(n_321) );
INVx1_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
OR2x2_ASAP7_75t_L g339 ( .A(n_243), .B(n_273), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_246), .B(n_288), .Y(n_287) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_247), .A2(n_270), .B1(n_275), .B2(n_279), .Y(n_269) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_250), .A2(n_312), .B1(n_319), .B2(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g396 ( .A(n_250), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_252), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g415 ( .A(n_252), .B(n_298), .Y(n_415) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .B(n_265), .Y(n_252) );
INVx1_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_255), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_257), .A2(n_266), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AOI21xp5_ASAP7_75t_SL g476 ( .A1(n_267), .A2(n_477), .B(n_478), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_281), .B1(n_282), .B2(n_287), .C(n_289), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_271), .B(n_273), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_271), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g290 ( .A(n_272), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_272), .A2(n_378), .B(n_379), .C(n_380), .Y(n_377) );
AND2x2_ASAP7_75t_L g382 ( .A(n_272), .B(n_362), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_SL g420 ( .A1(n_272), .A2(n_361), .B(n_421), .C(n_422), .Y(n_420) );
BUFx3_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_276), .B(n_333), .Y(n_376) );
AOI211xp5_ASAP7_75t_L g395 ( .A1(n_276), .A2(n_396), .B(n_398), .C(n_404), .Y(n_395) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVxp67_ASAP7_75t_L g356 ( .A(n_278), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_280), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AOI211xp5_ASAP7_75t_L g300 ( .A1(n_284), .A2(n_301), .B(n_302), .C(n_310), .Y(n_300) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g385 ( .A(n_288), .Y(n_385) );
OR2x2_ASAP7_75t_L g402 ( .A(n_288), .B(n_332), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_296), .B2(n_299), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g302 ( .A1(n_291), .A2(n_303), .B1(n_304), .B2(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
OR2x2_ASAP7_75t_L g389 ( .A(n_293), .B(n_333), .Y(n_389) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g344 ( .A(n_294), .B(n_334), .Y(n_344) );
INVx1_ASAP7_75t_L g352 ( .A(n_295), .Y(n_352) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_298), .B(n_312), .Y(n_360) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_308), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g417 ( .A(n_309), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B(n_316), .Y(n_310) );
INVx1_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_312), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_312), .B(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_312), .B(n_338), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_312), .B(n_359), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_312), .A2(n_322), .B(n_362), .C(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_322), .B1(n_324), .B2(n_328), .C(n_329), .Y(n_317) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_326), .B(n_334), .Y(n_408) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_328), .A2(n_343), .B(n_345), .C(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_331), .B(n_338), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_332), .B(n_385), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_333), .Y(n_332) );
INVxp33_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AOI21xp33_ASAP7_75t_SL g348 ( .A1(n_337), .A2(n_349), .B(n_351), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_337), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_338), .B(n_392), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_345), .B2(n_347), .C(n_348), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_344), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
NAND5xp2_ASAP7_75t_L g353 ( .A(n_354), .B(n_381), .C(n_395), .D(n_406), .E(n_419), .Y(n_353) );
AOI211xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_364), .C(n_377), .Y(n_354) );
INVx2_ASAP7_75t_SL g401 ( .A(n_355), .Y(n_401) );
NAND4xp25_ASAP7_75t_SL g357 ( .A(n_358), .B(n_360), .C(n_361), .D(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_363), .A2(n_365), .B(n_368), .C(n_374), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_407), .B1(n_409), .B2(n_411), .C(n_413), .Y(n_406) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_383), .B1(n_386), .B2(n_388), .C(n_390), .Y(n_381) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_412), .B1(n_414), .B2(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx4_ASAP7_75t_L g720 ( .A(n_427), .Y(n_720) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR5x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_585), .C(n_663), .D(n_687), .E(n_704), .Y(n_428) );
OAI211xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_462), .B(n_504), .C(n_562), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_441), .Y(n_430) );
AND2x2_ASAP7_75t_L g516 ( .A(n_431), .B(n_443), .Y(n_516) );
INVx5_ASAP7_75t_SL g544 ( .A(n_431), .Y(n_544) );
AND2x2_ASAP7_75t_L g580 ( .A(n_431), .B(n_565), .Y(n_580) );
OR2x2_ASAP7_75t_L g619 ( .A(n_431), .B(n_442), .Y(n_619) );
OR2x2_ASAP7_75t_L g650 ( .A(n_431), .B(n_541), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_431), .B(n_554), .Y(n_686) );
AND2x2_ASAP7_75t_L g698 ( .A(n_431), .B(n_541), .Y(n_698) );
OR2x6_ASAP7_75t_L g431 ( .A(n_432), .B(n_440), .Y(n_431) );
AND2x2_ASAP7_75t_L g697 ( .A(n_441), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g560 ( .A(n_442), .B(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_452), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_443), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_443), .Y(n_553) );
INVx3_ASAP7_75t_L g568 ( .A(n_443), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_443), .B(n_452), .Y(n_592) );
OR2x2_ASAP7_75t_L g601 ( .A(n_443), .B(n_544), .Y(n_601) );
AND2x2_ASAP7_75t_L g605 ( .A(n_443), .B(n_565), .Y(n_605) );
AND2x2_ASAP7_75t_L g611 ( .A(n_443), .B(n_612), .Y(n_611) );
INVxp67_ASAP7_75t_L g648 ( .A(n_443), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_443), .B(n_507), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_448), .A2(n_489), .B(n_490), .C(n_491), .Y(n_488) );
OR2x2_ASAP7_75t_L g554 ( .A(n_452), .B(n_507), .Y(n_554) );
AND2x2_ASAP7_75t_L g565 ( .A(n_452), .B(n_541), .Y(n_565) );
AND2x2_ASAP7_75t_L g577 ( .A(n_452), .B(n_568), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_452), .B(n_507), .Y(n_600) );
INVx1_ASAP7_75t_SL g612 ( .A(n_452), .Y(n_612) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g506 ( .A(n_453), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_453), .B(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B(n_461), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_461), .A2(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
AND2x2_ASAP7_75t_L g525 ( .A(n_464), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_464), .B(n_484), .Y(n_529) );
AND2x2_ASAP7_75t_L g532 ( .A(n_464), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_464), .B(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g557 ( .A(n_464), .B(n_548), .Y(n_557) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_464), .Y(n_576) );
AND2x2_ASAP7_75t_L g597 ( .A(n_464), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g607 ( .A(n_464), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g653 ( .A(n_464), .B(n_536), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_464), .B(n_559), .Y(n_680) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g550 ( .A(n_465), .Y(n_550) );
AND2x2_ASAP7_75t_L g616 ( .A(n_465), .B(n_548), .Y(n_616) );
AND2x2_ASAP7_75t_L g700 ( .A(n_465), .B(n_568), .Y(n_700) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_474), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_474), .Y(n_689) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
AND2x2_ASAP7_75t_L g519 ( .A(n_475), .B(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g528 ( .A(n_475), .B(n_526), .Y(n_528) );
INVx5_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
AND2x2_ASAP7_75t_L g559 ( .A(n_475), .B(n_495), .Y(n_559) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_475), .Y(n_596) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
INVx1_ASAP7_75t_L g637 ( .A(n_484), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_484), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g670 ( .A(n_484), .B(n_536), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_484), .A2(n_593), .B(n_700), .C(n_701), .Y(n_699) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .Y(n_484) );
BUFx2_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx2_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_492), .Y(n_486) );
INVx2_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
AND2x2_ASAP7_75t_L g533 ( .A(n_495), .B(n_524), .Y(n_533) );
AND2x2_ASAP7_75t_L g624 ( .A(n_495), .B(n_536), .Y(n_624) );
AOI211x1_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_517), .B(n_530), .C(n_555), .Y(n_504) );
INVx1_ASAP7_75t_L g621 ( .A(n_505), .Y(n_621) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_516), .Y(n_505) );
INVx5_ASAP7_75t_SL g541 ( .A(n_507), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_507), .B(n_611), .Y(n_610) );
AOI311xp33_ASAP7_75t_L g629 ( .A1(n_507), .A2(n_630), .A3(n_632), .B(n_633), .C(n_639), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_507), .A2(n_577), .B(n_665), .C(n_668), .Y(n_664) );
INVxp67_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
NAND4xp25_ASAP7_75t_SL g517 ( .A(n_518), .B(n_521), .C(n_527), .D(n_529), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_518), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g575 ( .A(n_519), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_522), .B(n_528), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_522), .B(n_535), .Y(n_655) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_523), .B(n_536), .Y(n_673) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g548 ( .A(n_524), .Y(n_548) );
INVxp67_ASAP7_75t_L g583 ( .A(n_525), .Y(n_583) );
AND2x4_ASAP7_75t_L g535 ( .A(n_526), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g609 ( .A(n_526), .B(n_548), .Y(n_609) );
INVx1_ASAP7_75t_L g636 ( .A(n_526), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_526), .B(n_623), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_527), .B(n_597), .Y(n_617) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_528), .B(n_550), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_528), .B(n_597), .Y(n_696) );
INVx1_ASAP7_75t_L g707 ( .A(n_529), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_534), .B(n_537), .C(n_545), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g549 ( .A(n_533), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g587 ( .A(n_533), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g569 ( .A(n_534), .Y(n_569) );
AND2x2_ASAP7_75t_L g546 ( .A(n_535), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_535), .B(n_597), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_535), .B(n_616), .Y(n_640) );
OR2x2_ASAP7_75t_L g556 ( .A(n_536), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g588 ( .A(n_536), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_536), .B(n_548), .Y(n_603) );
AND2x2_ASAP7_75t_L g660 ( .A(n_536), .B(n_616), .Y(n_660) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_536), .Y(n_667) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_538), .A2(n_550), .B1(n_672), .B2(n_674), .C(n_677), .Y(n_671) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g561 ( .A(n_541), .B(n_544), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_541), .B(n_611), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_541), .B(n_568), .Y(n_676) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g661 ( .A(n_543), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g675 ( .A(n_543), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_544), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g572 ( .A(n_544), .B(n_565), .Y(n_572) );
AND2x2_ASAP7_75t_L g642 ( .A(n_544), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_544), .B(n_591), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_544), .B(n_692), .Y(n_691) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_549), .B(n_551), .Y(n_545) );
INVx2_ASAP7_75t_L g578 ( .A(n_546), .Y(n_578) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g598 ( .A(n_548), .Y(n_598) );
OR2x2_ASAP7_75t_L g602 ( .A(n_550), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g705 ( .A(n_550), .B(n_673), .Y(n_705) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AOI21xp33_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_558), .B(n_560), .Y(n_555) );
INVx1_ASAP7_75t_L g709 ( .A(n_556), .Y(n_709) );
INVx2_ASAP7_75t_SL g623 ( .A(n_557), .Y(n_623) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_560), .A2(n_641), .B(n_705), .C(n_706), .Y(n_704) );
OAI322xp33_ASAP7_75t_SL g573 ( .A1(n_561), .A2(n_574), .A3(n_577), .B1(n_578), .B2(n_579), .C1(n_581), .C2(n_584), .Y(n_573) );
INVx2_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_569), .B1(n_570), .B2(n_572), .C(n_573), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI22xp33_ASAP7_75t_SL g639 ( .A1(n_564), .A2(n_640), .B1(n_641), .B2(n_644), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_565), .B(n_568), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_565), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g638 ( .A(n_567), .B(n_600), .Y(n_638) );
INVx1_ASAP7_75t_L g628 ( .A(n_568), .Y(n_628) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_572), .A2(n_682), .B(n_684), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g606 ( .A1(n_574), .A2(n_607), .B(n_610), .Y(n_606) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp67_ASAP7_75t_SL g635 ( .A(n_576), .B(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_576), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g692 ( .A(n_577), .Y(n_692) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_613), .C(n_629), .D(n_645), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_594), .C(n_606), .Y(n_586) );
INVx1_ASAP7_75t_L g678 ( .A(n_587), .Y(n_678) );
AND2x2_ASAP7_75t_L g626 ( .A(n_588), .B(n_609), .Y(n_626) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_593), .B(n_628), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B1(n_602), .B2(n_604), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_596), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_597), .A2(n_636), .B(n_659), .C(n_661), .Y(n_658) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g643 ( .A(n_600), .Y(n_643) );
INVx1_ASAP7_75t_L g703 ( .A(n_601), .Y(n_703) );
NAND2xp33_ASAP7_75t_SL g693 ( .A(n_602), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g632 ( .A(n_611), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B(n_618), .C(n_620), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_625), .B2(n_627), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_623), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_628), .B(n_649), .Y(n_711) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI21xp33_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_637), .B(n_638), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_651), .B1(n_654), .B2(n_656), .C(n_658), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_661), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_677) );
NAND3xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_671), .C(n_681), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B(n_690), .C(n_699), .Y(n_687) );
INVx1_ASAP7_75t_L g708 ( .A(n_688), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_695), .B2(n_697), .Y(n_690) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
NAND2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
NOR2xp33_ASAP7_75t_SL g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_SL g743 ( .A(n_724), .Y(n_743) );
INVx1_ASAP7_75t_L g742 ( .A(n_726), .Y(n_742) );
OA21x2_ASAP7_75t_L g745 ( .A1(n_726), .A2(n_743), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g733 ( .A(n_727), .Y(n_733) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g737 ( .A(n_729), .Y(n_737) );
BUFx2_ASAP7_75t_L g746 ( .A(n_729), .Y(n_746) );
OAI21xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_733), .B(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
CKINVDCx6p67_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
endmodule