module fake_netlist_6_3726_n_1850 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1850);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1850;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g178 ( 
.A(n_14),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_32),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_76),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_10),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_173),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_77),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_14),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_96),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_110),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_88),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_71),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_9),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_54),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_4),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_70),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_32),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_20),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_30),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_49),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_52),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_6),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_74),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_13),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_97),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_169),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_150),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_23),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_83),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_44),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_155),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_55),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_69),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_73),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_162),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_4),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_154),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_161),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_153),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_151),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_95),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_9),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_56),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_33),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_23),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_79),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_112),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_164),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_111),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_34),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_44),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_106),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_61),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_103),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_60),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_168),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_80),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_124),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_113),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_17),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_115),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_133),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_94),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_145),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_85),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_123),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_135),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_140),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_108),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_24),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_42),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_159),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_68),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_89),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_148),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_137),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_2),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_48),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_165),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_52),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_139),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_18),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_22),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_21),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_64),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_47),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_36),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_141),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_147),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_131),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_3),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_177),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_170),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_28),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_39),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_101),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_142),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_125),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_31),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_86),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_122),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_58),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_3),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_33),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_45),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_61),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_99),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_11),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_0),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_41),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_158),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_0),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_92),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_1),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_130),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_98),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_5),
.Y(n_335)
);

BUFx8_ASAP7_75t_SL g336 ( 
.A(n_65),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_172),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_50),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_116),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_1),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_156),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_81),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_93),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_49),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_43),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_24),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_117),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_51),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_59),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_62),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_54),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_22),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_27),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_42),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_202),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_181),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_179),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_180),
.B(n_6),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_187),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_187),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_200),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_182),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_186),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_293),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_185),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_190),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_200),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_180),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_209),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_222),
.B(n_7),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_203),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_304),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_213),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_304),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_214),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_218),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_283),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_310),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_227),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_203),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_225),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_220),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_206),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_331),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_206),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_178),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_336),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_208),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_228),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_183),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_215),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_208),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_225),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_232),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_178),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_184),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_236),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_210),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_189),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_210),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_211),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_246),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_211),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_248),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_256),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_257),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_224),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_273),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_259),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_194),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_284),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_224),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_215),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_226),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_226),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_233),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_233),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_234),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_234),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_195),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_197),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_284),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_R g430 ( 
.A(n_198),
.B(n_105),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_240),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_205),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_243),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_265),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_221),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_207),
.B(n_7),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_273),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_243),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_277),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_251),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_R g442 ( 
.A(n_229),
.B(n_107),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_255),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_251),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_192),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_394),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_397),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_222),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_388),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

AND3x2_ASAP7_75t_L g452 ( 
.A(n_372),
.B(n_267),
.C(n_230),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_362),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_362),
.B(n_192),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_403),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_376),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_355),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_376),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_406),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_378),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_417),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_398),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_427),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_420),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_364),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_357),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_368),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_402),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_415),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_383),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_415),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_279),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_SL g481 ( 
.A(n_359),
.B(n_204),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_428),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_357),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_355),
.B(n_366),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_356),
.B(n_223),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_374),
.B(n_223),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_358),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_437),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_360),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_430),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_384),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_365),
.B(n_278),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_361),
.B(n_307),
.Y(n_494)
);

AND3x1_ASAP7_75t_L g495 ( 
.A(n_386),
.B(n_216),
.C(n_207),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_437),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_363),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_370),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_375),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_433),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_387),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_399),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_R g506 ( 
.A(n_365),
.B(n_285),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_367),
.B(n_307),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_385),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_410),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_367),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_279),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_421),
.B(n_255),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_422),
.B(n_235),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_369),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_436),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_369),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_371),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_371),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_L g523 ( 
.A1(n_496),
.A2(n_400),
.B1(n_418),
.B2(n_429),
.Y(n_523)
);

AND3x2_ASAP7_75t_L g524 ( 
.A(n_457),
.B(n_271),
.C(n_230),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_496),
.A2(n_386),
.B1(n_193),
.B2(n_330),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_450),
.B(n_373),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_520),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_456),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_496),
.B(n_199),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_488),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_258),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_450),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_488),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_373),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_457),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_454),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_461),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_490),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_499),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_451),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_499),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_495),
.A2(n_270),
.B1(n_391),
.B2(n_340),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_451),
.B(n_423),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_513),
.B(n_199),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_489),
.A2(n_322),
.B1(n_351),
.B2(n_441),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_377),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_454),
.B(n_424),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_454),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_451),
.B(n_425),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_451),
.B(n_426),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_445),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_462),
.Y(n_561)
);

INVx4_ASAP7_75t_SL g562 ( 
.A(n_486),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_486),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_462),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_454),
.B(n_431),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_513),
.B(n_254),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_517),
.B(n_377),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_513),
.B(n_254),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

BUFx8_ASAP7_75t_SL g570 ( 
.A(n_469),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_470),
.B(n_281),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_456),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_445),
.B(n_258),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_470),
.B(n_281),
.Y(n_576)
);

BUFx4f_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_489),
.A2(n_351),
.B1(n_322),
.B2(n_439),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_445),
.B(n_261),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_466),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_480),
.B(n_516),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_448),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_486),
.B(n_219),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_503),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_466),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_503),
.B(n_219),
.Y(n_589)
);

INVx8_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_508),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_491),
.B(n_432),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_480),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_466),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_447),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_447),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_480),
.B(n_380),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_468),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_509),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_449),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_481),
.A2(n_434),
.B1(n_320),
.B2(n_348),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_518),
.B(n_380),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_503),
.Y(n_605)
);

INVx6_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_466),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_468),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_473),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_506),
.A2(n_404),
.B1(n_440),
.B2(n_435),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_503),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_495),
.B(n_219),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_518),
.A2(n_411),
.B1(n_440),
.B2(n_435),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_516),
.B(n_261),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_483),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_522),
.B(n_382),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_468),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_483),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_516),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_515),
.A2(n_300),
.B1(n_231),
.B2(n_217),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_515),
.B(n_268),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_475),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_522),
.B(n_382),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_493),
.B(n_389),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_389),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_453),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_446),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_453),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_497),
.B(n_396),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_491),
.B(n_396),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_458),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_458),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_460),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_485),
.B(n_401),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_491),
.B(n_401),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_475),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_452),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_460),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_475),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_484),
.B(n_216),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_494),
.A2(n_260),
.B1(n_262),
.B2(n_250),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_497),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_497),
.B(n_404),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_498),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_449),
.B(n_268),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_477),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_409),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_477),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_498),
.B(n_274),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_501),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_476),
.B(n_409),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_492),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_452),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_494),
.B(n_274),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_511),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_501),
.A2(n_250),
.B1(n_300),
.B2(n_245),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_501),
.B(n_411),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_491),
.B(n_412),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_502),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_502),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_502),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_519),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_504),
.B(n_412),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_504),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_507),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_507),
.B(n_282),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_507),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_530),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_600),
.A2(n_514),
.B(n_512),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_560),
.B(n_583),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_533),
.B(n_413),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_628),
.B(n_413),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_570),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_593),
.B(n_416),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_543),
.B(n_512),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_625),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_583),
.B(n_464),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_643),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_583),
.B(n_464),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_546),
.A2(n_514),
.B(n_512),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_525),
.B(n_247),
.C(n_467),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_514),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_551),
.B(n_282),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_628),
.B(n_286),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_539),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_532),
.A2(n_327),
.B1(n_260),
.B2(n_262),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_637),
.B(n_286),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_606),
.A2(n_306),
.B1(n_341),
.B2(n_337),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_541),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_637),
.B(n_191),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_606),
.A2(n_288),
.B1(n_287),
.B2(n_306),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_532),
.B(n_287),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_532),
.B(n_606),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_567),
.A2(n_325),
.B1(n_337),
.B2(n_333),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_632),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_535),
.B(n_467),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_611),
.B(n_459),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_526),
.B(n_463),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_647),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_537),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_542),
.Y(n_709)
);

INVx6_ASAP7_75t_L g710 ( 
.A(n_668),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_537),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_532),
.B(n_288),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_544),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_537),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_549),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_532),
.B(n_325),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_662),
.A2(n_333),
.B(n_341),
.C(n_478),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_535),
.B(n_465),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_643),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_627),
.A2(n_624),
.B1(n_552),
.B2(n_662),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_555),
.A2(n_472),
.B(n_471),
.Y(n_721)
);

BUFx8_ASAP7_75t_L g722 ( 
.A(n_536),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_R g723 ( 
.A(n_584),
.B(n_482),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_590),
.B(n_217),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_578),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_669),
.B(n_472),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_591),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_552),
.B(n_474),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_575),
.B(n_237),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_523),
.A2(n_296),
.B1(n_245),
.B2(n_313),
.C(n_299),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_552),
.B(n_474),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_643),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_642),
.B(n_478),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_597),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_579),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_642),
.B(n_479),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_622),
.B(n_196),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_579),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_665),
.B(n_479),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_665),
.B(n_269),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_670),
.B(n_275),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_615),
.A2(n_321),
.B1(n_296),
.B2(n_299),
.Y(n_742)
);

OAI221xp5_ASAP7_75t_L g743 ( 
.A1(n_645),
.A2(n_623),
.B1(n_601),
.B2(n_580),
.C(n_550),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_595),
.Y(n_744)
);

O2A1O1Ixp5_ASAP7_75t_L g745 ( 
.A1(n_529),
.A2(n_313),
.B(n_327),
.C(n_321),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_668),
.B(n_219),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_617),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_595),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_602),
.B(n_291),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_602),
.B(n_619),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_617),
.A2(n_231),
.B(n_320),
.C(n_346),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_627),
.B(n_500),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_619),
.B(n_292),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_626),
.B(n_295),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_626),
.B(n_298),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_644),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_668),
.B(n_238),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_571),
.B(n_302),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_559),
.B(n_629),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_616),
.B(n_442),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_571),
.B(n_303),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_554),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_599),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_608),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_554),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_618),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_576),
.B(n_308),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_239),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_633),
.B(n_638),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_634),
.B(n_241),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_635),
.B(n_242),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_636),
.B(n_565),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_529),
.B(n_244),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_639),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_590),
.B(n_346),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_623),
.A2(n_349),
.B1(n_352),
.B2(n_348),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_621),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_SL g778 ( 
.A(n_601),
.B(n_354),
.C(n_353),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_547),
.B(n_249),
.Y(n_779)
);

AND2x4_ASAP7_75t_SL g780 ( 
.A(n_667),
.B(n_215),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_554),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_558),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_615),
.B(n_352),
.C(n_349),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_596),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_547),
.B(n_252),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_596),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_576),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_624),
.A2(n_315),
.B1(n_347),
.B2(n_253),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_617),
.A2(n_318),
.B(n_272),
.C(n_276),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_598),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_641),
.B(n_311),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_658),
.B(n_651),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_566),
.A2(n_280),
.B1(n_266),
.B2(n_290),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_663),
.B(n_264),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_598),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_566),
.B(n_312),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_568),
.B(n_294),
.Y(n_797)
);

OAI221xp5_ASAP7_75t_L g798 ( 
.A1(n_645),
.A2(n_350),
.B1(n_345),
.B2(n_344),
.C(n_317),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_644),
.B(n_610),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_527),
.B(n_215),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_568),
.B(n_323),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_609),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_644),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_570),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_SL g805 ( 
.A(n_545),
.B(n_324),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_673),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_527),
.B(n_326),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_624),
.B(n_301),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_624),
.B(n_305),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_624),
.B(n_309),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_SL g811 ( 
.A(n_527),
.B(n_289),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_657),
.B(n_328),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_575),
.A2(n_343),
.B1(n_342),
.B2(n_339),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_575),
.B(n_334),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_550),
.A2(n_329),
.B1(n_319),
.B2(n_314),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_609),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_673),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_659),
.A2(n_219),
.B1(n_263),
.B2(n_297),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_654),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_524),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_575),
.A2(n_316),
.B1(n_297),
.B2(n_289),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_575),
.B(n_263),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_581),
.A2(n_316),
.B1(n_297),
.B2(n_289),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_655),
.B(n_338),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_585),
.A2(n_316),
.B(n_297),
.C(n_289),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_654),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_667),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_581),
.B(n_263),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_655),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_646),
.A2(n_335),
.B1(n_332),
.B2(n_263),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_581),
.B(n_263),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_648),
.B(n_316),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_654),
.B(n_171),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_580),
.B(n_8),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_581),
.B(n_143),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_581),
.B(n_659),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_592),
.B(n_138),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_620),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_556),
.B(n_8),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_664),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_666),
.B(n_10),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_838),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_708),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_698),
.B(n_659),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_790),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_584),
.C(n_661),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_690),
.A2(n_586),
.B(n_569),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_750),
.B(n_659),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_772),
.A2(n_586),
.B(n_569),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_726),
.B(n_659),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_678),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_819),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_819),
.A2(n_577),
.B(n_614),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_740),
.A2(n_577),
.B(n_614),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_679),
.B(n_649),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_703),
.B(n_556),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_792),
.A2(n_614),
.B(n_572),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_762),
.A2(n_574),
.B(n_572),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_762),
.A2(n_574),
.B(n_572),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_679),
.B(n_660),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_795),
.Y(n_862)
);

AND3x4_ASAP7_75t_L g863 ( 
.A(n_689),
.B(n_656),
.C(n_667),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_749),
.A2(n_671),
.B(n_613),
.C(n_661),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_778),
.A2(n_649),
.B1(n_672),
.B2(n_605),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_723),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_826),
.A2(n_594),
.B(n_604),
.Y(n_867)
);

CKINVDCx10_ASAP7_75t_R g868 ( 
.A(n_680),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_728),
.A2(n_594),
.B(n_604),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_766),
.B(n_590),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_691),
.B(n_649),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_749),
.B(n_556),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_753),
.B(n_649),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_708),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_731),
.A2(n_594),
.B(n_604),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_753),
.B(n_649),
.Y(n_876)
);

BUFx4f_ASAP7_75t_L g877 ( 
.A(n_827),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_674),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_747),
.B(n_603),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_720),
.A2(n_787),
.B1(n_743),
.B2(n_710),
.Y(n_880)
);

CKINVDCx10_ASAP7_75t_R g881 ( 
.A(n_804),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_708),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_757),
.A2(n_574),
.B(n_605),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_787),
.A2(n_585),
.B(n_589),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_692),
.A2(n_589),
.B(n_587),
.C(n_528),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_754),
.B(n_630),
.Y(n_886)
);

OAI321xp33_ASAP7_75t_L g887 ( 
.A1(n_702),
.A2(n_653),
.A3(n_652),
.B1(n_640),
.B2(n_620),
.C(n_564),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_676),
.Y(n_888)
);

OR2x6_ASAP7_75t_L g889 ( 
.A(n_685),
.B(n_630),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_693),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_707),
.B(n_630),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_754),
.B(n_603),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_695),
.A2(n_564),
.B(n_561),
.C(n_548),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_769),
.A2(n_558),
.B(n_563),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_722),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_697),
.Y(n_896)
);

CKINVDCx16_ASAP7_75t_R g897 ( 
.A(n_706),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_708),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_711),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_766),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_755),
.B(n_587),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_741),
.A2(n_653),
.B(n_652),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_710),
.A2(n_528),
.B1(n_553),
.B2(n_582),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_777),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_677),
.A2(n_563),
.B(n_612),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_755),
.B(n_528),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_739),
.A2(n_836),
.B(n_774),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_774),
.A2(n_563),
.B(n_612),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_758),
.A2(n_640),
.B(n_553),
.C(n_582),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_700),
.A2(n_538),
.B(n_531),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_774),
.A2(n_612),
.B(n_607),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_774),
.A2(n_612),
.B(n_607),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_777),
.B(n_582),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_710),
.A2(n_694),
.B1(n_803),
.B2(n_737),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_782),
.A2(n_540),
.B(n_607),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_758),
.A2(n_553),
.B(n_538),
.C(n_548),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_682),
.B(n_11),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_761),
.A2(n_573),
.B(n_561),
.C(n_531),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_712),
.A2(n_573),
.B(n_672),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_802),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_761),
.A2(n_767),
.B(n_796),
.C(n_801),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_711),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_716),
.A2(n_588),
.B(n_557),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_782),
.A2(n_588),
.B(n_557),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_782),
.A2(n_588),
.B(n_557),
.Y(n_926)
);

AOI221x1_ASAP7_75t_L g927 ( 
.A1(n_783),
.A2(n_717),
.B1(n_699),
.B2(n_696),
.C(n_789),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_782),
.A2(n_588),
.B(n_557),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_816),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_733),
.A2(n_607),
.B(n_540),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_722),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_834),
.A2(n_672),
.B(n_562),
.C(n_16),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_675),
.A2(n_562),
.B(n_650),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_711),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_812),
.B(n_12),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_737),
.B(n_672),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_736),
.A2(n_688),
.B(n_822),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_799),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_724),
.Y(n_939)
);

BUFx2_ASAP7_75t_SL g940 ( 
.A(n_705),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_742),
.A2(n_672),
.B(n_562),
.C(n_19),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_828),
.A2(n_540),
.B(n_650),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_709),
.B(n_650),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_735),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_711),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_807),
.B(n_15),
.Y(n_946)
);

AOI21x1_ASAP7_75t_L g947 ( 
.A1(n_831),
.A2(n_650),
.B(n_639),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_713),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_800),
.B(n_540),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_833),
.A2(n_639),
.B(n_136),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_833),
.A2(n_128),
.B1(n_127),
.B2(n_120),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_715),
.B(n_15),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_811),
.B(n_118),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_767),
.B(n_102),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_730),
.B(n_17),
.C(n_19),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_694),
.A2(n_90),
.B1(n_84),
.B2(n_82),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_806),
.A2(n_78),
.B(n_72),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_725),
.B(n_727),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_765),
.A2(n_66),
.B(n_63),
.Y(n_959)
);

NOR2x1p5_ASAP7_75t_SL g960 ( 
.A(n_686),
.B(n_25),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_824),
.A2(n_791),
.B(n_783),
.C(n_763),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_729),
.A2(n_25),
.B(n_26),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_746),
.A2(n_26),
.B(n_30),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_718),
.B(n_31),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_714),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_817),
.A2(n_34),
.B(n_35),
.Y(n_966)
);

NOR3xp33_ASAP7_75t_L g967 ( 
.A(n_704),
.B(n_35),
.C(n_36),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_742),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_764),
.B(n_37),
.Y(n_969)
);

NAND2x1p5_ASAP7_75t_L g970 ( 
.A(n_714),
.B(n_38),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_752),
.B(n_40),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_721),
.A2(n_41),
.B(n_43),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_824),
.B(n_45),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_745),
.A2(n_46),
.B(n_50),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_773),
.A2(n_46),
.B(n_51),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_751),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_830),
.A2(n_53),
.B(n_57),
.C(n_58),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_803),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_714),
.B(n_781),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_830),
.A2(n_841),
.B(n_760),
.C(n_745),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_832),
.A2(n_840),
.B(n_797),
.C(n_779),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_714),
.B(n_781),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_738),
.A2(n_744),
.B(n_786),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_748),
.A2(n_784),
.B(n_814),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_832),
.A2(n_785),
.B(n_841),
.C(n_821),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_794),
.A2(n_810),
.B(n_808),
.C(n_809),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_829),
.A2(n_719),
.B(n_732),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_798),
.A2(n_839),
.B(n_771),
.C(n_770),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_746),
.A2(n_768),
.B(n_835),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_756),
.B(n_687),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_781),
.A2(n_681),
.B(n_684),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_756),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_813),
.B(n_823),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_815),
.A2(n_776),
.B(n_793),
.C(n_825),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_776),
.B(n_818),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_724),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_818),
.A2(n_689),
.B(n_820),
.C(n_775),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_837),
.A2(n_788),
.B(n_805),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_724),
.A2(n_775),
.B(n_780),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_775),
.B(n_750),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_701),
.A2(n_577),
.B(n_569),
.Y(n_1001)
);

AO21x1_ASAP7_75t_L g1002 ( 
.A1(n_750),
.A2(n_698),
.B(n_691),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_701),
.A2(n_577),
.B(n_569),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_698),
.B(n_750),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_708),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_698),
.A2(n_750),
.B(n_753),
.C(n_749),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_701),
.A2(n_577),
.B(n_569),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_701),
.A2(n_577),
.B(n_569),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_698),
.B(n_750),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_708),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_675),
.A2(n_683),
.B(n_688),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_698),
.A2(n_720),
.B1(n_750),
.B2(n_787),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_750),
.B(n_698),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_819),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_838),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_698),
.A2(n_750),
.B1(n_720),
.B2(n_679),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_750),
.B(n_698),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_750),
.B(n_698),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_678),
.B(n_450),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_683),
.A2(n_701),
.B(n_759),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_678),
.B(n_450),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_698),
.A2(n_750),
.B1(n_720),
.B2(n_679),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_819),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_866),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_861),
.B(n_1006),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_1002),
.A2(n_909),
.A3(n_880),
.B(n_1012),
.Y(n_1033)
);

O2A1O1Ixp5_ASAP7_75t_L g1034 ( 
.A1(n_921),
.A2(n_973),
.B(n_985),
.C(n_993),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_843),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_1019),
.A2(n_1027),
.B(n_1013),
.Y(n_1036)
);

AND3x4_ASAP7_75t_L g1037 ( 
.A(n_967),
.B(n_863),
.C(n_897),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_868),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_916),
.A2(n_927),
.A3(n_849),
.B(n_844),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_900),
.Y(n_1040)
);

AO31x2_ASAP7_75t_L g1041 ( 
.A1(n_918),
.A2(n_876),
.A3(n_873),
.B(n_961),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_847),
.B(n_1017),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_902),
.A2(n_937),
.B(n_894),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_872),
.A2(n_856),
.B(n_848),
.C(n_886),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1018),
.A2(n_1024),
.B(n_1023),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_883),
.A2(n_984),
.B(n_947),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_965),
.B(n_874),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1018),
.A2(n_1024),
.B(n_1023),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_859),
.A2(n_860),
.B(n_869),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1025),
.B(n_995),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1025),
.B(n_892),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_904),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_901),
.B(n_906),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_875),
.A2(n_910),
.B(n_1001),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_1003),
.A2(n_1008),
.B(n_1007),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_989),
.A2(n_851),
.B(n_871),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_924),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_885),
.A2(n_907),
.B(n_893),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_994),
.A2(n_935),
.B(n_846),
.C(n_988),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_843),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_981),
.A2(n_936),
.B(n_919),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_972),
.A2(n_914),
.B1(n_966),
.B2(n_964),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_878),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_958),
.B(n_888),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_890),
.B(n_896),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_864),
.A2(n_848),
.A3(n_850),
.B(n_917),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_852),
.B(n_891),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_971),
.B(n_990),
.C(n_997),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_854),
.A2(n_991),
.B(n_986),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_853),
.A2(n_1028),
.B(n_1015),
.Y(n_1072)
);

INVx6_ASAP7_75t_L g1073 ( 
.A(n_843),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_948),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_965),
.B(n_874),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_854),
.A2(n_855),
.B(n_983),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_946),
.B(n_938),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_855),
.A2(n_950),
.B(n_850),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_SL g1079 ( 
.A1(n_950),
.A2(n_962),
.B(n_957),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_923),
.A2(n_867),
.B(n_942),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_952),
.A2(n_969),
.B(n_1000),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_923),
.A2(n_942),
.B(n_930),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_879),
.B(n_845),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_884),
.A2(n_998),
.B(n_887),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1016),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_858),
.A2(n_903),
.B(n_905),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_980),
.A2(n_865),
.B(n_932),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_879),
.B(n_929),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_922),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_862),
.B(n_944),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_992),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_928),
.B(n_926),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_954),
.A2(n_982),
.B(n_979),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_943),
.A2(n_949),
.B(n_974),
.Y(n_1094)
);

AOI221xp5_ASAP7_75t_L g1095 ( 
.A1(n_978),
.A2(n_977),
.B1(n_955),
.B2(n_968),
.C(n_975),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_920),
.B(n_913),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_925),
.A2(n_908),
.B(n_899),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_941),
.A2(n_975),
.B(n_951),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_956),
.A2(n_953),
.B(n_965),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_882),
.A2(n_899),
.B(n_898),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_882),
.B(n_898),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_911),
.A2(n_912),
.B(n_959),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_922),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_L g1104 ( 
.A(n_922),
.B(n_945),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_963),
.A2(n_970),
.B(n_996),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_965),
.B(n_1010),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_870),
.B(n_940),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_999),
.A2(n_960),
.B(n_976),
.C(n_996),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_889),
.A2(n_970),
.B1(n_934),
.B2(n_945),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_857),
.A2(n_1010),
.B(n_1005),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_889),
.B(n_934),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_889),
.A2(n_939),
.B(n_877),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_877),
.A2(n_881),
.B(n_895),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_931),
.B(n_853),
.Y(n_1114)
);

AOI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.Y(n_1115)
);

NOR2x1_ASAP7_75t_L g1116 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1022),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_878),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1121)
);

NAND2x1p5_ASAP7_75t_L g1122 ( 
.A(n_965),
.B(n_874),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_939),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1006),
.A2(n_1020),
.B(n_1014),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_842),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_L g1126 ( 
.A1(n_871),
.A2(n_848),
.B(n_989),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1002),
.A2(n_1006),
.A3(n_909),
.B(n_880),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_853),
.B(n_1015),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1130)
);

AO21x2_ASAP7_75t_L g1131 ( 
.A1(n_1006),
.A2(n_844),
.B(n_873),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.C(n_1006),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.C(n_1006),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_R g1134 ( 
.A(n_866),
.B(n_827),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_924),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_871),
.A2(n_848),
.B(n_989),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_900),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.C(n_1006),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1002),
.A2(n_1006),
.A3(n_909),
.B(n_880),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1022),
.B(n_533),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_871),
.A2(n_848),
.B(n_989),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.C(n_1006),
.Y(n_1150)
);

AO31x2_ASAP7_75t_L g1151 ( 
.A1(n_1002),
.A2(n_1006),
.A3(n_909),
.B(n_880),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_843),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_SL g1156 ( 
.A1(n_972),
.A2(n_950),
.B(n_966),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.C(n_1006),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1006),
.A2(n_1020),
.B(n_1014),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_849),
.A2(n_856),
.B(n_973),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1014),
.A2(n_1020),
.B1(n_1021),
.B2(n_1009),
.C(n_1004),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.C(n_1006),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_842),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_987),
.A2(n_933),
.B(n_1011),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_940),
.B(n_590),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1168)
);

AO21x1_ASAP7_75t_L g1169 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_878),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_878),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_900),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_847),
.A2(n_1017),
.B(n_1013),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1020),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_843),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1145),
.B(n_1066),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_1038),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_1123),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1129),
.B(n_1111),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1030),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1032),
.A2(n_1177),
.B1(n_1161),
.B2(n_1152),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1064),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1040),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1074),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1120),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1035),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1031),
.A2(n_1119),
.B(n_1118),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1052),
.A2(n_1043),
.B(n_1130),
.Y(n_1191)
);

INVx3_ASAP7_75t_SL g1192 ( 
.A(n_1114),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1173),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_1161),
.B(n_1133),
.C(n_1132),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1035),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1129),
.B(n_1112),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1138),
.A2(n_1176),
.B1(n_1152),
.B2(n_1170),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1138),
.A2(n_1176),
.B1(n_1170),
.B2(n_1146),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1121),
.A2(n_1135),
.B(n_1127),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1053),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1115),
.A2(n_1143),
.B(n_1158),
.C(n_1162),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1171),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1035),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1142),
.Y(n_1204)
);

NOR2x1_ASAP7_75t_L g1205 ( 
.A(n_1070),
.B(n_1167),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1115),
.A2(n_1150),
.B(n_1060),
.C(n_1063),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1077),
.B(n_1116),
.Y(n_1207)
);

OAI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_1124),
.A2(n_1159),
.B1(n_1029),
.B2(n_1063),
.C(n_1095),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1061),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1124),
.A2(n_1159),
.B1(n_1037),
.B2(n_1169),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1117),
.A2(n_1081),
.B1(n_1069),
.B2(n_1107),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1167),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1065),
.B(n_1036),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1034),
.A2(n_1156),
.B(n_1098),
.C(n_1036),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1058),
.B(n_1136),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1065),
.B(n_1054),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1172),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1167),
.B(n_1067),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1114),
.B(n_1083),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1073),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1054),
.B(n_1051),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1137),
.A2(n_1046),
.B(n_1168),
.Y(n_1222)
);

INVx3_ASAP7_75t_SL g1223 ( 
.A(n_1091),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1049),
.A2(n_1175),
.B(n_1174),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1048),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1061),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1051),
.B(n_1096),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1091),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1141),
.A2(n_1168),
.B(n_1174),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1085),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1141),
.A2(n_1175),
.B(n_1148),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1048),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1125),
.B(n_1165),
.Y(n_1233)
);

BUFx10_ASAP7_75t_L g1234 ( 
.A(n_1073),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1098),
.A2(n_1087),
.B1(n_1095),
.B2(n_1084),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1061),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1148),
.A2(n_1084),
.B(n_1042),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1083),
.B(n_1088),
.Y(n_1238)
);

INVxp33_ASAP7_75t_L g1239 ( 
.A(n_1134),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1087),
.A2(n_1109),
.B1(n_1108),
.B2(n_1096),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1090),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_1073),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1088),
.B(n_1072),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1042),
.A2(n_1062),
.B(n_1078),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1090),
.B(n_1154),
.Y(n_1245)
);

AND2x2_ASAP7_75t_SL g1246 ( 
.A(n_1104),
.B(n_1178),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1100),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1089),
.B(n_1154),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1101),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1113),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1089),
.B(n_1109),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1103),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1062),
.A2(n_1079),
.B(n_1057),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1045),
.B(n_1178),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1033),
.B(n_1151),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1075),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1110),
.B(n_1103),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1103),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1110),
.B(n_1033),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1105),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1033),
.B(n_1131),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1106),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1099),
.B(n_1144),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1131),
.B(n_1128),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1106),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_SL g1268 ( 
.A(n_1122),
.B(n_1094),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_1122),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1160),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1144),
.B(n_1068),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1093),
.A2(n_1126),
.B1(n_1139),
.B2(n_1147),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1144),
.B(n_1068),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1093),
.A2(n_1076),
.B1(n_1044),
.B2(n_1055),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1056),
.A2(n_1071),
.B1(n_1082),
.B2(n_1080),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1092),
.B(n_1086),
.Y(n_1276)
);

BUFx2_ASAP7_75t_SL g1277 ( 
.A(n_1041),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_SL g1278 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1102),
.B(n_1039),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1047),
.A2(n_1059),
.B1(n_1050),
.B2(n_1153),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1039),
.B(n_1140),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1149),
.B(n_1155),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_1163),
.Y(n_1283)
);

NAND2x1p5_ASAP7_75t_L g1284 ( 
.A(n_1164),
.B(n_1166),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1030),
.B(n_866),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1177),
.B(n_1014),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1064),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_SL g1288 ( 
.A1(n_1063),
.A2(n_972),
.B(n_1159),
.C(n_1124),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1167),
.B(n_590),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1066),
.B(n_1146),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1161),
.B(n_1014),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1040),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1129),
.B(n_1111),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1142),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1129),
.B(n_1111),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1032),
.B(n_1020),
.C(n_1014),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1053),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1129),
.B(n_1111),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1123),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1138),
.A2(n_1020),
.B1(n_1021),
.B2(n_1014),
.Y(n_1300)
);

NOR2x1_ASAP7_75t_SL g1301 ( 
.A(n_1167),
.B(n_1110),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1032),
.B(n_1020),
.C(n_1014),
.Y(n_1302)
);

AND2x6_ASAP7_75t_L g1303 ( 
.A(n_1032),
.B(n_1019),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1064),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1040),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1052),
.A2(n_1043),
.B(n_921),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1040),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1052),
.A2(n_1043),
.B(n_921),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1031),
.A2(n_1119),
.B(n_1118),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1030),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1032),
.A2(n_1014),
.B(n_1021),
.C(n_1020),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1048),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1048),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1161),
.B(n_1014),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1040),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1161),
.B(n_1014),
.Y(n_1316)
);

OR2x2_ASAP7_75t_SL g1317 ( 
.A(n_1138),
.B(n_897),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1129),
.B(n_1111),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1161),
.B(n_1014),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1161),
.B(n_1014),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1040),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1064),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1190),
.A2(n_1309),
.B(n_1199),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1229),
.A2(n_1231),
.B(n_1222),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1203),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1303),
.A2(n_1302),
.B1(n_1296),
.B2(n_1208),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1184),
.B(n_1210),
.Y(n_1327)
);

BUFx8_ASAP7_75t_L g1328 ( 
.A(n_1181),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1303),
.A2(n_1296),
.B1(n_1208),
.B2(n_1286),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1203),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1271),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1266),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1304),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1300),
.A2(n_1303),
.B1(n_1320),
.B2(n_1291),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1303),
.A2(n_1194),
.B1(n_1320),
.B2(n_1319),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1299),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1255),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1263),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1262),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1300),
.A2(n_1319),
.B1(n_1316),
.B2(n_1291),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1194),
.A2(n_1314),
.B1(n_1316),
.B2(n_1235),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1322),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1216),
.B(n_1238),
.Y(n_1343)
);

BUFx8_ASAP7_75t_SL g1344 ( 
.A(n_1180),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1314),
.A2(n_1235),
.B1(n_1250),
.B2(n_1240),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1240),
.A2(n_1207),
.B1(n_1219),
.B2(n_1218),
.Y(n_1346)
);

BUFx2_ASAP7_75t_R g1347 ( 
.A(n_1183),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1244),
.A2(n_1237),
.B(n_1253),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1277),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1263),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1290),
.B(n_1204),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1294),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1260),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1216),
.B(n_1198),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1249),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1228),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1270),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_1228),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1272),
.A2(n_1284),
.B(n_1244),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1281),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1205),
.A2(n_1213),
.B1(n_1218),
.B2(n_1197),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1213),
.A2(n_1179),
.B1(n_1182),
.B2(n_1318),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1251),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1185),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1206),
.A2(n_1201),
.B(n_1214),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1265),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1187),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1196),
.A2(n_1211),
.B1(n_1293),
.B2(n_1318),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1265),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1188),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1252),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1203),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1220),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1310),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1191),
.A2(n_1308),
.B(n_1306),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1202),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1225),
.Y(n_1377)
);

BUFx12f_ASAP7_75t_L g1378 ( 
.A(n_1212),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1241),
.B(n_1245),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1182),
.A2(n_1298),
.B1(n_1295),
.B2(n_1293),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1294),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1217),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1295),
.A2(n_1298),
.B1(n_1243),
.B2(n_1196),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1258),
.Y(n_1384)
);

INVx4_ASAP7_75t_SL g1385 ( 
.A(n_1273),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1221),
.B(n_1227),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1287),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1261),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1254),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1227),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1193),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1221),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1305),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1234),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1200),
.A2(n_1273),
.B1(n_1321),
.B2(n_1307),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1315),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1268),
.A2(n_1289),
.B1(n_1246),
.B2(n_1186),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1292),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1269),
.Y(n_1399)
);

BUFx4f_ASAP7_75t_SL g1400 ( 
.A(n_1223),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1230),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1233),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1273),
.Y(n_1403)
);

NOR2x1_ASAP7_75t_R g1404 ( 
.A(n_1236),
.B(n_1259),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1215),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1279),
.B(n_1247),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1233),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1257),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1248),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1272),
.A2(n_1282),
.B(n_1283),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1248),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1192),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1289),
.A2(n_1297),
.B1(n_1239),
.B2(n_1268),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1256),
.Y(n_1414)
);

BUFx12f_ASAP7_75t_L g1415 ( 
.A(n_1234),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1189),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1317),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1195),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1284),
.A2(n_1283),
.B(n_1282),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1273),
.Y(n_1420)
);

CKINVDCx11_ASAP7_75t_R g1421 ( 
.A(n_1242),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1278),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1278),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1276),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1276),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1288),
.B(n_1313),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1232),
.B(n_1313),
.Y(n_1427)
);

AO21x1_ASAP7_75t_SL g1428 ( 
.A1(n_1274),
.A2(n_1280),
.B(n_1275),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1242),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1269),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1301),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1289),
.A2(n_1285),
.B1(n_1267),
.B2(n_1312),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1264),
.B(n_1195),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1264),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1209),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1226),
.A2(n_1014),
.B1(n_1021),
.B2(n_1020),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1311),
.A2(n_1020),
.B1(n_1021),
.B2(n_1014),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1228),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1229),
.A2(n_1231),
.B(n_1224),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1303),
.A2(n_1014),
.B1(n_1021),
.B2(n_1020),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1184),
.B(n_1210),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1251),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1358),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1384),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1381),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1353),
.B(n_1331),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1358),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1384),
.B(n_1353),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1344),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1325),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1359),
.B(n_1338),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1352),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1391),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1331),
.B(n_1363),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1351),
.B(n_1398),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1379),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1389),
.A2(n_1423),
.A3(n_1422),
.B(n_1339),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1434),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1379),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1337),
.B(n_1332),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1434),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1359),
.A2(n_1323),
.B(n_1410),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1337),
.Y(n_1463)
);

AO21x1_ASAP7_75t_SL g1464 ( 
.A1(n_1431),
.A2(n_1326),
.B(n_1420),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1338),
.B(n_1350),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1343),
.B(n_1354),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1363),
.B(n_1442),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1442),
.B(n_1343),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1354),
.B(n_1335),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1388),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1365),
.A2(n_1324),
.B(n_1439),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1388),
.Y(n_1472)
);

AO21x2_ASAP7_75t_L g1473 ( 
.A1(n_1349),
.A2(n_1426),
.B(n_1419),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1428),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1406),
.A2(n_1375),
.B(n_1348),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1402),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1426),
.A2(n_1341),
.B(n_1329),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1405),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1403),
.A2(n_1420),
.B(n_1360),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1340),
.A2(n_1403),
.B(n_1437),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1355),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1327),
.B(n_1441),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1407),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1424),
.A2(n_1425),
.B(n_1441),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1405),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1416),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1361),
.A2(n_1424),
.B(n_1425),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1327),
.A2(n_1390),
.B(n_1392),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1370),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1386),
.B(n_1366),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_SL g1492 ( 
.A(n_1374),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1345),
.B(n_1369),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1387),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1387),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1433),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1369),
.B(n_1386),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1325),
.A2(n_1330),
.B(n_1372),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1390),
.B(n_1392),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1385),
.B(n_1377),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1364),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1367),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1376),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1382),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1418),
.Y(n_1505)
);

OAI21xp33_ASAP7_75t_L g1506 ( 
.A1(n_1436),
.A2(n_1346),
.B(n_1362),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1395),
.B(n_1417),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1457),
.B(n_1333),
.Y(n_1508)
);

NAND2xp33_ASAP7_75t_R g1509 ( 
.A(n_1449),
.B(n_1393),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1444),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1497),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1497),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1457),
.B(n_1342),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1448),
.B(n_1468),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1465),
.B(n_1385),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1457),
.B(n_1342),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1470),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1457),
.B(n_1408),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1470),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1472),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1448),
.B(n_1468),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1457),
.B(n_1413),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1497),
.B(n_1325),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1454),
.B(n_1428),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1466),
.B(n_1401),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_L g1527 ( 
.A(n_1443),
.B(n_1447),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1445),
.B(n_1368),
.Y(n_1528)
);

INVx5_ASAP7_75t_L g1529 ( 
.A(n_1474),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1506),
.A2(n_1397),
.B1(n_1373),
.B2(n_1383),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1497),
.Y(n_1531)
);

AOI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1488),
.A2(n_1432),
.B1(n_1411),
.B2(n_1409),
.C(n_1414),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1465),
.B(n_1385),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1472),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1444),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1461),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1489),
.B(n_1373),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1443),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1453),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1465),
.B(n_1433),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1467),
.B(n_1433),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1412),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1489),
.B(n_1435),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1497),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1467),
.B(n_1435),
.Y(n_1545)
);

NOR3xp33_ASAP7_75t_L g1546 ( 
.A(n_1506),
.B(n_1399),
.C(n_1404),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1465),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1463),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1465),
.B(n_1357),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1452),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1463),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1479),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1469),
.B(n_1427),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1501),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1492),
.B(n_1393),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1539),
.B(n_1458),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1530),
.A2(n_1522),
.B(n_1482),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1552),
.A2(n_1462),
.B(n_1475),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1522),
.A2(n_1507),
.B1(n_1482),
.B2(n_1485),
.C(n_1478),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1514),
.B(n_1491),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1546),
.A2(n_1474),
.B(n_1507),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1456),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1459),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1528),
.A2(n_1474),
.B(n_1493),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1510),
.B(n_1504),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1532),
.A2(n_1486),
.B1(n_1505),
.B2(n_1455),
.C(n_1502),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1511),
.B(n_1512),
.Y(n_1567)
);

AOI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1537),
.B2(n_1542),
.C(n_1526),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1504),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1501),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1537),
.B(n_1357),
.C(n_1477),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1503),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1529),
.B(n_1347),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1541),
.B(n_1480),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1545),
.B(n_1480),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1545),
.B(n_1480),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1508),
.B(n_1357),
.C(n_1477),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1544),
.B(n_1479),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1554),
.B(n_1517),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1508),
.B(n_1357),
.C(n_1477),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1519),
.B(n_1480),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1540),
.A2(n_1474),
.B1(n_1493),
.B2(n_1477),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1518),
.B(n_1476),
.C(n_1483),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1520),
.B(n_1490),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1534),
.B(n_1490),
.Y(n_1588)
);

NOR3xp33_ASAP7_75t_L g1589 ( 
.A(n_1555),
.B(n_1399),
.C(n_1450),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1551),
.B(n_1494),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1549),
.B(n_1474),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1548),
.B(n_1494),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1548),
.B(n_1495),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1549),
.B(n_1527),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1544),
.B(n_1484),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1529),
.A2(n_1471),
.B1(n_1500),
.B2(n_1487),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1549),
.A2(n_1464),
.B1(n_1378),
.B2(n_1496),
.Y(n_1597)
);

OAI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1543),
.A2(n_1380),
.B1(n_1430),
.B2(n_1356),
.C(n_1438),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1518),
.A2(n_1446),
.B1(n_1499),
.B2(n_1460),
.C(n_1451),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1524),
.B(n_1481),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1538),
.B(n_1396),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1582),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1592),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1593),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1557),
.A2(n_1471),
.B1(n_1464),
.B2(n_1515),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1571),
.B(n_1525),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1580),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1543),
.Y(n_1608)
);

AND2x2_ASAP7_75t_SL g1609 ( 
.A(n_1585),
.B(n_1547),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1580),
.B(n_1547),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1581),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1513),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1573),
.B(n_1515),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1558),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1595),
.Y(n_1615)
);

INVx3_ASAP7_75t_R g1616 ( 
.A(n_1575),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1577),
.B(n_1513),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1596),
.B(n_1523),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1565),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1578),
.B(n_1516),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1558),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1533),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1558),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1558),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1567),
.B(n_1576),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1587),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1588),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1586),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1557),
.A2(n_1533),
.B1(n_1378),
.B2(n_1487),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1603),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1600),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1612),
.B(n_1579),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1604),
.Y(n_1636)
);

OA211x2_ASAP7_75t_L g1637 ( 
.A1(n_1630),
.A2(n_1575),
.B(n_1601),
.C(n_1594),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1609),
.B(n_1559),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1627),
.B(n_1591),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1627),
.B(n_1560),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1628),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1612),
.B(n_1583),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1617),
.B(n_1583),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1623),
.B(n_1572),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1628),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1622),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1627),
.B(n_1562),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1628),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1617),
.B(n_1572),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1602),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1629),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1613),
.B(n_1563),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1608),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1621),
.B(n_1556),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1622),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1629),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1622),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1613),
.B(n_1574),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1629),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1632),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1630),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1632),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1620),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1613),
.B(n_1524),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1643),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1667),
.B(n_1608),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1615),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1646),
.B(n_1615),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1643),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1657),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1647),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1646),
.B(n_1623),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1615),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1650),
.Y(n_1684)
);

AOI21xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1656),
.A2(n_1609),
.B(n_1509),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1637),
.A2(n_1605),
.B1(n_1609),
.B2(n_1631),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1656),
.B(n_1620),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1650),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1654),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1642),
.B(n_1652),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1653),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1644),
.B(n_1606),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1670),
.B(n_1623),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1670),
.B(n_1623),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1642),
.B(n_1634),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1648),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1654),
.B(n_1623),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1648),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1659),
.B(n_1619),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1659),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1662),
.B(n_1564),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

OAI22xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1640),
.A2(n_1611),
.B1(n_1614),
.B2(n_1599),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1663),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1610),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1663),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1666),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1641),
.B(n_1655),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1644),
.A2(n_1609),
.B(n_1561),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1658),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1666),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1671),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1682),
.B(n_1668),
.Y(n_1716)
);

CKINVDCx16_ASAP7_75t_R g1717 ( 
.A(n_1687),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1692),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_SL g1719 ( 
.A1(n_1705),
.A2(n_1619),
.B1(n_1637),
.B2(n_1645),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1703),
.B(n_1374),
.Y(n_1720)
);

NOR2x1_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1651),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1711),
.A2(n_1619),
.B1(n_1631),
.B2(n_1605),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1685),
.B(n_1328),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1678),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1691),
.B(n_1661),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1712),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1671),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1682),
.A2(n_1589),
.B1(n_1651),
.B2(n_1598),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1673),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1697),
.B(n_1661),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1682),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1328),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1681),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1713),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1710),
.B(n_1655),
.Y(n_1735)
);

AND3x2_ASAP7_75t_L g1736 ( 
.A(n_1673),
.B(n_1664),
.C(n_1607),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1676),
.B(n_1669),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1677),
.B(n_1669),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1674),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1712),
.Y(n_1740)
);

CKINVDCx16_ASAP7_75t_R g1741 ( 
.A(n_1674),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1710),
.B(n_1668),
.Y(n_1742)
);

BUFx2_ASAP7_75t_SL g1743 ( 
.A(n_1683),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1681),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1684),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1684),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1712),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1706),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1696),
.B(n_1613),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1715),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1724),
.B(n_1680),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1720),
.B(n_1696),
.Y(n_1753)
);

NAND4xp25_ASAP7_75t_L g1754 ( 
.A(n_1719),
.B(n_1683),
.C(n_1566),
.D(n_1701),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1734),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1715),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1717),
.B(n_1693),
.C(n_1706),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1718),
.B(n_1686),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1727),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1717),
.B(n_1701),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1721),
.A2(n_1701),
.B(n_1561),
.Y(n_1761)
);

NAND4xp75_ASAP7_75t_L g1762 ( 
.A(n_1723),
.B(n_1732),
.C(n_1733),
.D(n_1727),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1722),
.A2(n_1679),
.B(n_1675),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1731),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1733),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1736),
.A2(n_1564),
.B(n_1694),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1741),
.B(n_1695),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1729),
.A2(n_1694),
.B1(n_1695),
.B2(n_1699),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1693),
.C(n_1690),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1739),
.B(n_1707),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1735),
.B(n_1699),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1731),
.A2(n_1725),
.B(n_1735),
.Y(n_1772)
);

AOI31xp33_ASAP7_75t_L g1773 ( 
.A1(n_1714),
.A2(n_1396),
.A3(n_1328),
.B(n_1336),
.Y(n_1773)
);

OAI32xp33_ASAP7_75t_L g1774 ( 
.A1(n_1742),
.A2(n_1614),
.A3(n_1625),
.B1(n_1624),
.B2(n_1702),
.Y(n_1774)
);

OAI21xp33_ASAP7_75t_L g1775 ( 
.A1(n_1730),
.A2(n_1699),
.B(n_1694),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1755),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1767),
.B(n_1743),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1755),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1757),
.A2(n_1743),
.B1(n_1716),
.B2(n_1749),
.Y(n_1779)
);

INVxp33_ASAP7_75t_L g1780 ( 
.A(n_1760),
.Y(n_1780)
);

NAND2x1_ASAP7_75t_L g1781 ( 
.A(n_1767),
.B(n_1716),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1764),
.B(n_1716),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1750),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1764),
.B(n_1772),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1750),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1753),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.B(n_1749),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1752),
.B(n_1737),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1758),
.B(n_1737),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1761),
.B(n_1616),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1754),
.B(n_1738),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1751),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1762),
.B(n_1738),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1763),
.B(n_1744),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1773),
.B(n_1744),
.Y(n_1795)
);

XOR2x2_ASAP7_75t_L g1796 ( 
.A(n_1793),
.B(n_1769),
.Y(n_1796)
);

AOI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1791),
.A2(n_1766),
.B(n_1775),
.C(n_1774),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1779),
.A2(n_1768),
.B(n_1756),
.C(n_1759),
.Y(n_1798)
);

AOI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1780),
.A2(n_1770),
.B(n_1765),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1781),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1780),
.B(n_1771),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1794),
.A2(n_1746),
.B(n_1745),
.Y(n_1802)
);

NOR4xp25_ASAP7_75t_L g1803 ( 
.A(n_1784),
.B(n_1748),
.C(n_1745),
.D(n_1746),
.Y(n_1803)
);

AOI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1790),
.A2(n_1748),
.B(n_1747),
.C(n_1726),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1777),
.A2(n_1740),
.B(n_1726),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1790),
.A2(n_1747),
.B(n_1740),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1776),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1786),
.A2(n_1689),
.B1(n_1709),
.B2(n_1708),
.C(n_1704),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1807),
.Y(n_1809)
);

NAND4xp75_ASAP7_75t_L g1810 ( 
.A(n_1800),
.B(n_1778),
.C(n_1777),
.D(n_1795),
.Y(n_1810)
);

AND4x1_ASAP7_75t_L g1811 ( 
.A(n_1801),
.B(n_1782),
.C(n_1789),
.D(n_1792),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1799),
.B(n_1783),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1798),
.B(n_1785),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1805),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1806),
.B(n_1788),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1796),
.A2(n_1788),
.B(n_1787),
.Y(n_1816)
);

AOI211x1_ASAP7_75t_SL g1817 ( 
.A1(n_1802),
.A2(n_1698),
.B(n_1700),
.C(n_1648),
.Y(n_1817)
);

NOR2x1_ASAP7_75t_L g1818 ( 
.A(n_1803),
.B(n_1787),
.Y(n_1818)
);

NOR3xp33_ASAP7_75t_L g1819 ( 
.A(n_1797),
.B(n_1429),
.C(n_1421),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1818),
.A2(n_1808),
.B(n_1804),
.Y(n_1820)
);

NOR3x2_ASAP7_75t_L g1821 ( 
.A(n_1810),
.B(n_1336),
.C(n_1400),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1813),
.A2(n_1713),
.B(n_1700),
.Y(n_1822)
);

OAI211xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1819),
.A2(n_1336),
.B(n_1438),
.C(n_1356),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1815),
.B(n_1698),
.Y(n_1824)
);

CKINVDCx16_ASAP7_75t_R g1825 ( 
.A(n_1821),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1824),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1820),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_SL g1828 ( 
.A(n_1822),
.B(n_1816),
.C(n_1811),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1823),
.B(n_1812),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1824),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1825),
.B(n_1814),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1829),
.B(n_1809),
.Y(n_1832)
);

NOR2x1p5_ASAP7_75t_L g1833 ( 
.A(n_1828),
.B(n_1371),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1827),
.B(n_1817),
.Y(n_1834)
);

NAND4xp25_ASAP7_75t_L g1835 ( 
.A(n_1828),
.B(n_1371),
.C(n_1597),
.D(n_1415),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1831),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1832),
.Y(n_1837)
);

AOI22x1_ASAP7_75t_L g1838 ( 
.A1(n_1833),
.A2(n_1830),
.B1(n_1826),
.B2(n_1415),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1836),
.B(n_1835),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_SL g1840 ( 
.A1(n_1839),
.A2(n_1837),
.B1(n_1834),
.B2(n_1838),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1840),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1840),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1842),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1841),
.B(n_1394),
.C(n_1665),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1843),
.A2(n_1394),
.B(n_1665),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1844),
.B(n_1613),
.Y(n_1846)
);

OA22x2_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1665),
.B1(n_1660),
.B2(n_1658),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1847),
.A2(n_1845),
.B1(n_1660),
.B2(n_1538),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1848),
.A2(n_1639),
.B1(n_1638),
.B2(n_1636),
.C(n_1633),
.Y(n_1849)
);

AOI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1430),
.B(n_1498),
.C(n_1330),
.Y(n_1850)
);


endmodule