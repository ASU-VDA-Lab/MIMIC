module real_aes_10368_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1931;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1916;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AO221x1_ASAP7_75t_L g1608 ( .A1(n_0), .A2(n_151), .B1(n_1560), .B2(n_1609), .C(n_1611), .Y(n_1608) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_1), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_1), .A2(n_11), .B1(n_691), .B2(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_2), .A2(n_94), .B1(n_793), .B2(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1450 ( .A(n_2), .Y(n_1450) );
INVx1_ASAP7_75t_L g944 ( .A(n_3), .Y(n_944) );
INVx1_ASAP7_75t_L g1180 ( .A(n_4), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1585 ( .A1(n_5), .A2(n_134), .B1(n_1560), .B2(n_1566), .Y(n_1585) );
INVx1_ASAP7_75t_L g1319 ( .A(n_6), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_7), .A2(n_251), .B1(n_535), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_7), .A2(n_251), .B1(n_631), .B2(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_8), .A2(n_188), .B1(n_570), .B2(n_631), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_8), .A2(n_188), .B1(n_640), .B2(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g655 ( .A(n_9), .Y(n_655) );
INVx1_ASAP7_75t_L g1422 ( .A(n_10), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_10), .A2(n_279), .B1(n_691), .B2(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g664 ( .A(n_11), .Y(n_664) );
INVxp33_ASAP7_75t_SL g1281 ( .A(n_12), .Y(n_1281) );
AOI22xp5_ASAP7_75t_SL g1306 ( .A1(n_12), .A2(n_309), .B1(n_703), .B2(n_963), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g1365 ( .A(n_13), .Y(n_1365) );
INVx1_ASAP7_75t_L g1893 ( .A(n_14), .Y(n_1893) );
AO22x1_ASAP7_75t_L g1263 ( .A1(n_15), .A2(n_1264), .B1(n_1265), .B2(n_1310), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_15), .Y(n_1264) );
AOI22xp33_ASAP7_75t_SL g1289 ( .A1(n_16), .A2(n_249), .B1(n_537), .B2(n_1290), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_16), .A2(n_249), .B1(n_1303), .B2(n_1305), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1930 ( .A1(n_17), .A2(n_241), .B1(n_601), .B2(n_1931), .Y(n_1930) );
AOI22xp33_ASAP7_75t_L g1936 ( .A1(n_17), .A2(n_241), .B1(n_920), .B2(n_1937), .Y(n_1936) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_18), .A2(n_269), .B1(n_523), .B2(n_745), .Y(n_1086) );
AOI221xp5_ASAP7_75t_SL g1095 ( .A1(n_18), .A2(n_558), .B1(n_1096), .B2(n_1097), .C(n_1105), .Y(n_1095) );
INVx1_ASAP7_75t_L g654 ( .A(n_19), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_19), .A2(n_69), .B1(n_636), .B2(n_684), .Y(n_694) );
INVx1_ASAP7_75t_L g1612 ( .A(n_20), .Y(n_1612) );
INVx1_ASAP7_75t_L g1925 ( .A(n_21), .Y(n_1925) );
OAI22xp5_ASAP7_75t_L g1944 ( .A1(n_21), .A2(n_263), .B1(n_670), .B2(n_1005), .Y(n_1944) );
INVx1_ASAP7_75t_L g782 ( .A(n_22), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_22), .A2(n_340), .B1(n_581), .B2(n_586), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1441 ( .A1(n_23), .A2(n_367), .B1(n_590), .B2(n_751), .Y(n_1441) );
INVx1_ASAP7_75t_L g1447 ( .A(n_23), .Y(n_1447) );
INVx1_ASAP7_75t_L g832 ( .A(n_24), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_25), .A2(n_83), .B1(n_511), .B2(n_514), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_25), .A2(n_83), .B1(n_552), .B2(n_555), .Y(n_551) );
INVxp67_ASAP7_75t_SL g1332 ( .A(n_26), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_26), .A2(n_238), .B1(n_963), .B2(n_1258), .Y(n_1354) );
INVx1_ASAP7_75t_L g436 ( .A(n_27), .Y(n_436) );
INVx1_ASAP7_75t_L g740 ( .A(n_28), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_28), .A2(n_220), .B1(n_570), .B2(n_571), .Y(n_756) );
CKINVDCx5p33_ASAP7_75t_R g1403 ( .A(n_29), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_30), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g1525 ( .A1(n_31), .A2(n_99), .B1(n_601), .B2(n_1526), .Y(n_1525) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_31), .A2(n_99), .B1(n_1258), .B2(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g826 ( .A(n_32), .Y(n_826) );
INVx1_ASAP7_75t_L g1156 ( .A(n_33), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_33), .A2(n_242), .B1(n_581), .B2(n_596), .Y(n_1160) );
CKINVDCx5p33_ASAP7_75t_R g1404 ( .A(n_34), .Y(n_1404) );
INVx1_ASAP7_75t_L g1373 ( .A(n_35), .Y(n_1373) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_35), .A2(n_204), .B1(n_640), .B2(n_644), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_36), .A2(n_150), .B1(n_963), .B2(n_1129), .Y(n_1128) );
INVxp67_ASAP7_75t_SL g1141 ( .A(n_36), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1940 ( .A1(n_37), .A2(n_363), .B1(n_1195), .B2(n_1203), .Y(n_1940) );
INVxp67_ASAP7_75t_SL g1947 ( .A(n_37), .Y(n_1947) );
OAI211xp5_ASAP7_75t_L g1059 ( .A1(n_38), .A2(n_449), .B(n_1060), .C(n_1062), .Y(n_1059) );
INVx1_ASAP7_75t_L g1090 ( .A(n_38), .Y(n_1090) );
INVx1_ASAP7_75t_L g382 ( .A(n_39), .Y(n_382) );
XNOR2xp5_ASAP7_75t_L g1359 ( .A(n_40), .B(n_1360), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_41), .A2(n_253), .B1(n_601), .B2(n_602), .C(n_603), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_41), .A2(n_253), .B1(n_570), .B2(n_571), .Y(n_626) );
OAI211xp5_ASAP7_75t_L g1116 ( .A1(n_42), .A2(n_449), .B(n_1117), .C(n_1118), .Y(n_1116) );
INVx1_ASAP7_75t_L g1134 ( .A(n_42), .Y(n_1134) );
XNOR2xp5_ASAP7_75t_L g1172 ( .A(n_43), .B(n_1173), .Y(n_1172) );
INVxp67_ASAP7_75t_L g1238 ( .A(n_44), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_44), .A2(n_299), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
INVx1_ASAP7_75t_L g1275 ( .A(n_45), .Y(n_1275) );
AOI22xp5_ASAP7_75t_L g1581 ( .A1(n_46), .A2(n_162), .B1(n_1560), .B2(n_1566), .Y(n_1581) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_47), .A2(n_131), .B1(n_581), .B2(n_596), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_47), .A2(n_131), .B1(n_520), .B2(n_1025), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1229 ( .A(n_48), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_48), .A2(n_375), .B1(n_670), .B2(n_671), .Y(n_1235) );
AOI22xp33_ASAP7_75t_SL g1929 ( .A1(n_49), .A2(n_208), .B1(n_519), .B2(n_1294), .Y(n_1929) );
AOI22xp33_ASAP7_75t_SL g1938 ( .A1(n_49), .A2(n_208), .B1(n_1193), .B2(n_1200), .Y(n_1938) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_50), .A2(n_356), .B1(n_1018), .B2(n_1020), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_50), .A2(n_254), .B1(n_1037), .B2(n_1039), .Y(n_1036) );
INVxp33_ASAP7_75t_L g1522 ( .A(n_51), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1544 ( .A1(n_51), .A2(n_312), .B1(n_710), .B2(n_860), .Y(n_1544) );
INVxp33_ASAP7_75t_SL g1286 ( .A(n_52), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_52), .A2(n_307), .B1(n_1303), .B2(n_1308), .Y(n_1307) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_53), .A2(n_351), .B1(n_581), .B2(n_596), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_53), .A2(n_266), .B1(n_532), .B2(n_897), .Y(n_1189) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_54), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_55), .A2(n_214), .B1(n_636), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_55), .A2(n_214), .B1(n_590), .B2(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g1846 ( .A(n_56), .Y(n_1846) );
INVxp33_ASAP7_75t_SL g1320 ( .A(n_57), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_57), .A2(n_218), .B1(n_691), .B2(n_1028), .Y(n_1337) );
INVxp33_ASAP7_75t_SL g1334 ( .A(n_58), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_58), .A2(n_79), .B1(n_487), .B2(n_1350), .Y(n_1353) );
AO221x2_ASAP7_75t_L g1707 ( .A1(n_59), .A2(n_289), .B1(n_1609), .B2(n_1708), .C(n_1710), .Y(n_1707) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_60), .A2(n_64), .B1(n_1030), .B2(n_1244), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_60), .A2(n_64), .B1(n_1041), .B2(n_1252), .Y(n_1251) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_61), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_61), .A2(n_77), .B1(n_568), .B2(n_571), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_62), .A2(n_121), .B1(n_640), .B2(n_644), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_62), .A2(n_110), .B1(n_926), .B2(n_927), .Y(n_925) );
INVxp33_ASAP7_75t_SL g1008 ( .A(n_63), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_63), .A2(n_182), .B1(n_1039), .B2(n_1043), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_65), .A2(n_370), .B1(n_640), .B2(n_644), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_65), .A2(n_370), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
INVxp67_ASAP7_75t_SL g1467 ( .A(n_66), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_66), .A2(n_237), .B1(n_532), .B2(n_602), .Y(n_1479) );
OAI22xp33_ASAP7_75t_L g1063 ( .A1(n_67), .A2(n_156), .B1(n_391), .B2(n_410), .Y(n_1063) );
INVx1_ASAP7_75t_L g1089 ( .A(n_67), .Y(n_1089) );
INVx1_ASAP7_75t_L g628 ( .A(n_68), .Y(n_628) );
INVx1_ASAP7_75t_L g657 ( .A(n_69), .Y(n_657) );
INVx1_ASAP7_75t_L g668 ( .A(n_70), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_70), .A2(n_273), .B1(n_575), .B2(n_710), .Y(n_709) );
OAI211xp5_ASAP7_75t_L g587 ( .A1(n_71), .A2(n_588), .B(n_591), .C(n_592), .Y(n_587) );
INVx1_ASAP7_75t_L g616 ( .A(n_71), .Y(n_616) );
XNOR2xp5_ASAP7_75t_L g1414 ( .A(n_72), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g947 ( .A(n_73), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_74), .A2(n_1047), .B1(n_1107), .B2(n_1108), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_74), .Y(n_1108) );
INVx1_ASAP7_75t_L g939 ( .A(n_75), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_75), .A2(n_178), .B1(n_486), .B2(n_963), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_76), .A2(n_322), .B1(n_1560), .B2(n_1566), .Y(n_1559) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_77), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g1584 ( .A1(n_78), .A2(n_347), .B1(n_1568), .B2(n_1574), .Y(n_1584) );
INVxp67_ASAP7_75t_SL g1328 ( .A(n_79), .Y(n_1328) );
INVxp33_ASAP7_75t_SL g1813 ( .A(n_80), .Y(n_1813) );
AOI22xp33_ASAP7_75t_L g1863 ( .A1(n_80), .A2(n_364), .B1(n_552), .B2(n_1136), .Y(n_1863) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_81), .A2(n_160), .B1(n_897), .B2(n_1242), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_81), .A2(n_160), .B1(n_825), .B2(n_920), .Y(n_1254) );
INVx1_ASAP7_75t_L g823 ( .A(n_82), .Y(n_823) );
AO22x2_ASAP7_75t_L g871 ( .A1(n_84), .A2(n_872), .B1(n_873), .B2(n_929), .Y(n_871) );
INVxp67_ASAP7_75t_L g929 ( .A(n_84), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_85), .Y(n_808) );
AO22x1_ASAP7_75t_L g1600 ( .A1(n_86), .A2(n_272), .B1(n_1566), .B2(n_1601), .Y(n_1600) );
INVxp33_ASAP7_75t_SL g955 ( .A(n_87), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_87), .A2(n_169), .B1(n_511), .B2(n_905), .Y(n_979) );
XOR2xp5_ASAP7_75t_L g988 ( .A(n_88), .B(n_989), .Y(n_988) );
AO22x1_ASAP7_75t_L g1602 ( .A1(n_88), .A2(n_270), .B1(n_1568), .B2(n_1574), .Y(n_1602) );
INVx1_ASAP7_75t_L g995 ( .A(n_89), .Y(n_995) );
OAI222xp33_ASAP7_75t_L g1004 ( .A1(n_89), .A2(n_195), .B1(n_291), .B2(n_438), .C1(n_607), .C2(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1274 ( .A(n_90), .Y(n_1274) );
AOI22xp33_ASAP7_75t_SL g1293 ( .A1(n_90), .A2(n_129), .B1(n_1290), .B2(n_1294), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_91), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_91), .A2(n_106), .B1(n_1100), .B2(n_1103), .Y(n_1099) );
INVx1_ASAP7_75t_L g1126 ( .A(n_92), .Y(n_1126) );
OAI21xp33_ASAP7_75t_SL g993 ( .A1(n_93), .A2(n_789), .B(n_994), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_93), .A2(n_326), .B1(n_1028), .B2(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g1451 ( .A(n_94), .Y(n_1451) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_95), .A2(n_105), .B1(n_1345), .B2(n_1347), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_95), .A2(n_105), .B1(n_487), .B2(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1271 ( .A(n_96), .Y(n_1271) );
INVxp67_ASAP7_75t_SL g1838 ( .A(n_97), .Y(n_1838) );
AOI221xp5_ASAP7_75t_L g1880 ( .A1(n_97), .A2(n_368), .B1(n_1881), .B2(n_1882), .C(n_1883), .Y(n_1880) );
CKINVDCx5p33_ASAP7_75t_R g1418 ( .A(n_98), .Y(n_1418) );
BUFx2_ASAP7_75t_L g454 ( .A(n_100), .Y(n_454) );
BUFx2_ASAP7_75t_L g507 ( .A(n_100), .Y(n_507) );
INVx1_ASAP7_75t_L g542 ( .A(n_100), .Y(n_542) );
OR2x2_ASAP7_75t_L g1822 ( .A(n_100), .B(n_1823), .Y(n_1822) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_101), .A2(n_204), .B1(n_700), .B2(n_1375), .Y(n_1374) );
OAI211xp5_ASAP7_75t_L g1401 ( .A1(n_101), .A2(n_449), .B(n_913), .C(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1923 ( .A(n_102), .Y(n_1923) );
AOI22xp33_ASAP7_75t_SL g1934 ( .A1(n_102), .A2(n_213), .B1(n_519), .B2(n_1481), .Y(n_1934) );
AOI22xp33_ASAP7_75t_SL g1186 ( .A1(n_103), .A2(n_258), .B1(n_519), .B2(n_731), .Y(n_1186) );
AOI22xp33_ASAP7_75t_SL g1192 ( .A1(n_103), .A2(n_258), .B1(n_1041), .B2(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1322 ( .A(n_104), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_104), .A2(n_126), .B1(n_523), .B2(n_684), .Y(n_1338) );
INVxp67_ASAP7_75t_SL g1085 ( .A(n_106), .Y(n_1085) );
INVx1_ASAP7_75t_L g722 ( .A(n_107), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_107), .A2(n_365), .B1(n_513), .B2(n_535), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_108), .A2(n_297), .B1(n_691), .B2(n_1341), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_108), .A2(n_297), .B1(n_1092), .B2(n_1301), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_109), .A2(n_330), .B1(n_519), .B2(n_523), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_109), .A2(n_330), .B1(n_547), .B2(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g882 ( .A(n_110), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g1815 ( .A1(n_111), .A2(n_200), .B1(n_1816), .B2(n_1824), .C(n_1828), .Y(n_1815) );
OAI22xp5_ASAP7_75t_L g1868 ( .A1(n_111), .A2(n_200), .B1(n_1869), .B2(n_1874), .Y(n_1868) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_112), .A2(n_268), .B1(n_596), .B2(n_597), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_112), .A2(n_268), .B1(n_511), .B2(n_533), .C(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_113), .A2(n_254), .B1(n_1012), .B2(n_1015), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_113), .A2(n_356), .B1(n_1033), .B2(n_1035), .Y(n_1032) );
INVx1_ASAP7_75t_L g1398 ( .A(n_114), .Y(n_1398) );
OAI211xp5_ASAP7_75t_SL g1409 ( .A1(n_114), .A2(n_497), .B(n_887), .C(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g861 ( .A(n_115), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_116), .A2(n_117), .B1(n_640), .B2(n_644), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_116), .A2(n_117), .B1(n_801), .B2(n_1136), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_118), .A2(n_128), .B1(n_662), .B2(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_118), .A2(n_128), .B1(n_671), .B2(n_735), .Y(n_734) );
AO221x1_ASAP7_75t_L g1595 ( .A1(n_119), .A2(n_138), .B1(n_1560), .B2(n_1566), .C(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1278 ( .A(n_120), .Y(n_1278) );
INVx1_ASAP7_75t_L g924 ( .A(n_121), .Y(n_924) );
AO221x1_ASAP7_75t_L g1587 ( .A1(n_122), .A2(n_334), .B1(n_1560), .B2(n_1566), .C(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1592 ( .A(n_123), .Y(n_1592) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_124), .A2(n_154), .B1(n_968), .B2(n_971), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_124), .A2(n_154), .B1(n_905), .B2(n_940), .Y(n_977) );
INVx1_ASAP7_75t_L g604 ( .A(n_125), .Y(n_604) );
INVxp33_ASAP7_75t_SL g1316 ( .A(n_126), .Y(n_1316) );
INVx1_ASAP7_75t_L g854 ( .A(n_127), .Y(n_854) );
INVxp33_ASAP7_75t_SL g1268 ( .A(n_129), .Y(n_1268) );
INVxp33_ASAP7_75t_SL g936 ( .A(n_130), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_130), .A2(n_181), .B1(n_962), .B2(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g836 ( .A(n_132), .Y(n_836) );
OAI22xp33_ASAP7_75t_SL g867 ( .A1(n_132), .A2(n_240), .B1(n_391), .B2(n_640), .Y(n_867) );
INVx1_ASAP7_75t_L g1598 ( .A(n_133), .Y(n_1598) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_135), .A2(n_248), .B1(n_1203), .B2(n_1205), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_135), .A2(n_248), .B1(n_640), .B2(n_644), .Y(n_1215) );
INVx1_ASAP7_75t_L g594 ( .A(n_136), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_137), .A2(n_168), .B1(n_1568), .B2(n_1574), .Y(n_1580) );
INVxp33_ASAP7_75t_SL g1519 ( .A(n_139), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_139), .A2(n_239), .B1(n_1546), .B2(n_1547), .Y(n_1545) );
AOI22xp33_ASAP7_75t_L g1486 ( .A1(n_140), .A2(n_275), .B1(n_547), .B2(n_1252), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g1491 ( .A(n_140), .Y(n_1491) );
INVxp67_ASAP7_75t_SL g1232 ( .A(n_141), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_141), .A2(n_321), .B1(n_710), .B2(n_1252), .Y(n_1256) );
XOR2xp5_ASAP7_75t_L g758 ( .A(n_142), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g1711 ( .A(n_143), .Y(n_1711) );
INVx1_ASAP7_75t_L g1421 ( .A(n_144), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_144), .A2(n_282), .B1(n_523), .B2(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1471 ( .A(n_145), .Y(n_1471) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_145), .A2(n_323), .B1(n_670), .B2(n_1005), .Y(n_1492) );
INVxp33_ASAP7_75t_L g457 ( .A(n_146), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_146), .A2(n_203), .B1(n_519), .B2(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_147), .A2(n_266), .B1(n_586), .B2(n_597), .Y(n_1176) );
INVxp33_ASAP7_75t_SL g1214 ( .A(n_147), .Y(n_1214) );
AOI22xp33_ASAP7_75t_SL g1527 ( .A1(n_148), .A2(n_319), .B1(n_1528), .B2(n_1530), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_148), .A2(n_319), .B1(n_860), .B2(n_1538), .Y(n_1537) );
INVxp33_ASAP7_75t_SL g1506 ( .A(n_149), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_149), .A2(n_353), .B1(n_1018), .B2(n_1533), .Y(n_1532) );
INVxp67_ASAP7_75t_SL g1145 ( .A(n_150), .Y(n_1145) );
INVx1_ASAP7_75t_L g850 ( .A(n_152), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_152), .A2(n_161), .B1(n_581), .B2(n_596), .Y(n_856) );
XNOR2xp5_ASAP7_75t_L g1216 ( .A(n_153), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g414 ( .A(n_155), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_156), .A2(n_355), .B1(n_586), .B2(n_597), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_157), .A2(n_231), .B1(n_1367), .B2(n_1369), .Y(n_1366) );
INVx1_ASAP7_75t_L g1385 ( .A(n_157), .Y(n_1385) );
INVx1_ASAP7_75t_L g780 ( .A(n_158), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_158), .A2(n_313), .B1(n_596), .B2(n_597), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_159), .A2(n_201), .B1(n_391), .B2(n_410), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_159), .A2(n_291), .B1(n_1035), .B2(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g853 ( .A(n_161), .Y(n_853) );
XOR2xp5_ASAP7_75t_L g1798 ( .A(n_162), .B(n_1799), .Y(n_1798) );
AOI22xp33_ASAP7_75t_L g1906 ( .A1(n_162), .A2(n_1907), .B1(n_1911), .B2(n_1950), .Y(n_1906) );
INVx1_ASAP7_75t_L g1565 ( .A(n_163), .Y(n_1565) );
INVxp33_ASAP7_75t_SL g1463 ( .A(n_164), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g1480 ( .A1(n_164), .A2(n_209), .B1(n_519), .B2(n_1481), .Y(n_1480) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_165), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_166), .A2(n_372), .B1(n_391), .B2(n_410), .Y(n_1115) );
INVx1_ASAP7_75t_L g1132 ( .A(n_166), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_167), .A2(n_264), .B1(n_684), .B2(n_687), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_167), .A2(n_264), .B1(n_699), .B2(n_700), .Y(n_698) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_169), .Y(n_957) );
INVx1_ASAP7_75t_L g1589 ( .A(n_170), .Y(n_1589) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_171), .Y(n_422) );
INVx1_ASAP7_75t_L g1512 ( .A(n_172), .Y(n_1512) );
OAI22xp5_ASAP7_75t_L g1517 ( .A1(n_172), .A2(n_303), .B1(n_438), .B2(n_1005), .Y(n_1517) );
OAI211xp5_ASAP7_75t_L g886 ( .A1(n_173), .A2(n_591), .B(n_887), .C(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g911 ( .A(n_173), .Y(n_911) );
AO22x2_ASAP7_75t_SL g1458 ( .A1(n_174), .A2(n_1459), .B1(n_1460), .B2(n_1498), .Y(n_1458) );
CKINVDCx16_ASAP7_75t_R g1459 ( .A(n_174), .Y(n_1459) );
INVx1_ASAP7_75t_L g796 ( .A(n_175), .Y(n_796) );
OAI22xp33_ASAP7_75t_SL g817 ( .A1(n_175), .A2(n_186), .B1(n_391), .B2(n_640), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_176), .A2(n_316), .B1(n_511), .B2(n_1147), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_176), .A2(n_316), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
INVx1_ASAP7_75t_L g1563 ( .A(n_177), .Y(n_1563) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_177), .B(n_1571), .Y(n_1576) );
INVxp67_ASAP7_75t_SL g937 ( .A(n_178), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_179), .A2(n_247), .B1(n_432), .B2(n_1431), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1438 ( .A1(n_179), .A2(n_247), .B1(n_590), .B2(n_751), .Y(n_1438) );
INVxp33_ASAP7_75t_SL g1269 ( .A(n_180), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_180), .A2(n_260), .B1(n_511), .B2(n_692), .Y(n_1292) );
INVxp33_ASAP7_75t_SL g946 ( .A(n_181), .Y(n_946) );
INVxp33_ASAP7_75t_L g1007 ( .A(n_182), .Y(n_1007) );
INVxp67_ASAP7_75t_SL g1224 ( .A(n_183), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1246 ( .A1(n_183), .A2(n_244), .B1(n_1242), .B2(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_L g394 ( .A(n_184), .Y(n_394) );
INVxp33_ASAP7_75t_L g1505 ( .A(n_185), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1535 ( .A1(n_185), .A2(n_343), .B1(n_432), .B2(n_1244), .Y(n_1535) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_186), .A2(n_302), .B1(n_631), .B2(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_SL g1939 ( .A1(n_187), .A2(n_327), .B1(n_487), .B2(n_547), .Y(n_1939) );
INVxp33_ASAP7_75t_SL g1949 ( .A(n_187), .Y(n_1949) );
BUFx3_ASAP7_75t_L g466 ( .A(n_189), .Y(n_466) );
INVx1_ASAP7_75t_L g483 ( .A(n_189), .Y(n_483) );
INVx1_ASAP7_75t_L g1151 ( .A(n_190), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g1163 ( .A1(n_190), .A2(n_372), .B1(n_586), .B2(n_597), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_191), .A2(n_194), .B1(n_1193), .B2(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1213 ( .A(n_191), .Y(n_1213) );
XNOR2xp5_ASAP7_75t_L g1912 ( .A(n_192), .B(n_1913), .Y(n_1912) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_193), .A2(n_256), .B1(n_535), .B2(n_682), .Y(n_743) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_193), .A2(n_256), .B1(n_570), .B2(n_631), .Y(n_753) );
INVx1_ASAP7_75t_L g1210 ( .A(n_194), .Y(n_1210) );
INVx1_ASAP7_75t_L g996 ( .A(n_195), .Y(n_996) );
INVxp33_ASAP7_75t_SL g1808 ( .A(n_196), .Y(n_1808) );
AOI221xp5_ASAP7_75t_L g1856 ( .A1(n_196), .A2(n_311), .B1(n_1857), .B2(n_1858), .C(n_1860), .Y(n_1856) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_197), .A2(n_348), .B1(n_581), .B2(n_596), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_197), .A2(n_348), .B1(n_511), .B2(n_905), .C(n_908), .Y(n_904) );
INVx1_ASAP7_75t_L g718 ( .A(n_198), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_198), .A2(n_328), .B1(n_636), .B2(n_745), .Y(n_748) );
INVxp33_ASAP7_75t_L g443 ( .A(n_199), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_199), .A2(n_262), .B1(n_547), .B2(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g998 ( .A(n_201), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_202), .A2(n_252), .B1(n_511), .B2(n_1477), .Y(n_1476) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_202), .A2(n_252), .B1(n_1039), .B2(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g485 ( .A(n_203), .Y(n_485) );
INVx1_ASAP7_75t_L g1157 ( .A(n_205), .Y(n_1157) );
OAI211xp5_ASAP7_75t_L g1161 ( .A1(n_205), .A2(n_591), .B(n_789), .C(n_1162), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_206), .A2(n_339), .B1(n_532), .B2(n_1184), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_206), .A2(n_339), .B1(n_1033), .B2(n_1195), .Y(n_1194) );
AOI22xp33_ASAP7_75t_SL g1475 ( .A1(n_207), .A2(n_366), .B1(n_519), .B2(n_1294), .Y(n_1475) );
AOI22xp33_ASAP7_75t_SL g1485 ( .A1(n_207), .A2(n_366), .B1(n_487), .B2(n_1041), .Y(n_1485) );
INVx1_ASAP7_75t_L g1469 ( .A(n_209), .Y(n_1469) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_210), .A2(n_306), .B1(n_962), .B2(n_963), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_210), .A2(n_306), .B1(n_511), .B2(n_897), .Y(n_978) );
INVx1_ASAP7_75t_L g1226 ( .A(n_211), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_211), .A2(n_216), .B1(n_731), .B2(n_1244), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_212), .A2(n_1113), .B1(n_1164), .B2(n_1165), .Y(n_1112) );
INVx1_ASAP7_75t_L g1165 ( .A(n_212), .Y(n_1165) );
INVxp33_ASAP7_75t_SL g1917 ( .A(n_213), .Y(n_1917) );
INVx1_ASAP7_75t_L g837 ( .A(n_215), .Y(n_837) );
OAI211xp5_ASAP7_75t_SL g865 ( .A1(n_215), .A2(n_449), .B(n_814), .C(n_866), .Y(n_865) );
INVxp33_ASAP7_75t_SL g1220 ( .A(n_216), .Y(n_1220) );
INVx1_ASAP7_75t_L g1713 ( .A(n_217), .Y(n_1713) );
INVxp33_ASAP7_75t_SL g1317 ( .A(n_218), .Y(n_1317) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_219), .A2(n_308), .B1(n_581), .B2(n_586), .Y(n_580) );
INVx1_ASAP7_75t_L g638 ( .A(n_219), .Y(n_638) );
INVx1_ASAP7_75t_L g738 ( .A(n_220), .Y(n_738) );
INVx1_ASAP7_75t_L g505 ( .A(n_221), .Y(n_505) );
INVx1_ASAP7_75t_L g1867 ( .A(n_221), .Y(n_1867) );
INVx1_ASAP7_75t_L g1127 ( .A(n_222), .Y(n_1127) );
INVxp67_ASAP7_75t_L g677 ( .A(n_223), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_223), .A2(n_315), .B1(n_570), .B2(n_571), .Y(n_711) );
INVx1_ASAP7_75t_L g1426 ( .A(n_224), .Y(n_1426) );
OAI22xp33_ASAP7_75t_L g1448 ( .A1(n_224), .A2(n_341), .B1(n_438), .B2(n_1005), .Y(n_1448) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_225), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_225), .A2(n_342), .B1(n_631), .B2(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g1848 ( .A(n_226), .Y(n_1848) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_227), .A2(n_362), .B1(n_535), .B2(n_682), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_227), .A2(n_362), .B1(n_1129), .B2(n_1301), .Y(n_1439) );
INVx1_ASAP7_75t_L g1392 ( .A(n_228), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_228), .A2(n_233), .B1(n_581), .B2(n_596), .Y(n_1407) );
INVx1_ASAP7_75t_L g1597 ( .A(n_229), .Y(n_1597) );
INVxp67_ASAP7_75t_SL g1840 ( .A(n_230), .Y(n_1840) );
AOI22xp33_ASAP7_75t_L g1884 ( .A1(n_230), .A2(n_317), .B1(n_555), .B2(n_1885), .Y(n_1884) );
INVx1_ASAP7_75t_L g1381 ( .A(n_231), .Y(n_1381) );
AOI22xp5_ASAP7_75t_L g1567 ( .A1(n_232), .A2(n_374), .B1(n_1568), .B2(n_1574), .Y(n_1567) );
INVx1_ASAP7_75t_L g1389 ( .A(n_233), .Y(n_1389) );
CKINVDCx14_ASAP7_75t_R g577 ( .A(n_234), .Y(n_577) );
INVx1_ASAP7_75t_L g593 ( .A(n_235), .Y(n_593) );
INVx1_ASAP7_75t_L g1920 ( .A(n_236), .Y(n_1920) );
INVxp33_ASAP7_75t_SL g1464 ( .A(n_237), .Y(n_1464) );
INVxp33_ASAP7_75t_L g1331 ( .A(n_238), .Y(n_1331) );
INVxp67_ASAP7_75t_SL g1520 ( .A(n_239), .Y(n_1520) );
INVx1_ASAP7_75t_L g839 ( .A(n_240), .Y(n_839) );
INVx1_ASAP7_75t_L g1149 ( .A(n_242), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_243), .Y(n_900) );
INVxp33_ASAP7_75t_SL g1221 ( .A(n_244), .Y(n_1221) );
INVx1_ASAP7_75t_L g1466 ( .A(n_245), .Y(n_1466) );
INVx1_ASAP7_75t_L g769 ( .A(n_246), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_250), .A2(n_324), .B1(n_581), .B2(n_596), .Y(n_1056) );
INVx1_ASAP7_75t_L g1074 ( .A(n_250), .Y(n_1074) );
INVx1_ASAP7_75t_L g606 ( .A(n_255), .Y(n_606) );
INVx1_ASAP7_75t_L g1055 ( .A(n_257), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_259), .Y(n_1364) );
INVxp33_ASAP7_75t_SL g1272 ( .A(n_260), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_261), .A2(n_265), .B1(n_586), .B2(n_597), .Y(n_891) );
INVx1_ASAP7_75t_L g909 ( .A(n_261), .Y(n_909) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_262), .Y(n_430) );
INVx1_ASAP7_75t_L g1926 ( .A(n_263), .Y(n_1926) );
INVx1_ASAP7_75t_L g883 ( .A(n_265), .Y(n_883) );
INVx1_ASAP7_75t_L g953 ( .A(n_267), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_267), .A2(n_314), .B1(n_432), .B2(n_602), .Y(n_980) );
INVxp67_ASAP7_75t_SL g1098 ( .A(n_269), .Y(n_1098) );
INVx1_ASAP7_75t_L g841 ( .A(n_271), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_271), .A2(n_281), .B1(n_410), .B2(n_644), .Y(n_864) );
INVxp33_ASAP7_75t_L g673 ( .A(n_273), .Y(n_673) );
INVx1_ASAP7_75t_L g943 ( .A(n_274), .Y(n_943) );
INVxp33_ASAP7_75t_L g1497 ( .A(n_275), .Y(n_1497) );
BUFx3_ASAP7_75t_L g468 ( .A(n_276), .Y(n_468) );
INVx1_ASAP7_75t_L g474 ( .A(n_276), .Y(n_474) );
INVxp67_ASAP7_75t_SL g1921 ( .A(n_277), .Y(n_1921) );
AOI22xp33_ASAP7_75t_L g1933 ( .A1(n_277), .A2(n_285), .B1(n_511), .B2(n_602), .Y(n_1933) );
INVx1_ASAP7_75t_L g629 ( .A(n_278), .Y(n_629) );
INVx1_ASAP7_75t_L g1419 ( .A(n_279), .Y(n_1419) );
INVx1_ASAP7_75t_L g1372 ( .A(n_280), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_280), .A2(n_336), .B1(n_391), .B2(n_410), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_281), .A2(n_287), .B1(n_586), .B2(n_597), .Y(n_857) );
INVx1_ASAP7_75t_L g1424 ( .A(n_282), .Y(n_1424) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_283), .Y(n_390) );
INVx1_ASAP7_75t_L g544 ( .A(n_283), .Y(n_544) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_283), .B(n_413), .Y(n_1807) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_283), .B(n_346), .Y(n_1823) );
AOI221xp5_ASAP7_75t_SL g896 ( .A1(n_284), .A2(n_294), .B1(n_897), .B2(n_898), .C(n_899), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_284), .A2(n_294), .B1(n_919), .B2(n_920), .Y(n_918) );
INVxp33_ASAP7_75t_SL g1918 ( .A(n_285), .Y(n_1918) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_286), .Y(n_809) );
INVx1_ASAP7_75t_L g851 ( .A(n_287), .Y(n_851) );
INVx1_ASAP7_75t_L g1054 ( .A(n_288), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_290), .B(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g461 ( .A(n_292), .Y(n_461) );
OR2x2_ASAP7_75t_L g1866 ( .A(n_292), .B(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g650 ( .A(n_293), .Y(n_650) );
INVx1_ASAP7_75t_L g1508 ( .A(n_295), .Y(n_1508) );
INVx1_ASAP7_75t_L g1324 ( .A(n_296), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_296), .A2(n_332), .B1(n_670), .B2(n_671), .Y(n_1329) );
INVx1_ASAP7_75t_L g862 ( .A(n_298), .Y(n_862) );
INVxp67_ASAP7_75t_L g1237 ( .A(n_299), .Y(n_1237) );
OAI211xp5_ASAP7_75t_L g1050 ( .A1(n_300), .A2(n_591), .B(n_1051), .C(n_1053), .Y(n_1050) );
INVx1_ASAP7_75t_L g1075 ( .A(n_300), .Y(n_1075) );
OAI211xp5_ASAP7_75t_L g1177 ( .A1(n_301), .A2(n_591), .B(n_797), .C(n_1178), .Y(n_1177) );
AOI22xp33_ASAP7_75t_SL g1190 ( .A1(n_301), .A2(n_351), .B1(n_520), .B2(n_731), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_302), .A2(n_340), .B1(n_410), .B2(n_644), .Y(n_812) );
INVx1_ASAP7_75t_L g1513 ( .A(n_303), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_304), .Y(n_901) );
INVx1_ASAP7_75t_L g1843 ( .A(n_305), .Y(n_1843) );
INVx1_ASAP7_75t_L g1284 ( .A(n_307), .Y(n_1284) );
INVx1_ASAP7_75t_L g613 ( .A(n_308), .Y(n_613) );
INVxp33_ASAP7_75t_SL g1282 ( .A(n_309), .Y(n_1282) );
INVx1_ASAP7_75t_L g1223 ( .A(n_310), .Y(n_1223) );
INVxp33_ASAP7_75t_L g1811 ( .A(n_311), .Y(n_1811) );
INVxp67_ASAP7_75t_SL g1516 ( .A(n_312), .Y(n_1516) );
INVx1_ASAP7_75t_L g778 ( .A(n_313), .Y(n_778) );
INVxp33_ASAP7_75t_SL g951 ( .A(n_314), .Y(n_951) );
INVx1_ASAP7_75t_L g674 ( .A(n_315), .Y(n_674) );
INVxp33_ASAP7_75t_L g1832 ( .A(n_317), .Y(n_1832) );
INVx1_ASAP7_75t_L g799 ( .A(n_318), .Y(n_799) );
OAI211xp5_ASAP7_75t_SL g813 ( .A1(n_318), .A2(n_449), .B(n_814), .C(n_816), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_320), .A2(n_344), .B1(n_659), .B2(n_662), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_320), .A2(n_344), .B1(n_670), .B2(n_671), .Y(n_669) );
INVxp67_ASAP7_75t_SL g1234 ( .A(n_321), .Y(n_1234) );
INVx1_ASAP7_75t_L g1472 ( .A(n_323), .Y(n_1472) );
INVx1_ASAP7_75t_L g1067 ( .A(n_324), .Y(n_1067) );
INVx1_ASAP7_75t_L g737 ( .A(n_325), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_325), .A2(n_350), .B1(n_575), .B2(n_751), .Y(n_755) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_326), .Y(n_999) );
INVxp67_ASAP7_75t_SL g1943 ( .A(n_327), .Y(n_1943) );
INVx1_ASAP7_75t_L g725 ( .A(n_328), .Y(n_725) );
INVx1_ASAP7_75t_L g405 ( .A(n_329), .Y(n_405) );
INVx1_ASAP7_75t_L g829 ( .A(n_331), .Y(n_829) );
INVx1_ASAP7_75t_L g1323 ( .A(n_332), .Y(n_1323) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_333), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_333), .A2(n_349), .B1(n_532), .B2(n_533), .Y(n_531) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_335), .Y(n_384) );
AND3x2_ASAP7_75t_L g1564 ( .A(n_335), .B(n_382), .C(n_1565), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_335), .B(n_382), .Y(n_1573) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_336), .A2(n_359), .B1(n_586), .B2(n_597), .Y(n_1408) );
INVx2_ASAP7_75t_L g395 ( .A(n_337), .Y(n_395) );
INVx1_ASAP7_75t_L g1121 ( .A(n_338), .Y(n_1121) );
INVx1_ASAP7_75t_L g1425 ( .A(n_341), .Y(n_1425) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_342), .Y(n_771) );
INVxp67_ASAP7_75t_SL g1511 ( .A(n_343), .Y(n_1511) );
INVx1_ASAP7_75t_L g766 ( .A(n_345), .Y(n_766) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
INVx2_ASAP7_75t_L g413 ( .A(n_346), .Y(n_413) );
XNOR2xp5_ASAP7_75t_L g714 ( .A(n_347), .B(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_349), .Y(n_479) );
INVx1_ASAP7_75t_L g730 ( .A(n_350), .Y(n_730) );
INVx1_ASAP7_75t_L g1849 ( .A(n_352), .Y(n_1849) );
INVxp33_ASAP7_75t_L g1509 ( .A(n_353), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_354), .Y(n_880) );
INVx1_ASAP7_75t_L g1070 ( .A(n_355), .Y(n_1070) );
AO22x2_ASAP7_75t_L g931 ( .A1(n_357), .A2(n_932), .B1(n_933), .B2(n_981), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_357), .Y(n_932) );
INVx1_ASAP7_75t_L g1119 ( .A(n_358), .Y(n_1119) );
INVx1_ASAP7_75t_L g1397 ( .A(n_359), .Y(n_1397) );
INVx1_ASAP7_75t_L g1179 ( .A(n_360), .Y(n_1179) );
XOR2x2_ASAP7_75t_L g1312 ( .A(n_361), .B(n_1313), .Y(n_1312) );
INVxp33_ASAP7_75t_SL g1946 ( .A(n_363), .Y(n_1946) );
INVxp33_ASAP7_75t_SL g1803 ( .A(n_364), .Y(n_1803) );
INVx1_ASAP7_75t_L g723 ( .A(n_365), .Y(n_723) );
INVx1_ASAP7_75t_L g1453 ( .A(n_367), .Y(n_1453) );
INVxp33_ASAP7_75t_SL g1834 ( .A(n_368), .Y(n_1834) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_369), .A2(n_373), .B1(n_923), .B2(n_1488), .Y(n_1487) );
INVxp33_ASAP7_75t_L g1494 ( .A(n_369), .Y(n_1494) );
INVx1_ASAP7_75t_L g784 ( .A(n_371), .Y(n_784) );
INVxp67_ASAP7_75t_SL g1495 ( .A(n_373), .Y(n_1495) );
AO22x1_ASAP7_75t_L g1500 ( .A1(n_374), .A2(n_1501), .B1(n_1502), .B2(n_1548), .Y(n_1500) );
INVxp67_ASAP7_75t_L g1501 ( .A(n_374), .Y(n_1501) );
INVxp67_ASAP7_75t_SL g1227 ( .A(n_375), .Y(n_1227) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_398), .B(n_1551), .Y(n_376) );
BUFx12f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_385), .Y(n_379) );
AND2x4_ASAP7_75t_L g1905 ( .A(n_380), .B(n_386), .Y(n_1905) );
NOR2xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_SL g1910 ( .A(n_381), .Y(n_1910) );
NAND2xp5_ASAP7_75t_L g1955 ( .A(n_381), .B(n_383), .Y(n_1955) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g1909 ( .A(n_383), .B(n_1910), .Y(n_1909) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_391), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x6_ASAP7_75t_L g453 ( .A(n_388), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g678 ( .A(n_388), .B(n_454), .Y(n_678) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g529 ( .A(n_389), .B(n_397), .Y(n_529) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g763 ( .A(n_390), .B(n_412), .Y(n_763) );
INVx8_ASAP7_75t_L g442 ( .A(n_391), .Y(n_442) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
OR2x6_ASAP7_75t_L g410 ( .A(n_392), .B(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_392), .Y(n_605) );
INVx2_ASAP7_75t_SL g615 ( .A(n_392), .Y(n_615) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_392), .Y(n_765) );
INVx2_ASAP7_75t_SL g846 ( .A(n_392), .Y(n_846) );
INVx1_ASAP7_75t_L g1155 ( .A(n_392), .Y(n_1155) );
OR2x2_ASAP7_75t_L g1896 ( .A(n_392), .B(n_1822), .Y(n_1896) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
INVx1_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
INVx1_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
AND2x4_ASAP7_75t_L g447 ( .A(n_394), .B(n_435), .Y(n_447) );
AND2x2_ASAP7_75t_L g522 ( .A(n_394), .B(n_395), .Y(n_522) );
INVx1_ASAP7_75t_L g419 ( .A(n_395), .Y(n_419) );
INVx2_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
INVx1_ASAP7_75t_L g609 ( .A(n_395), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_395), .B(n_417), .Y(n_643) );
AND2x4_ASAP7_75t_L g439 ( .A(n_396), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g671 ( .A(n_397), .B(n_425), .Y(n_671) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_397), .B(n_425), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_1167), .B1(n_1168), .B2(n_1550), .Y(n_398) );
INVx1_ASAP7_75t_L g1550 ( .A(n_399), .Y(n_1550) );
AO22x2_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_983), .B2(n_984), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XOR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_870), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_646), .Y(n_402) );
XNOR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_576), .Y(n_403) );
XNOR2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_452), .B1(n_455), .B2(n_501), .C(n_508), .Y(n_406) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_408), .B(n_421), .C(n_441), .D(n_449), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_414), .B1(n_415), .B2(n_420), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_409), .A2(n_442), .B1(n_628), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_409), .A2(n_442), .B1(n_946), .B2(n_947), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_409), .A2(n_442), .B1(n_1213), .B2(n_1214), .Y(n_1212) );
AOI22xp33_ASAP7_75t_SL g1452 ( .A1(n_409), .A2(n_442), .B1(n_1418), .B2(n_1453), .Y(n_1452) );
AOI22xp33_ASAP7_75t_SL g1948 ( .A1(n_409), .A2(n_442), .B1(n_1920), .B2(n_1949), .Y(n_1948) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx5_ASAP7_75t_L g676 ( .A(n_410), .Y(n_676) );
AND2x4_ASAP7_75t_L g415 ( .A(n_411), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g444 ( .A(n_411), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g641 ( .A(n_411), .Y(n_641) );
AND2x4_ASAP7_75t_L g645 ( .A(n_411), .B(n_445), .Y(n_645) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g429 ( .A(n_413), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_414), .A2(n_476), .B1(n_479), .B2(n_480), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_415), .A2(n_442), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_415), .A2(n_442), .B1(n_737), .B2(n_738), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_415), .A2(n_645), .B1(n_936), .B2(n_937), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_415), .A2(n_444), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
AOI22xp5_ASAP7_75t_SL g1236 ( .A1(n_415), .A2(n_645), .B1(n_1237), .B2(n_1238), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_415), .A2(n_645), .B1(n_1281), .B2(n_1282), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_415), .A2(n_444), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
AOI22xp33_ASAP7_75t_SL g1449 ( .A1(n_415), .A2(n_444), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_415), .A2(n_645), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_415), .A2(n_444), .B1(n_1519), .B2(n_1520), .Y(n_1518) );
AOI22xp33_ASAP7_75t_L g1945 ( .A1(n_415), .A2(n_645), .B1(n_1946), .B2(n_1947), .Y(n_1945) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_416), .Y(n_513) );
BUFx2_ASAP7_75t_L g532 ( .A(n_416), .Y(n_532) );
BUFx2_ASAP7_75t_L g601 ( .A(n_416), .Y(n_601) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_416), .Y(n_682) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_416), .Y(n_691) );
INVx1_ASAP7_75t_L g1019 ( .A(n_416), .Y(n_1019) );
INVx1_ASAP7_75t_L g1026 ( .A(n_416), .Y(n_1026) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g1827 ( .A(n_417), .Y(n_1827) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_430), .B2(n_431), .C1(n_436), .C2(n_437), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g484 ( .A1(n_422), .A2(n_436), .B1(n_485), .B2(n_486), .C1(n_490), .C2(n_495), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_423), .A2(n_439), .B1(n_593), .B2(n_594), .C1(n_629), .C2(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_423), .A2(n_439), .B1(n_808), .B2(n_809), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_423), .A2(n_439), .B1(n_861), .B2(n_862), .Y(n_866) );
AOI222xp33_ASAP7_75t_L g877 ( .A1(n_423), .A2(n_432), .B1(n_439), .B2(n_878), .C1(n_879), .C2(n_880), .Y(n_877) );
AOI222xp33_ASAP7_75t_L g938 ( .A1(n_423), .A2(n_439), .B1(n_939), .B2(n_940), .C1(n_943), .C2(n_944), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_423), .A2(n_437), .B1(n_1054), .B2(n_1055), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_423), .A2(n_1119), .B1(n_1120), .B2(n_1121), .Y(n_1118) );
AOI222xp33_ASAP7_75t_L g1283 ( .A1(n_423), .A2(n_439), .B1(n_731), .B2(n_1275), .C1(n_1278), .C2(n_1284), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_423), .A2(n_439), .B1(n_1403), .B2(n_1404), .Y(n_1402) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
AND2x4_ASAP7_75t_L g1211 ( .A(n_424), .B(n_427), .Y(n_1211) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g608 ( .A(n_426), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_426), .B(n_609), .Y(n_768) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g451 ( .A(n_428), .Y(n_451) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_429), .B(n_544), .Y(n_543) );
AOI211xp5_ASAP7_75t_L g1446 ( .A1(n_431), .A2(n_450), .B(n_1447), .C(n_1448), .Y(n_1446) );
AOI211xp5_ASAP7_75t_L g1515 ( .A1(n_431), .A2(n_450), .B(n_1516), .C(n_1517), .Y(n_1515) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g538 ( .A(n_432), .Y(n_538) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g450 ( .A(n_433), .B(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g524 ( .A(n_433), .Y(n_524) );
BUFx3_ASAP7_75t_L g636 ( .A(n_433), .Y(n_636) );
INVx1_ASAP7_75t_L g688 ( .A(n_433), .Y(n_688) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_433), .Y(n_733) );
BUFx2_ASAP7_75t_L g942 ( .A(n_433), .Y(n_942) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g670 ( .A(n_439), .Y(n_670) );
INVx2_ASAP7_75t_L g735 ( .A(n_439), .Y(n_735) );
AOI222xp33_ASAP7_75t_L g1209 ( .A1(n_439), .A2(n_733), .B1(n_1179), .B2(n_1180), .C1(n_1210), .C2(n_1211), .Y(n_1209) );
INVx1_ASAP7_75t_L g1820 ( .A(n_440), .Y(n_1820) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .B1(n_444), .B2(n_448), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_442), .A2(n_676), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g1231 ( .A1(n_442), .A2(n_676), .B1(n_1223), .B2(n_1232), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_442), .A2(n_676), .B1(n_1271), .B2(n_1286), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_442), .A2(n_676), .B1(n_1319), .B2(n_1334), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_442), .A2(n_676), .B1(n_1466), .B2(n_1497), .Y(n_1496) );
AOI22xp33_ASAP7_75t_SL g1521 ( .A1(n_442), .A2(n_676), .B1(n_1508), .B2(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_446), .Y(n_693) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g517 ( .A(n_447), .Y(n_517) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_447), .Y(n_535) );
INVx1_ASAP7_75t_L g1023 ( .A(n_447), .Y(n_1023) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_449), .B(n_634), .C(n_637), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_449), .B(n_877), .C(n_881), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g934 ( .A(n_449), .B(n_935), .C(n_938), .D(n_945), .Y(n_934) );
NAND3xp33_ASAP7_75t_L g1208 ( .A(n_449), .B(n_1209), .C(n_1212), .Y(n_1208) );
NAND4xp25_ASAP7_75t_SL g1279 ( .A(n_449), .B(n_1280), .C(n_1283), .D(n_1285), .Y(n_1279) );
CKINVDCx11_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_450), .A2(n_635), .B(n_668), .C(n_669), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_450), .A2(n_730), .B(n_731), .C(n_734), .Y(n_729) );
NOR3xp33_ASAP7_75t_L g1002 ( .A(n_450), .B(n_1003), .C(n_1004), .Y(n_1002) );
AOI211xp5_ASAP7_75t_L g1233 ( .A1(n_450), .A2(n_687), .B(n_1234), .C(n_1235), .Y(n_1233) );
AOI211xp5_ASAP7_75t_L g1326 ( .A1(n_450), .A2(n_1327), .B(n_1328), .C(n_1329), .Y(n_1326) );
AOI211xp5_ASAP7_75t_L g1490 ( .A1(n_450), .A2(n_523), .B(n_1491), .C(n_1492), .Y(n_1490) );
AOI211xp5_ASAP7_75t_SL g1942 ( .A1(n_450), .A2(n_687), .B(n_1943), .C(n_1944), .Y(n_1942) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_452), .A2(n_633), .B(n_639), .Y(n_632) );
OAI31xp33_ASAP7_75t_SL g811 ( .A1(n_452), .A2(n_812), .A3(n_813), .B(n_817), .Y(n_811) );
OAI31xp33_ASAP7_75t_SL g863 ( .A1(n_452), .A2(n_864), .A3(n_865), .B(n_867), .Y(n_863) );
O2A1O1Ixp33_ASAP7_75t_L g874 ( .A1(n_452), .A2(n_875), .B(n_876), .C(n_884), .Y(n_874) );
AOI221x1_ASAP7_75t_L g933 ( .A1(n_452), .A2(n_503), .B1(n_934), .B2(n_948), .C(n_958), .Y(n_933) );
OAI31xp33_ASAP7_75t_L g1057 ( .A1(n_452), .A2(n_1058), .A3(n_1059), .B(n_1063), .Y(n_1057) );
OAI31xp33_ASAP7_75t_L g1114 ( .A1(n_452), .A2(n_1115), .A3(n_1116), .B(n_1122), .Y(n_1114) );
OAI21xp5_ASAP7_75t_L g1207 ( .A1(n_452), .A2(n_1208), .B(n_1215), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_452), .A2(n_503), .B1(n_1266), .B2(n_1279), .C(n_1287), .Y(n_1265) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_452), .A2(n_503), .B1(n_1314), .B2(n_1325), .C(n_1335), .Y(n_1313) );
OAI31xp33_ASAP7_75t_SL g1399 ( .A1(n_452), .A2(n_1400), .A3(n_1401), .B(n_1405), .Y(n_1399) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
AOI31xp33_ASAP7_75t_L g1230 ( .A1(n_453), .A2(n_1231), .A3(n_1233), .B(n_1236), .Y(n_1230) );
AOI31xp33_ASAP7_75t_L g1445 ( .A1(n_453), .A2(n_1446), .A3(n_1449), .B(n_1452), .Y(n_1445) );
AOI31xp33_ASAP7_75t_L g1489 ( .A1(n_453), .A2(n_1490), .A3(n_1493), .B(n_1496), .Y(n_1489) );
AOI31xp33_ASAP7_75t_L g1514 ( .A1(n_453), .A2(n_1515), .A3(n_1518), .B(n_1521), .Y(n_1514) );
AOI31xp33_ASAP7_75t_L g1941 ( .A1(n_453), .A2(n_1942), .A3(n_1945), .B(n_1948), .Y(n_1941) );
AND2x4_ASAP7_75t_L g564 ( .A(n_454), .B(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g712 ( .A(n_454), .B(n_565), .Y(n_712) );
AND2x4_ASAP7_75t_L g1898 ( .A(n_454), .B(n_1899), .Y(n_1898) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_475), .C(n_484), .D(n_497), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_469), .B2(n_470), .Y(n_456) );
AOI22xp5_ASAP7_75t_SL g653 ( .A1(n_458), .A2(n_476), .B1(n_654), .B2(n_655), .Y(n_653) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_458), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_458), .A2(n_470), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_458), .A2(n_470), .B1(n_1268), .B2(n_1269), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_458), .A2(n_470), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_458), .A2(n_470), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_458), .A2(n_470), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_462), .Y(n_458) );
AND2x6_ASAP7_75t_L g480 ( .A(n_459), .B(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g719 ( .A(n_459), .B(n_462), .Y(n_719) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g660 ( .A(n_460), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g472 ( .A(n_461), .Y(n_472) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_461), .Y(n_478) );
AND2x2_ASAP7_75t_L g560 ( .A(n_461), .B(n_505), .Y(n_560) );
INVx2_ASAP7_75t_L g566 ( .A(n_461), .Y(n_566) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g548 ( .A(n_463), .Y(n_548) );
INVx1_ASAP7_75t_L g699 ( .A(n_463), .Y(n_699) );
INVx2_ASAP7_75t_L g970 ( .A(n_463), .Y(n_970) );
BUFx6f_ASAP7_75t_L g1038 ( .A(n_463), .Y(n_1038) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_463), .Y(n_1201) );
INVx2_ASAP7_75t_SL g1540 ( .A(n_463), .Y(n_1540) );
INVx6_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g476 ( .A(n_464), .B(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g710 ( .A(n_464), .Y(n_710) );
INVx2_ASAP7_75t_L g752 ( .A(n_464), .Y(n_752) );
AND2x2_ASAP7_75t_L g1899 ( .A(n_464), .B(n_1871), .Y(n_1899) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g496 ( .A(n_465), .Y(n_496) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g473 ( .A(n_466), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g489 ( .A(n_466), .B(n_468), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g482 ( .A(n_468), .B(n_483), .Y(n_482) );
CKINVDCx6p67_ASAP7_75t_R g596 ( .A(n_470), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_470), .A2(n_480), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_470), .A2(n_480), .B1(n_722), .B2(n_723), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_470), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1504 ( .A1(n_470), .A2(n_719), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
AOI22xp33_ASAP7_75t_L g1916 ( .A1(n_470), .A2(n_719), .B1(n_1917), .B2(n_1918), .Y(n_1916) );
AND2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
INVx1_ASAP7_75t_L g582 ( .A(n_471), .Y(n_582) );
AND2x2_ASAP7_75t_L g589 ( .A(n_471), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x6_ASAP7_75t_L g495 ( .A(n_472), .B(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
BUFx3_ASAP7_75t_L g570 ( .A(n_473), .Y(n_570) );
INVx2_ASAP7_75t_SL g704 ( .A(n_473), .Y(n_704) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_473), .Y(n_793) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_473), .Y(n_801) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_473), .Y(n_825) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_473), .Y(n_1043) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_473), .Y(n_1092) );
HB1xp67_ASAP7_75t_L g1484 ( .A(n_473), .Y(n_1484) );
HB1xp67_ASAP7_75t_L g1546 ( .A(n_473), .Y(n_1546) );
INVx1_ASAP7_75t_L g585 ( .A(n_474), .Y(n_585) );
INVx4_ASAP7_75t_L g586 ( .A(n_476), .Y(n_586) );
AOI22xp5_ASAP7_75t_SL g717 ( .A1(n_476), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_476), .A2(n_480), .B1(n_947), .B2(n_951), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_476), .A2(n_480), .B1(n_998), .B2(n_999), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_476), .A2(n_480), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_476), .A2(n_480), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_476), .A2(n_480), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
AOI22xp5_ASAP7_75t_L g1417 ( .A1(n_476), .A2(n_480), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g1465 ( .A1(n_476), .A2(n_480), .B1(n_1466), .B2(n_1467), .Y(n_1465) );
AOI22xp33_ASAP7_75t_L g1507 ( .A1(n_476), .A2(n_480), .B1(n_1508), .B2(n_1509), .Y(n_1507) );
AOI22xp33_ASAP7_75t_L g1919 ( .A1(n_476), .A2(n_480), .B1(n_1920), .B2(n_1921), .Y(n_1919) );
AND2x4_ASAP7_75t_L g491 ( .A(n_477), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_SL g1228 ( .A(n_477), .B(n_492), .Y(n_1228) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g597 ( .A(n_480), .Y(n_597) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_481), .Y(n_571) );
INVx2_ASAP7_75t_L g840 ( .A(n_481), .Y(n_840) );
INVx1_ASAP7_75t_L g1094 ( .A(n_481), .Y(n_1094) );
INVx1_ASAP7_75t_L g1260 ( .A(n_481), .Y(n_1260) );
BUFx6f_ASAP7_75t_L g1301 ( .A(n_481), .Y(n_1301) );
INVx1_ASAP7_75t_L g1444 ( .A(n_481), .Y(n_1444) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g556 ( .A(n_482), .Y(n_556) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_482), .Y(n_631) );
INVx2_ASAP7_75t_L g966 ( .A(n_482), .Y(n_966) );
INVx1_ASAP7_75t_L g584 ( .A(n_483), .Y(n_584) );
AOI222xp33_ASAP7_75t_L g952 ( .A1(n_486), .A2(n_490), .B1(n_495), .B2(n_943), .C1(n_944), .C2(n_953), .Y(n_952) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx4f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_488), .Y(n_575) );
INVx2_ASAP7_75t_SL g807 ( .A(n_488), .Y(n_807) );
BUFx3_ASAP7_75t_L g1193 ( .A(n_488), .Y(n_1193) );
INVx1_ASAP7_75t_L g1309 ( .A(n_488), .Y(n_1309) );
AND2x4_ASAP7_75t_L g1879 ( .A(n_488), .B(n_1865), .Y(n_1879) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_489), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_490), .A2(n_495), .B1(n_878), .B2(n_880), .Y(n_889) );
AOI222xp33_ASAP7_75t_L g1468 ( .A1(n_490), .A2(n_495), .B1(n_1469), .B2(n_1470), .C1(n_1471), .C2(n_1472), .Y(n_1468) );
AOI222xp33_ASAP7_75t_L g1922 ( .A1(n_490), .A2(n_495), .B1(n_1923), .B2(n_1924), .C1(n_1925), .C2(n_1926), .Y(n_1922) );
BUFx4f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_491), .A2(n_495), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_491), .A2(n_495), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_491), .A2(n_495), .B1(n_1119), .B2(n_1121), .Y(n_1162) );
AOI22xp33_ASAP7_75t_SL g1178 ( .A1(n_491), .A2(n_495), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
INVx1_ASAP7_75t_L g1277 ( .A(n_491), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_491), .A2(n_495), .B1(n_1403), .B2(n_1404), .Y(n_1410) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g661 ( .A(n_493), .Y(n_661) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g1102 ( .A(n_494), .Y(n_1102) );
INVx3_ASAP7_75t_L g662 ( .A(n_495), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g805 ( .A1(n_495), .A2(n_660), .B1(n_784), .B2(n_806), .C1(n_808), .C2(n_809), .Y(n_805) );
AOI222xp33_ASAP7_75t_L g859 ( .A1(n_495), .A2(n_660), .B1(n_854), .B2(n_860), .C1(n_861), .C2(n_862), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_495), .A2(n_660), .B1(n_995), .B2(n_996), .Y(n_994) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_495), .A2(n_573), .B1(n_1226), .B2(n_1227), .C1(n_1228), .C2(n_1229), .Y(n_1225) );
AOI222xp33_ASAP7_75t_L g1273 ( .A1(n_495), .A2(n_1193), .B1(n_1274), .B2(n_1275), .C1(n_1276), .C2(n_1278), .Y(n_1273) );
AOI222xp33_ASAP7_75t_L g1321 ( .A1(n_495), .A2(n_1228), .B1(n_1252), .B2(n_1322), .C1(n_1323), .C2(n_1324), .Y(n_1321) );
AOI222xp33_ASAP7_75t_L g1423 ( .A1(n_495), .A2(n_1193), .B1(n_1228), .B2(n_1424), .C1(n_1425), .C2(n_1426), .Y(n_1423) );
AOI222xp33_ASAP7_75t_L g1510 ( .A1(n_495), .A2(n_575), .B1(n_1228), .B2(n_1511), .C1(n_1512), .C2(n_1513), .Y(n_1510) );
BUFx3_ASAP7_75t_L g1104 ( .A(n_496), .Y(n_1104) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_497), .B(n_653), .C(n_656), .D(n_663), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_497), .B(n_717), .C(n_721), .D(n_724), .Y(n_716) );
BUFx2_ASAP7_75t_L g949 ( .A(n_497), .Y(n_949) );
NAND4xp25_ASAP7_75t_L g1266 ( .A(n_497), .B(n_1267), .C(n_1270), .D(n_1273), .Y(n_1266) );
NAND4xp25_ASAP7_75t_L g1416 ( .A(n_497), .B(n_1417), .C(n_1420), .D(n_1423), .Y(n_1416) );
NAND4xp25_ASAP7_75t_SL g1461 ( .A(n_497), .B(n_1462), .C(n_1465), .D(n_1468), .Y(n_1461) );
NAND4xp25_ASAP7_75t_SL g1503 ( .A(n_497), .B(n_1504), .C(n_1507), .D(n_1510), .Y(n_1503) );
NAND4xp25_ASAP7_75t_SL g1915 ( .A(n_497), .B(n_1916), .C(n_1919), .D(n_1922), .Y(n_1915) );
INVx5_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
CKINVDCx8_ASAP7_75t_R g591 ( .A(n_498), .Y(n_591) );
NOR2xp33_ASAP7_75t_SL g992 ( .A(n_498), .B(n_993), .Y(n_992) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g550 ( .A(n_500), .Y(n_550) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_500), .Y(n_590) );
INVx1_ASAP7_75t_L g701 ( .A(n_500), .Y(n_701) );
BUFx6f_ASAP7_75t_L g1253 ( .A(n_500), .Y(n_1253) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_503), .Y(n_894) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_503), .A2(n_991), .B(n_1000), .Y(n_990) );
AO211x2_ASAP7_75t_L g1217 ( .A1(n_503), .A2(n_1218), .B(n_1230), .C(n_1239), .Y(n_1217) );
OAI31xp33_ASAP7_75t_SL g1406 ( .A1(n_503), .A2(n_1407), .A3(n_1408), .B(n_1409), .Y(n_1406) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x4_ASAP7_75t_L g598 ( .A(n_504), .B(n_506), .Y(n_598) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g565 ( .A(n_505), .B(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
OR2x6_ASAP7_75t_L g762 ( .A(n_507), .B(n_763), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_530), .C(n_545), .D(n_561), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .C(n_525), .Y(n_509) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g1814 ( .A(n_513), .B(n_1806), .Y(n_1814) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g779 ( .A(n_516), .Y(n_779) );
BUFx3_ASAP7_75t_L g897 ( .A(n_516), .Y(n_897) );
AND2x4_ASAP7_75t_L g1805 ( .A(n_516), .B(n_1806), .Y(n_1805) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g776 ( .A(n_517), .Y(n_776) );
BUFx6f_ASAP7_75t_L g1029 ( .A(n_517), .Y(n_1029) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_521), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_521), .Y(n_1529) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_522), .Y(n_686) );
HB1xp67_ASAP7_75t_L g1327 ( .A(n_523), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1016 ( .A(n_524), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_525), .A2(n_896), .B1(n_904), .B2(n_914), .C(n_916), .Y(n_895) );
AOI33xp33_ASAP7_75t_L g976 ( .A1(n_525), .A2(n_914), .A3(n_977), .B1(n_978), .B2(n_979), .B3(n_980), .Y(n_976) );
AOI33xp33_ASAP7_75t_L g1474 ( .A1(n_525), .A2(n_617), .A3(n_1475), .B1(n_1476), .B2(n_1479), .B3(n_1480), .Y(n_1474) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g610 ( .A(n_527), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_527), .B(n_681), .C(n_683), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_527), .B(n_743), .C(n_744), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g1240 ( .A(n_527), .B(n_1241), .C(n_1243), .Y(n_1240) );
NAND3xp33_ASAP7_75t_L g1339 ( .A(n_527), .B(n_1340), .C(n_1344), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g1428 ( .A(n_527), .B(n_1429), .C(n_1430), .Y(n_1428) );
NAND3xp33_ASAP7_75t_L g1524 ( .A(n_527), .B(n_1525), .C(n_1527), .Y(n_1524) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
OR2x6_ASAP7_75t_L g558 ( .A(n_528), .B(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g619 ( .A(n_528), .B(n_559), .Y(n_619) );
AND2x2_ASAP7_75t_L g695 ( .A(n_528), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g706 ( .A(n_528), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_528), .B(n_529), .Y(n_1010) );
INVx2_ASAP7_75t_L g1853 ( .A(n_528), .Y(n_1853) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .C(n_539), .Y(n_530) );
HB1xp67_ASAP7_75t_L g898 ( .A(n_532), .Y(n_898) );
INVxp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
INVx4_ASAP7_75t_L g1185 ( .A(n_535), .Y(n_1185) );
INVx2_ASAP7_75t_SL g1478 ( .A(n_535), .Y(n_1478) );
INVx2_ASAP7_75t_SL g1932 ( .A(n_535), .Y(n_1932) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_538), .Y(n_1294) );
CKINVDCx8_ASAP7_75t_R g915 ( .A(n_539), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g1188 ( .A(n_539), .B(n_1189), .C(n_1190), .Y(n_1188) );
NAND3xp33_ASAP7_75t_L g1245 ( .A(n_539), .B(n_1246), .C(n_1249), .Y(n_1245) );
NAND3xp33_ASAP7_75t_L g1336 ( .A(n_539), .B(n_1337), .C(n_1338), .Y(n_1336) );
NAND3xp33_ASAP7_75t_L g1531 ( .A(n_539), .B(n_1532), .C(n_1535), .Y(n_1531) );
INVx5_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx6_ASAP7_75t_L g617 ( .A(n_540), .Y(n_617) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g1806 ( .A(n_542), .B(n_1807), .Y(n_1806) );
INVx2_ASAP7_75t_L g696 ( .A(n_543), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .C(n_557), .Y(n_545) );
BUFx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_548), .Y(n_926) );
HB1xp67_ASAP7_75t_L g1885 ( .A(n_548), .Y(n_1885) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g860 ( .A(n_550), .Y(n_860) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_553), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_838) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g919 ( .A(n_554), .Y(n_919) );
INVx2_ASAP7_75t_SL g1368 ( .A(n_554), .Y(n_1368) );
AND2x4_ASAP7_75t_L g1864 ( .A(n_554), .B(n_1865), .Y(n_1864) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g1039 ( .A(n_556), .Y(n_1039) );
INVx1_ASAP7_75t_L g1205 ( .A(n_556), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g916 ( .A1(n_558), .A2(n_563), .B1(n_917), .B2(n_921), .Y(n_916) );
INVx2_ASAP7_75t_L g960 ( .A(n_558), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_558), .A2(n_1087), .B1(n_1125), .B2(n_1130), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_558), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_558), .A2(n_563), .B1(n_1363), .B2(n_1370), .Y(n_1362) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g707 ( .A(n_560), .Y(n_707) );
INVx1_ASAP7_75t_L g1883 ( .A(n_560), .Y(n_1883) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_567), .C(n_572), .Y(n_561) );
AOI33xp33_ASAP7_75t_L g959 ( .A1(n_562), .A2(n_960), .A3(n_961), .B1(n_967), .B2(n_972), .B3(n_973), .Y(n_959) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_SL g618 ( .A1(n_563), .A2(n_619), .B1(n_620), .B2(n_627), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g786 ( .A1(n_563), .A2(n_706), .B1(n_787), .B2(n_794), .Y(n_786) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx4f_ASAP7_75t_L g1044 ( .A(n_564), .Y(n_1044) );
BUFx4f_ASAP7_75t_L g1206 ( .A(n_564), .Y(n_1206) );
AOI33xp33_ASAP7_75t_L g1295 ( .A1(n_564), .A2(n_1296), .A3(n_1297), .B1(n_1302), .B2(n_1306), .B3(n_1307), .Y(n_1295) );
INVx2_ASAP7_75t_SL g1862 ( .A(n_565), .Y(n_1862) );
AND2x4_ASAP7_75t_L g1871 ( .A(n_566), .B(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
BUFx3_ASAP7_75t_L g1298 ( .A(n_570), .Y(n_1298) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g1305 ( .A(n_574), .Y(n_1305) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_575), .Y(n_971) );
BUFx2_ASAP7_75t_SL g1882 ( .A(n_575), .Y(n_1882) );
XNOR2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND3x1_ASAP7_75t_SL g578 ( .A(n_579), .B(n_599), .C(n_632), .Y(n_578) );
OAI31xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_587), .A3(n_595), .B(n_598), .Y(n_579) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g622 ( .A(n_583), .Y(n_622) );
INVx1_ASAP7_75t_L g831 ( .A(n_583), .Y(n_831) );
INVx1_ASAP7_75t_L g1106 ( .A(n_583), .Y(n_1106) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_583), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1890 ( .A(n_583), .B(n_1866), .Y(n_1890) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g625 ( .A(n_584), .B(n_585), .Y(n_625) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_589), .A2(n_657), .B(n_658), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_589), .A2(n_725), .B(n_726), .Y(n_724) );
HB1xp67_ASAP7_75t_L g1470 ( .A(n_590), .Y(n_1470) );
HB1xp67_ASAP7_75t_L g1924 ( .A(n_590), .Y(n_1924) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_591), .B(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g858 ( .A(n_591), .B(n_859), .Y(n_858) );
NAND4xp25_ASAP7_75t_SL g1218 ( .A(n_591), .B(n_1219), .C(n_1222), .D(n_1225), .Y(n_1218) );
NAND4xp25_ASAP7_75t_L g1314 ( .A(n_591), .B(n_1315), .C(n_1318), .D(n_1321), .Y(n_1314) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_598), .A2(n_652), .B(n_666), .C(n_679), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g715 ( .A1(n_598), .A2(n_716), .B(n_728), .C(n_741), .Y(n_715) );
OAI31xp33_ASAP7_75t_SL g802 ( .A1(n_598), .A2(n_803), .A3(n_804), .B(n_810), .Y(n_802) );
OAI31xp33_ASAP7_75t_L g855 ( .A1(n_598), .A2(n_856), .A3(n_857), .B(n_858), .Y(n_855) );
OAI31xp33_ASAP7_75t_SL g1159 ( .A1(n_598), .A2(n_1160), .A3(n_1161), .B(n_1163), .Y(n_1159) );
OAI31xp33_ASAP7_75t_L g1174 ( .A1(n_598), .A2(n_1175), .A3(n_1176), .B(n_1177), .Y(n_1174) );
AOI211xp5_ASAP7_75t_L g1415 ( .A1(n_598), .A2(n_1416), .B(n_1427), .C(n_1445), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_610), .B1(n_611), .B2(n_617), .C(n_618), .Y(n_599) );
INVx1_ASAP7_75t_L g910 ( .A(n_602), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_604), .A2(n_606), .B1(n_621), .B2(n_623), .C(n_626), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_605), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
OAI22xp33_ASAP7_75t_SL g612 ( .A1(n_607), .A2(n_613), .B1(n_614), .B2(n_616), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_607), .A2(n_845), .B1(n_853), .B2(n_854), .Y(n_852) );
INVx1_ASAP7_75t_L g1061 ( .A(n_607), .Y(n_1061) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_607), .Y(n_1117) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g783 ( .A(n_608), .Y(n_783) );
BUFx2_ASAP7_75t_L g815 ( .A(n_608), .Y(n_815) );
INVx2_ASAP7_75t_L g1836 ( .A(n_608), .Y(n_1836) );
AOI33xp33_ASAP7_75t_L g1288 ( .A1(n_610), .A2(n_617), .A3(n_1289), .B1(n_1291), .B2(n_1292), .B3(n_1293), .Y(n_1288) );
OAI22xp5_ASAP7_75t_SL g899 ( .A1(n_614), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI33xp33_ASAP7_75t_L g1009 ( .A1(n_617), .A2(n_1010), .A3(n_1011), .B1(n_1017), .B2(n_1024), .B3(n_1027), .Y(n_1009) );
INVx2_ASAP7_75t_L g1077 ( .A(n_617), .Y(n_1077) );
INVx1_ASAP7_75t_L g1158 ( .A(n_617), .Y(n_1158) );
AOI33xp33_ASAP7_75t_L g1928 ( .A1(n_617), .A2(n_1010), .A3(n_1929), .B1(n_1930), .B2(n_1933), .B3(n_1934), .Y(n_1928) );
OAI33xp33_ASAP7_75t_L g821 ( .A1(n_619), .A2(n_822), .A3(n_828), .B1(n_835), .B2(n_838), .B3(n_842), .Y(n_821) );
INVx1_ASAP7_75t_SL g1197 ( .A(n_619), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_621), .A2(n_623), .B1(n_628), .B2(n_629), .C(n_630), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_621), .A2(n_887), .B1(n_1089), .B2(n_1090), .C(n_1091), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_621), .A2(n_887), .B1(n_1126), .B2(n_1127), .C(n_1128), .Y(n_1125) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g788 ( .A(n_622), .Y(n_788) );
INVx2_ASAP7_75t_L g795 ( .A(n_622), .Y(n_795) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_623), .A2(n_795), .B1(n_900), .B2(n_901), .C(n_918), .Y(n_917) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_623), .A2(n_879), .B1(n_922), .B2(n_924), .C(n_925), .Y(n_921) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g888 ( .A(n_624), .Y(n_888) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g791 ( .A(n_625), .Y(n_791) );
BUFx2_ASAP7_75t_L g798 ( .A(n_625), .Y(n_798) );
BUFx4f_ASAP7_75t_L g834 ( .A(n_625), .Y(n_834) );
INVx1_ASAP7_75t_L g1052 ( .A(n_625), .Y(n_1052) );
INVx1_ASAP7_75t_L g827 ( .A(n_631), .Y(n_827) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_631), .Y(n_920) );
INVx1_ASAP7_75t_L g928 ( .A(n_631), .Y(n_928) );
INVx1_ASAP7_75t_L g1196 ( .A(n_631), .Y(n_1196) );
BUFx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x6_ASAP7_75t_L g1809 ( .A(n_636), .B(n_1806), .Y(n_1809) );
NAND2x1p5_ASAP7_75t_L g1829 ( .A(n_636), .B(n_1821), .Y(n_1829) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g1081 ( .A(n_642), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1842 ( .A(n_642), .Y(n_1842) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g773 ( .A(n_643), .Y(n_773) );
INVx1_ASAP7_75t_L g1144 ( .A(n_643), .Y(n_1144) );
INVx5_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_645), .A2(n_655), .B1(n_676), .B2(n_677), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_645), .A2(n_676), .B1(n_720), .B2(n_740), .Y(n_739) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_757), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_713), .B2(n_714), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g727 ( .A(n_660), .Y(n_727) );
AOI31xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_672), .A3(n_675), .B(n_678), .Y(n_666) );
AOI31xp33_ASAP7_75t_L g728 ( .A1(n_678), .A2(n_729), .A3(n_736), .B(n_739), .Y(n_728) );
AO21x1_ASAP7_75t_SL g1001 ( .A1(n_678), .A2(n_1002), .B(n_1006), .Y(n_1001) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_689), .C(n_697), .D(n_708), .Y(n_679) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g745 ( .A(n_685), .Y(n_745) );
INVx2_ASAP7_75t_SL g1431 ( .A(n_685), .Y(n_1431) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_686), .Y(n_907) );
BUFx2_ASAP7_75t_L g1436 ( .A(n_686), .Y(n_1436) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_694), .C(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g746 ( .A(n_695), .B(n_747), .C(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g785 ( .A(n_695), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g1432 ( .A(n_695), .B(n_1433), .C(n_1435), .Y(n_1432) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_702), .C(n_705), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g1129 ( .A(n_704), .Y(n_1129) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_705), .B(n_750), .C(n_753), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g1348 ( .A(n_705), .B(n_1349), .C(n_1351), .Y(n_1348) );
NAND3xp33_ASAP7_75t_L g1437 ( .A(n_705), .B(n_1438), .C(n_1439), .Y(n_1437) );
NAND3xp33_ASAP7_75t_L g1536 ( .A(n_705), .B(n_1537), .C(n_1541), .Y(n_1536) );
INVx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .C(n_712), .Y(n_708) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_710), .Y(n_1096) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_712), .B(n_755), .C(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g842 ( .A(n_712), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g1352 ( .A(n_712), .B(n_1353), .C(n_1354), .Y(n_1352) );
NAND3xp33_ASAP7_75t_L g1440 ( .A(n_712), .B(n_1441), .C(n_1442), .Y(n_1440) );
NAND3xp33_ASAP7_75t_L g1543 ( .A(n_712), .B(n_1544), .C(n_1545), .Y(n_1543) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g1347 ( .A(n_732), .Y(n_1347) );
INVx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_733), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1530 ( .A(n_733), .Y(n_1530) );
INVx1_ASAP7_75t_L g1120 ( .A(n_735), .Y(n_1120) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_742), .B(n_746), .C(n_749), .D(n_754), .Y(n_741) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_SL g975 ( .A(n_752), .Y(n_975) );
INVx1_ASAP7_75t_L g1857 ( .A(n_752), .Y(n_1857) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_818), .B1(n_868), .B2(n_869), .Y(n_757) );
INVx1_ASAP7_75t_L g868 ( .A(n_758), .Y(n_868) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_802), .C(n_811), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_786), .Y(n_760) );
OAI33xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .A3(n_770), .B1(n_777), .B2(n_781), .B3(n_785), .Y(n_761) );
OAI33xp33_ASAP7_75t_L g843 ( .A1(n_762), .A2(n_785), .A3(n_844), .B1(n_847), .B2(n_848), .B3(n_852), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_762), .A2(n_1079), .B1(n_1087), .B2(n_1088), .Y(n_1078) );
OAI33xp33_ASAP7_75t_L g1137 ( .A1(n_762), .A2(n_1138), .A3(n_1140), .B1(n_1148), .B2(n_1153), .B3(n_1158), .Y(n_1137) );
INVx1_ASAP7_75t_L g1379 ( .A(n_762), .Y(n_1379) );
OAI33xp33_ASAP7_75t_L g1830 ( .A1(n_762), .A2(n_915), .A3(n_1831), .B1(n_1837), .B2(n_1841), .B3(n_1847), .Y(n_1830) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_767), .B2(n_769), .Y(n_764) );
OAI22xp33_ASAP7_75t_SL g1073 ( .A1(n_765), .A2(n_1074), .B1(n_1075), .B2(n_1076), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g1138 ( .A1(n_765), .A2(n_1126), .B1(n_1127), .B2(n_1139), .Y(n_1138) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_766), .A2(n_769), .B1(n_788), .B2(n_789), .C(n_792), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_767), .A2(n_829), .B1(n_832), .B2(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g903 ( .A(n_767), .Y(n_903) );
BUFx3_ASAP7_75t_L g913 ( .A(n_767), .Y(n_913) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI22xp33_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_772), .B1(n_774), .B2(n_775), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_772), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g847 ( .A1(n_772), .A2(n_779), .B1(n_823), .B2(n_826), .Y(n_847) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g849 ( .A(n_773), .Y(n_849) );
INVx1_ASAP7_75t_L g1069 ( .A(n_773), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_773), .Y(n_1391) );
INVx1_ASAP7_75t_L g1384 ( .A(n_775), .Y(n_1384) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g1248 ( .A(n_776), .Y(n_1248) );
INVx2_ASAP7_75t_L g1396 ( .A(n_776), .Y(n_1396) );
INVx2_ASAP7_75t_L g1534 ( .A(n_776), .Y(n_1534) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_779), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g1153 ( .A1(n_783), .A2(n_1154), .B1(n_1156), .B2(n_1157), .Y(n_1153) );
OAI221xp5_ASAP7_75t_L g1363 ( .A1(n_789), .A2(n_1131), .B1(n_1364), .B2(n_1365), .C(n_1366), .Y(n_1363) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
BUFx2_ASAP7_75t_L g1133 ( .A(n_791), .Y(n_1133) );
BUFx3_ASAP7_75t_L g923 ( .A(n_793), .Y(n_923) );
BUFx2_ASAP7_75t_L g962 ( .A(n_793), .Y(n_962) );
INVx2_ASAP7_75t_L g1034 ( .A(n_793), .Y(n_1034) );
INVx1_ASAP7_75t_L g1376 ( .A(n_793), .Y(n_1376) );
OAI221xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .B1(n_797), .B2(n_799), .C(n_800), .Y(n_794) );
INVx2_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g1204 ( .A(n_801), .Y(n_1204) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g1035 ( .A(n_807), .Y(n_1035) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g1076 ( .A(n_815), .Y(n_1076) );
INVx1_ASAP7_75t_L g1139 ( .A(n_815), .Y(n_1139) );
INVx1_ASAP7_75t_L g869 ( .A(n_818), .Y(n_869) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_855), .C(n_863), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_843), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B1(n_826), .B2(n_827), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
BUFx4f_ASAP7_75t_L g1258 ( .A(n_825), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B1(n_832), .B2(n_833), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_830), .A2(n_833), .B1(n_836), .B2(n_837), .Y(n_835) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g1369 ( .A(n_840), .Y(n_1369) );
OAI22xp33_ASAP7_75t_L g1386 ( .A1(n_845), .A2(n_1364), .B1(n_1365), .B2(n_1387), .Y(n_1386) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_845), .A2(n_1389), .B1(n_1390), .B2(n_1392), .Y(n_1388) );
BUFx2_ASAP7_75t_L g1833 ( .A(n_845), .Y(n_1833) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_930), .B1(n_931), .B2(n_982), .Y(n_870) );
INVx1_ASAP7_75t_L g982 ( .A(n_871), .Y(n_982) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_895), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_890), .B(n_893), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OAI21xp33_ASAP7_75t_SL g1097 ( .A1(n_887), .A2(n_1098), .B(n_1099), .Y(n_1097) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
OAI31xp33_ASAP7_75t_L g1048 ( .A1(n_894), .A2(n_1049), .A3(n_1050), .B(n_1056), .Y(n_1048) );
AOI211x1_ASAP7_75t_SL g1460 ( .A1(n_894), .A2(n_1461), .B(n_1473), .C(n_1489), .Y(n_1460) );
AOI211xp5_ASAP7_75t_L g1502 ( .A1(n_894), .A2(n_1503), .B(n_1514), .C(n_1523), .Y(n_1502) );
AOI211xp5_ASAP7_75t_SL g1914 ( .A1(n_894), .A2(n_1915), .B(n_1927), .C(n_1941), .Y(n_1914) );
OAI22xp33_ASAP7_75t_L g1847 ( .A1(n_902), .A2(n_1833), .B1(n_1848), .B2(n_1849), .Y(n_1847) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_907), .Y(n_1290) );
OAI22xp33_ASAP7_75t_SL g908 ( .A1(n_909), .A2(n_910), .B1(n_911), .B2(n_912), .Y(n_908) );
BUFx3_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OAI33xp33_ASAP7_75t_L g1377 ( .A1(n_915), .A2(n_1378), .A3(n_1380), .B1(n_1386), .B2(n_1388), .B3(n_1393), .Y(n_1377) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_SL g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g981 ( .A(n_933), .Y(n_981) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g1481 ( .A(n_941), .Y(n_1481) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
NAND4xp25_ASAP7_75t_SL g948 ( .A(n_949), .B(n_950), .C(n_952), .D(n_954), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_976), .Y(n_958) );
AOI33xp33_ASAP7_75t_L g1031 ( .A1(n_960), .A2(n_1032), .A3(n_1036), .B1(n_1040), .B2(n_1042), .B3(n_1044), .Y(n_1031) );
NAND3xp33_ASAP7_75t_L g1250 ( .A(n_960), .B(n_1251), .C(n_1254), .Y(n_1250) );
INVx2_ASAP7_75t_SL g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g1547 ( .A(n_964), .Y(n_1547) );
INVx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
BUFx2_ASAP7_75t_L g1136 ( .A(n_965), .Y(n_1136) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g1488 ( .A(n_966), .Y(n_1488) );
OR2x2_ASAP7_75t_L g1892 ( .A(n_966), .B(n_1866), .Y(n_1892) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g1304 ( .A(n_970), .Y(n_1304) );
BUFx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_984), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B1(n_1111), .B2(n_1166), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_1045), .B1(n_1109), .B2(n_1110), .Y(n_986) );
INVx1_ASAP7_75t_L g1110 ( .A(n_987), .Y(n_1110) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
NAND4xp25_ASAP7_75t_L g989 ( .A(n_990), .B(n_1001), .C(n_1009), .D(n_1031), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_997), .Y(n_991) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_1010), .Y(n_1187) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_1014), .Y(n_1244) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1014), .Y(n_1346) );
AND2x4_ASAP7_75t_L g1812 ( .A(n_1014), .B(n_1806), .Y(n_1812) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1023), .Y(n_1343) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1026), .Y(n_1242) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1028), .Y(n_1152) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1029), .Y(n_1072) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1029), .Y(n_1084) );
INVx3_ASAP7_75t_L g1147 ( .A(n_1029), .Y(n_1147) );
INVx2_ASAP7_75t_SL g1434 ( .A(n_1029), .Y(n_1434) );
INVx2_ASAP7_75t_L g1845 ( .A(n_1029), .Y(n_1845) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx4_ASAP7_75t_L g1041 ( .A(n_1038), .Y(n_1041) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1038), .Y(n_1350) );
CKINVDCx5p33_ASAP7_75t_R g1087 ( .A(n_1044), .Y(n_1087) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_1044), .B(n_1256), .C(n_1257), .Y(n_1255) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1045), .Y(n_1109) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1047), .Y(n_1107) );
NAND3xp33_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1057), .C(n_1064), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1061), .Y(n_1387) );
NOR3xp33_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1078), .C(n_1095), .Y(n_1064) );
NOR3xp33_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1073), .C(n_1077), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1068), .B1(n_1070), .B2(n_1071), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_1076), .A2(n_1394), .B1(n_1397), .B2(n_1398), .Y(n_1393) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1082), .B1(n_1083), .B2(n_1085), .C(n_1086), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1094), .Y(n_1542) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx2_ASAP7_75t_L g1873 ( .A(n_1102), .Y(n_1873) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx2_ASAP7_75t_L g1876 ( .A(n_1104), .Y(n_1876) );
BUFx2_ASAP7_75t_L g1371 ( .A(n_1105), .Y(n_1371) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1111), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1113), .Y(n_1164) );
NAND3xp33_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1123), .C(n_1159), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1137), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1132), .B1(n_1133), .B2(n_1134), .C(n_1135), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1142), .B1(n_1145), .B2(n_1146), .Y(n_1140) );
INVx2_ASAP7_75t_SL g1142 ( .A(n_1143), .Y(n_1142) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1143), .Y(n_1150) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1143), .Y(n_1382) );
INVx2_ASAP7_75t_L g1839 ( .A(n_1143), .Y(n_1839) );
BUFx3_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
OAI22xp5_ASAP7_75t_SL g1148 ( .A1(n_1149), .A2(n_1150), .B1(n_1151), .B2(n_1152), .Y(n_1148) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
OAI22xp33_ASAP7_75t_L g1611 ( .A1(n_1165), .A2(n_1590), .B1(n_1612), .B2(n_1613), .Y(n_1611) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1170), .B1(n_1355), .B2(n_1356), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
XNOR2xp5_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1261), .Y(n_1170) );
XOR2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1216), .Y(n_1171) );
NAND3x1_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1181), .C(n_1207), .Y(n_1173) );
AND4x1_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1188), .C(n_1191), .D(n_1198), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1186), .C(n_1187), .Y(n_1182) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
NAND3xp33_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1194), .C(n_1197), .Y(n_1191) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
NAND3xp33_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1202), .C(n_1206), .Y(n_1198) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1937 ( .A(n_1204), .Y(n_1937) );
AOI33xp33_ASAP7_75t_L g1482 ( .A1(n_1206), .A2(n_1296), .A3(n_1483), .B1(n_1485), .B2(n_1486), .B3(n_1487), .Y(n_1482) );
AOI33xp33_ASAP7_75t_L g1935 ( .A1(n_1206), .A2(n_1296), .A3(n_1936), .B1(n_1938), .B2(n_1939), .B3(n_1940), .Y(n_1935) );
NAND4xp25_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1245), .C(n_1250), .D(n_1255), .Y(n_1239) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx2_ASAP7_75t_SL g1526 ( .A(n_1248), .Y(n_1526) );
BUFx6f_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1253), .Y(n_1859) );
AND2x4_ASAP7_75t_L g1886 ( .A(n_1253), .B(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1263), .B1(n_1311), .B2(n_1312), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1265), .Y(n_1310) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1295), .Y(n_1287) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_1300), .A2(n_1371), .B1(n_1372), .B2(n_1373), .C(n_1374), .Y(n_1370) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
NAND3xp33_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1330), .C(n_1333), .Y(n_1325) );
NAND4xp25_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1339), .C(n_1348), .D(n_1352), .Y(n_1335) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
XNOR2xp5_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1456), .Y(n_1356) );
AOI22xp5_ASAP7_75t_L g1357 ( .A1(n_1358), .A2(n_1411), .B1(n_1454), .B2(n_1455), .Y(n_1357) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1358), .Y(n_1454) );
HB1xp67_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
NAND3xp33_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1399), .C(n_1406), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1377), .Y(n_1361) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1368), .Y(n_1881) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1382), .B1(n_1383), .B2(n_1385), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1837 ( .A1(n_1383), .A2(n_1838), .B1(n_1839), .B2(n_1840), .Y(n_1837) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVx2_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1411), .Y(n_1455) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
NAND4xp25_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1432), .C(n_1437), .D(n_1440), .Y(n_1427) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
HB1xp67_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1499), .B1(n_1500), .B2(n_1549), .Y(n_1457) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1458), .Y(n_1549) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1460), .Y(n_1498) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1482), .Y(n_1473) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1502), .Y(n_1548) );
NAND4xp25_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1531), .C(n_1536), .D(n_1543), .Y(n_1523) );
BUFx2_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx2_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx2_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
OAI221xp5_ASAP7_75t_L g1551 ( .A1(n_1552), .A2(n_1795), .B1(n_1797), .B2(n_1900), .C(n_1906), .Y(n_1551) );
AOI21xp5_ASAP7_75t_L g1552 ( .A1(n_1553), .A2(n_1716), .B(n_1761), .Y(n_1552) );
NAND3xp33_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1634), .C(n_1655), .Y(n_1553) );
O2A1O1Ixp33_ASAP7_75t_L g1554 ( .A1(n_1555), .A2(n_1603), .B(n_1617), .C(n_1619), .Y(n_1554) );
O2A1O1Ixp33_ASAP7_75t_L g1634 ( .A1(n_1555), .A2(n_1635), .B(n_1638), .C(n_1640), .Y(n_1634) );
NOR2xp33_ASAP7_75t_SL g1555 ( .A(n_1556), .B(n_1599), .Y(n_1555) );
NOR2xp33_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1577), .Y(n_1556) );
OAI21xp33_ASAP7_75t_L g1635 ( .A1(n_1557), .A2(n_1604), .B(n_1636), .Y(n_1635) );
INVx3_ASAP7_75t_L g1644 ( .A(n_1557), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1557), .B(n_1637), .Y(n_1740) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1557), .B(n_1672), .Y(n_1774) );
CKINVDCx5p33_ASAP7_75t_R g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1558), .Y(n_1618) );
INVx1_ASAP7_75t_SL g1628 ( .A(n_1558), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1558), .B(n_1626), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1558), .B(n_1637), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1558), .B(n_1599), .Y(n_1683) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1558), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1558), .B(n_1579), .Y(n_1746) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1558), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1567), .Y(n_1558) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1560), .Y(n_1709) );
BUFx3_ASAP7_75t_L g1796 ( .A(n_1560), .Y(n_1796) );
AND2x4_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1564), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1561), .B(n_1564), .Y(n_1601) );
HB1xp67_ASAP7_75t_L g1954 ( .A(n_1561), .Y(n_1954) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
AND2x4_ASAP7_75t_L g1566 ( .A(n_1562), .B(n_1564), .Y(n_1566) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1563), .B(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1565), .Y(n_1571) );
INVx2_ASAP7_75t_L g1610 ( .A(n_1566), .Y(n_1610) );
AND2x4_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1572), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
OR2x2_ASAP7_75t_L g1591 ( .A(n_1570), .B(n_1573), .Y(n_1591) );
HB1xp67_ASAP7_75t_L g1953 ( .A(n_1571), .Y(n_1953) );
AND2x4_ASAP7_75t_L g1574 ( .A(n_1572), .B(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1573), .B(n_1576), .Y(n_1593) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1577), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1586), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1782 ( .A(n_1578), .B(n_1615), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1582), .Y(n_1578) );
INVx4_ASAP7_75t_L g1626 ( .A(n_1579), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1579), .B(n_1586), .Y(n_1639) );
INVx3_ASAP7_75t_L g1653 ( .A(n_1579), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1579), .B(n_1615), .Y(n_1695) );
NOR2xp33_ASAP7_75t_L g1704 ( .A(n_1579), .B(n_1648), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1579), .B(n_1627), .Y(n_1725) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1579), .B(n_1659), .Y(n_1757) );
AND2x4_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1581), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1582), .B(n_1664), .Y(n_1663) );
OR2x2_ASAP7_75t_L g1666 ( .A(n_1582), .B(n_1667), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1582), .B(n_1594), .Y(n_1687) );
OAI322xp33_ASAP7_75t_L g1723 ( .A1(n_1582), .A2(n_1645), .A3(n_1695), .B1(n_1724), .B2(n_1726), .C1(n_1727), .C2(n_1730), .Y(n_1723) );
NOR2xp33_ASAP7_75t_L g1736 ( .A(n_1582), .B(n_1594), .Y(n_1736) );
OR2x2_ASAP7_75t_L g1764 ( .A(n_1582), .B(n_1639), .Y(n_1764) );
OR2x2_ASAP7_75t_L g1772 ( .A(n_1582), .B(n_1631), .Y(n_1772) );
BUFx3_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1583), .B(n_1615), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1583), .B(n_1586), .Y(n_1621) );
INVx2_ASAP7_75t_L g1632 ( .A(n_1583), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1583), .B(n_1659), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1583), .B(n_1649), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1583), .B(n_1631), .Y(n_1731) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1583), .B(n_1698), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1585), .Y(n_1583) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1586), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1586), .B(n_1679), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1750 ( .A(n_1586), .B(n_1653), .Y(n_1750) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1594), .Y(n_1586) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1587), .Y(n_1616) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1587), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1587), .B(n_1595), .Y(n_1649) );
OAI22xp33_ASAP7_75t_L g1588 ( .A1(n_1589), .A2(n_1590), .B1(n_1592), .B2(n_1593), .Y(n_1588) );
OAI22xp5_ASAP7_75t_L g1596 ( .A1(n_1590), .A2(n_1593), .B1(n_1597), .B2(n_1598), .Y(n_1596) );
BUFx3_ASAP7_75t_L g1712 ( .A(n_1590), .Y(n_1712) );
BUFx6f_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
HB1xp67_ASAP7_75t_L g1613 ( .A(n_1593), .Y(n_1613) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1593), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1594), .B(n_1616), .Y(n_1659) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1594), .Y(n_1664) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1595), .B(n_1616), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1599), .B(n_1607), .Y(n_1606) );
CKINVDCx5p33_ASAP7_75t_R g1622 ( .A(n_1599), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1599), .B(n_1628), .Y(n_1627) );
CKINVDCx6p67_ASAP7_75t_R g1637 ( .A(n_1599), .Y(n_1637) );
OR2x6_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1602), .Y(n_1599) );
INVxp67_ASAP7_75t_SL g1603 ( .A(n_1604), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1614), .Y(n_1604) );
OAI221xp5_ASAP7_75t_L g1701 ( .A1(n_1605), .A2(n_1644), .B1(n_1702), .B2(n_1703), .C(n_1705), .Y(n_1701) );
INVx2_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1606), .B(n_1729), .Y(n_1728) );
AOI221xp5_ASAP7_75t_L g1732 ( .A1(n_1606), .A2(n_1665), .B1(n_1733), .B2(n_1735), .C(n_1737), .Y(n_1732) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1607), .B(n_1637), .Y(n_1636) );
AND2x4_ASAP7_75t_SL g1672 ( .A(n_1607), .B(n_1637), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1607), .B(n_1644), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1756 ( .A(n_1607), .B(n_1626), .Y(n_1756) );
INVx2_ASAP7_75t_SL g1607 ( .A(n_1608), .Y(n_1607) );
INVx2_ASAP7_75t_L g1633 ( .A(n_1608), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1608), .B(n_1637), .Y(n_1647) );
OR2x2_ASAP7_75t_L g1726 ( .A(n_1608), .B(n_1644), .Y(n_1726) );
INVx2_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1614), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1615), .B(n_1626), .Y(n_1642) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1615), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1615), .B(n_1679), .Y(n_1718) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
O2A1O1Ixp33_ASAP7_75t_L g1619 ( .A1(n_1620), .A2(n_1622), .B(n_1623), .C(n_1633), .Y(n_1619) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1621), .B(n_1683), .Y(n_1794) );
AOI21xp33_ASAP7_75t_L g1747 ( .A1(n_1622), .A2(n_1748), .B(n_1751), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1624), .B(n_1629), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1624), .B(n_1662), .Y(n_1688) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
NOR2xp33_ASAP7_75t_L g1697 ( .A(n_1625), .B(n_1698), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1627), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1626), .B(n_1632), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1626), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1626), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1627), .B(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1627), .Y(n_1742) );
NAND2xp5_ASAP7_75t_L g1646 ( .A(n_1628), .B(n_1647), .Y(n_1646) );
NAND3xp33_ASAP7_75t_L g1744 ( .A(n_1629), .B(n_1637), .C(n_1745), .Y(n_1744) );
AOI322xp5_ASAP7_75t_L g1785 ( .A1(n_1629), .A2(n_1647), .A3(n_1733), .B1(n_1745), .B2(n_1786), .C1(n_1788), .C2(n_1790), .Y(n_1785) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1632), .Y(n_1630) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1632), .B(n_1649), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1632), .B(n_1659), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1632), .B(n_1694), .Y(n_1693) );
OR2x2_ASAP7_75t_L g1749 ( .A(n_1632), .B(n_1750), .Y(n_1749) );
OAI321xp33_ASAP7_75t_L g1751 ( .A1(n_1632), .A2(n_1643), .A3(n_1706), .B1(n_1752), .B2(n_1755), .C(n_1757), .Y(n_1751) );
INVx2_ASAP7_75t_L g1645 ( .A(n_1633), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1633), .B(n_1683), .Y(n_1691) );
NAND3xp33_ASAP7_75t_L g1700 ( .A(n_1633), .B(n_1654), .C(n_1674), .Y(n_1700) );
INVx2_ASAP7_75t_L g1734 ( .A(n_1633), .Y(n_1734) );
AOI221xp5_ASAP7_75t_L g1775 ( .A1(n_1633), .A2(n_1676), .B1(n_1776), .B2(n_1777), .C(n_1783), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1637), .B(n_1780), .Y(n_1779) );
A2O1A1Ixp33_ASAP7_75t_L g1767 ( .A1(n_1638), .A2(n_1672), .B(n_1718), .C(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
OAI221xp5_ASAP7_75t_L g1640 ( .A1(n_1641), .A2(n_1643), .B1(n_1646), .B2(n_1648), .C(n_1650), .Y(n_1640) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
NAND2xp5_ASAP7_75t_L g1643 ( .A(n_1644), .B(n_1645), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1781 ( .A(n_1644), .B(n_1782), .Y(n_1781) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1645), .B(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1646), .Y(n_1790) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1647), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1668 ( .A(n_1647), .B(n_1653), .Y(n_1668) );
AOI32xp33_ASAP7_75t_L g1758 ( .A1(n_1647), .A2(n_1654), .A3(n_1674), .B1(n_1683), .B2(n_1759), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_1648), .B(n_1754), .Y(n_1753) );
OAI21xp33_ASAP7_75t_L g1788 ( .A1(n_1648), .A2(n_1653), .B(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
INVxp67_ASAP7_75t_SL g1765 ( .A(n_1650), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1654), .Y(n_1651) );
INVx2_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
OR2x2_ASAP7_75t_L g1657 ( .A(n_1653), .B(n_1658), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1653), .B(n_1720), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1653), .B(n_1736), .Y(n_1735) );
O2A1O1Ixp33_ASAP7_75t_SL g1783 ( .A1(n_1653), .A2(n_1690), .B(n_1703), .C(n_1784), .Y(n_1783) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1654), .Y(n_1686) );
NOR5xp2_ASAP7_75t_L g1655 ( .A(n_1656), .B(n_1680), .C(n_1689), .D(n_1699), .E(n_1701), .Y(n_1655) );
OAI221xp5_ASAP7_75t_L g1656 ( .A1(n_1657), .A2(n_1660), .B1(n_1661), .B2(n_1668), .C(n_1669), .Y(n_1656) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1657), .Y(n_1776) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1659), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1659), .B(n_1679), .Y(n_1760) );
NOR2xp33_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1665), .Y(n_1661) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
OAI21xp33_ASAP7_75t_L g1777 ( .A1(n_1663), .A2(n_1778), .B(n_1781), .Y(n_1777) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
AOI22xp33_ASAP7_75t_SL g1669 ( .A1(n_1670), .A2(n_1675), .B1(n_1676), .B2(n_1677), .Y(n_1669) );
NAND2xp33_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1673), .Y(n_1670) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1675), .Y(n_1784) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
OAI211xp5_ASAP7_75t_L g1770 ( .A1(n_1679), .A2(n_1771), .B(n_1772), .C(n_1773), .Y(n_1770) );
OAI21xp5_ASAP7_75t_L g1680 ( .A1(n_1681), .A2(n_1684), .B(n_1688), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
AOI221xp5_ASAP7_75t_L g1762 ( .A1(n_1683), .A2(n_1728), .B1(n_1763), .B2(n_1765), .C(n_1766), .Y(n_1762) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
NAND2xp5_ASAP7_75t_SL g1685 ( .A(n_1686), .B(n_1687), .Y(n_1685) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1687), .Y(n_1792) );
OAI21xp5_ASAP7_75t_L g1689 ( .A1(n_1690), .A2(n_1692), .B(n_1696), .Y(n_1689) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
NOR2xp33_ASAP7_75t_L g1741 ( .A(n_1695), .B(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVxp67_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVx2_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
BUFx3_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
OAI22xp33_ASAP7_75t_L g1710 ( .A1(n_1711), .A2(n_1712), .B1(n_1713), .B2(n_1714), .Y(n_1710) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
NAND5xp2_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1732), .C(n_1739), .D(n_1747), .E(n_1758), .Y(n_1716) );
O2A1O1Ixp33_ASAP7_75t_L g1717 ( .A1(n_1718), .A2(n_1719), .B(n_1721), .C(n_1723), .Y(n_1717) );
AOI211xp5_ASAP7_75t_L g1739 ( .A1(n_1718), .A2(n_1740), .B(n_1741), .C(n_1743), .Y(n_1739) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1720), .Y(n_1789) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
A2O1A1Ixp33_ASAP7_75t_L g1791 ( .A1(n_1725), .A2(n_1734), .B(n_1792), .C(n_1793), .Y(n_1791) );
NOR2xp33_ASAP7_75t_L g1737 ( .A(n_1726), .B(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1750), .Y(n_1771) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
NAND4xp25_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1775), .C(n_1785), .D(n_1791), .Y(n_1761) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
NAND2xp5_ASAP7_75t_SL g1766 ( .A(n_1767), .B(n_1770), .Y(n_1766) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
INVxp33_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
INVxp67_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
HB1xp67_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
NAND2xp5_ASAP7_75t_L g1799 ( .A(n_1800), .B(n_1850), .Y(n_1799) );
NOR3xp33_ASAP7_75t_L g1800 ( .A(n_1801), .B(n_1815), .C(n_1830), .Y(n_1800) );
NAND2xp5_ASAP7_75t_L g1801 ( .A(n_1802), .B(n_1810), .Y(n_1801) );
AOI22xp33_ASAP7_75t_L g1802 ( .A1(n_1803), .A2(n_1804), .B1(n_1808), .B2(n_1809), .Y(n_1802) );
BUFx2_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
AOI22xp33_ASAP7_75t_L g1810 ( .A1(n_1811), .A2(n_1812), .B1(n_1813), .B2(n_1814), .Y(n_1810) );
INVx2_ASAP7_75t_SL g1816 ( .A(n_1817), .Y(n_1816) );
INVx2_ASAP7_75t_L g1817 ( .A(n_1818), .Y(n_1817) );
NAND2x1_ASAP7_75t_SL g1818 ( .A(n_1819), .B(n_1821), .Y(n_1818) );
INVx2_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
NAND2x1p5_ASAP7_75t_L g1825 ( .A(n_1821), .B(n_1826), .Y(n_1825) );
INVx3_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
BUFx4f_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
BUFx2_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
OAI22xp33_ASAP7_75t_L g1831 ( .A1(n_1832), .A2(n_1833), .B1(n_1834), .B2(n_1835), .Y(n_1831) );
HB1xp67_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
OAI22xp5_ASAP7_75t_L g1841 ( .A1(n_1842), .A2(n_1843), .B1(n_1844), .B2(n_1846), .Y(n_1841) );
AOI221xp5_ASAP7_75t_L g1855 ( .A1(n_1843), .A2(n_1856), .B1(n_1863), .B2(n_1864), .C(n_1868), .Y(n_1855) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
AOI22xp33_ASAP7_75t_L g1888 ( .A1(n_1846), .A2(n_1848), .B1(n_1889), .B2(n_1891), .Y(n_1888) );
AOI221xp5_ASAP7_75t_L g1877 ( .A1(n_1849), .A2(n_1878), .B1(n_1880), .B2(n_1884), .C(n_1886), .Y(n_1877) );
AOI22xp33_ASAP7_75t_L g1850 ( .A1(n_1851), .A2(n_1854), .B1(n_1893), .B2(n_1894), .Y(n_1850) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx2_ASAP7_75t_L g1852 ( .A(n_1853), .Y(n_1852) );
NAND3xp33_ASAP7_75t_L g1854 ( .A(n_1855), .B(n_1877), .C(n_1888), .Y(n_1854) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
INVx2_ASAP7_75t_L g1865 ( .A(n_1866), .Y(n_1865) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1867), .Y(n_1872) );
INVx2_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
AND2x4_ASAP7_75t_L g1870 ( .A(n_1871), .B(n_1873), .Y(n_1870) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1871), .Y(n_1875) );
OR2x2_ASAP7_75t_L g1874 ( .A(n_1875), .B(n_1876), .Y(n_1874) );
INVx1_ASAP7_75t_SL g1887 ( .A(n_1875), .Y(n_1887) );
BUFx6f_ASAP7_75t_L g1878 ( .A(n_1879), .Y(n_1878) );
INVx6_ASAP7_75t_L g1889 ( .A(n_1890), .Y(n_1889) );
INVx4_ASAP7_75t_L g1891 ( .A(n_1892), .Y(n_1891) );
INVx5_ASAP7_75t_L g1894 ( .A(n_1895), .Y(n_1894) );
AND2x4_ASAP7_75t_L g1895 ( .A(n_1896), .B(n_1897), .Y(n_1895) );
INVx2_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
INVx1_ASAP7_75t_SL g1900 ( .A(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g1901 ( .A(n_1902), .Y(n_1901) );
INVx1_ASAP7_75t_L g1902 ( .A(n_1903), .Y(n_1902) );
INVx1_ASAP7_75t_L g1903 ( .A(n_1904), .Y(n_1903) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
CKINVDCx5p33_ASAP7_75t_R g1908 ( .A(n_1909), .Y(n_1908) );
A2O1A1Ixp33_ASAP7_75t_L g1951 ( .A1(n_1910), .A2(n_1952), .B(n_1954), .C(n_1955), .Y(n_1951) );
INVxp33_ASAP7_75t_SL g1911 ( .A(n_1912), .Y(n_1911) );
HB1xp67_ASAP7_75t_L g1913 ( .A(n_1914), .Y(n_1913) );
NAND2xp5_ASAP7_75t_L g1927 ( .A(n_1928), .B(n_1935), .Y(n_1927) );
INVx1_ASAP7_75t_L g1931 ( .A(n_1932), .Y(n_1931) );
HB1xp67_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
INVx1_ASAP7_75t_L g1952 ( .A(n_1953), .Y(n_1952) );
endmodule