module real_jpeg_20424_n_5 (n_17, n_4, n_0, n_18, n_1, n_2, n_16, n_3, n_5);

input n_17;
input n_4;
input n_0;
input n_18;
input n_1;
input n_2;
input n_16;
input n_3;

output n_5;

wire n_8;
wire n_11;
wire n_14;
wire n_7;
wire n_10;
wire n_9;
wire n_12;
wire n_6;
wire n_13;

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_17),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_18),
.Y(n_12)
);

AOI221xp5_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.C(n_13),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_L g5 ( 
.A1(n_2),
.A2(n_6),
.B1(n_7),
.B2(n_14),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_16),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_11),
.B(n_12),
.Y(n_9)
);


endmodule