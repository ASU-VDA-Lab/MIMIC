module fake_jpeg_9169_n_272 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_26),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_37),
.B(n_38),
.C(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_45),
.B1(n_24),
.B2(n_19),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_24),
.B1(n_18),
.B2(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_18),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_67),
.Y(n_85)
);

AOI22x1_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_63),
.Y(n_92)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_71),
.B1(n_35),
.B2(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_29),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_53),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_73),
.B1(n_19),
.B2(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_42),
.B1(n_53),
.B2(n_44),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_42),
.Y(n_82)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_39),
.Y(n_90)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_71),
.B1(n_65),
.B2(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_38),
.B1(n_52),
.B2(n_36),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_83),
.B1(n_87),
.B2(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_89),
.B1(n_59),
.B2(n_67),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_54),
.B(n_25),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_35),
.B1(n_32),
.B2(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_94),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_26),
.B(n_33),
.C(n_55),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_73),
.B1(n_66),
.B2(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_101),
.B1(n_108),
.B2(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_71),
.B1(n_32),
.B2(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_60),
.C(n_74),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_90),
.C(n_93),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_80),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_20),
.B(n_22),
.Y(n_125)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_68),
.B(n_25),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_94),
.B(n_85),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_128),
.C(n_30),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_86),
.B(n_85),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_131),
.B(n_114),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_125),
.B(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_83),
.B1(n_75),
.B2(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_75),
.B1(n_17),
.B2(n_30),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_100),
.C(n_102),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_33),
.B(n_54),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_34),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_138),
.B(n_147),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_112),
.B(n_114),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_109),
.C(n_99),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_116),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_112),
.B1(n_98),
.B2(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_20),
.B1(n_28),
.B2(n_16),
.Y(n_180)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_150),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_113),
.B1(n_34),
.B2(n_31),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_117),
.B1(n_135),
.B2(n_133),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_33),
.B1(n_34),
.B2(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_155),
.B1(n_156),
.B2(n_121),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_33),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_34),
.B(n_31),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_121),
.B(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_152),
.C(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_173),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_171),
.C(n_172),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_165),
.B1(n_169),
.B2(n_23),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_144),
.B1(n_158),
.B2(n_154),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_167),
.B(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_134),
.B1(n_123),
.B2(n_128),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_125),
.B(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_138),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_115),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_117),
.C(n_126),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_22),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_23),
.C(n_20),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_176),
.C(n_145),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_22),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_0),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_187),
.B(n_175),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_192),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_151),
.C(n_139),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_191),
.C(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_197),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_141),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_198),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_141),
.C(n_156),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_155),
.B1(n_16),
.B2(n_23),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_166),
.B(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_20),
.C(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_20),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_7),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_165),
.B1(n_160),
.B2(n_161),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_215),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_216),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_179),
.B(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_185),
.B1(n_198),
.B2(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_176),
.C(n_20),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_0),
.C(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_7),
.C(n_11),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_228),
.C(n_209),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_6),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_5),
.C(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_5),
.C(n_10),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_204),
.C(n_210),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_13),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_212),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_237),
.C(n_219),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_10),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_211),
.B(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_212),
.C(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_9),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_9),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_242),
.B(n_10),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_230),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_247),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_221),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_249),
.B(n_251),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_243),
.A2(n_1),
.B(n_2),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_252),
.A2(n_2),
.B(n_3),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_236),
.C(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_254),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_244),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_248),
.B(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_2),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_2),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_259),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_3),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_264),
.B(n_266),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_261),
.C(n_247),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_245),
.B(n_4),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_4),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_4),
.Y(n_272)
);


endmodule