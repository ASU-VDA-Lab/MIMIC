module fake_jpeg_29983_n_454 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_454);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_454;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_48),
.B(n_72),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_49),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_2),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_2),
.C(n_3),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_75),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_37),
.A2(n_2),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_4),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_35),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_19),
.B1(n_43),
.B2(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_83),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_6),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_49),
.B(n_27),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_113),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_44),
.B(n_28),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_110),
.B(n_93),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_126),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_130),
.B1(n_131),
.B2(n_80),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_46),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_129),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_51),
.A2(n_28),
.B1(n_44),
.B2(n_43),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_50),
.A2(n_28),
.B1(n_43),
.B2(n_19),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_26),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_68),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_45),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_46),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_62),
.B(n_20),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_20),
.Y(n_189)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_96),
.A2(n_40),
.B1(n_39),
.B2(n_86),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_157),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_108),
.A2(n_53),
.B1(n_92),
.B2(n_90),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_177),
.B1(n_181),
.B2(n_199),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_40),
.B1(n_28),
.B2(n_19),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_159),
.A2(n_168),
.B1(n_192),
.B2(n_197),
.Y(n_218)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_167),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_97),
.A2(n_40),
.B1(n_32),
.B2(n_30),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_193),
.B1(n_100),
.B2(n_135),
.Y(n_208)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_176),
.Y(n_209)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_122),
.A2(n_141),
.B1(n_137),
.B2(n_139),
.Y(n_177)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_114),
.A2(n_84),
.B1(n_82),
.B2(n_79),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_132),
.B(n_74),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_184),
.C(n_187),
.Y(n_224)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_189),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_98),
.B(n_69),
.C(n_67),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_196),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_99),
.B(n_66),
.C(n_63),
.Y(n_187)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_97),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_106),
.A2(n_55),
.B1(n_60),
.B2(n_29),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

BUFx4f_ASAP7_75t_SL g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_195),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_135),
.A2(n_33),
.B1(n_8),
.B2(n_9),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_198),
.A2(n_201),
.B1(n_8),
.B2(n_9),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_114),
.A2(n_33),
.B1(n_8),
.B2(n_9),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_11),
.Y(n_245)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_116),
.B(n_7),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_7),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_208),
.A2(n_215),
.B1(n_227),
.B2(n_185),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_100),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_209),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_106),
.B1(n_147),
.B2(n_111),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_147),
.B1(n_111),
.B2(n_120),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_200),
.B1(n_197),
.B2(n_194),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_172),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_149),
.B1(n_116),
.B2(n_134),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_225),
.A2(n_237),
.B1(n_212),
.B2(n_238),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_134),
.B1(n_102),
.B2(n_129),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_102),
.B1(n_144),
.B2(n_33),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_199),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_182),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_153),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_170),
.A2(n_10),
.B(n_11),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_241),
.A2(n_244),
.B(n_12),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_187),
.A2(n_10),
.B(n_11),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_247),
.B(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_184),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_251),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_178),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_162),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_256),
.Y(n_301)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_255),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_179),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_150),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_268),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_267),
.B1(n_215),
.B2(n_278),
.Y(n_288)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_SL g261 ( 
.A(n_222),
.B(n_185),
.C(n_181),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_262),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_265),
.B1(n_242),
.B2(n_223),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_206),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_208),
.A2(n_155),
.B1(n_171),
.B2(n_175),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_213),
.A2(n_173),
.B1(n_191),
.B2(n_190),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_267),
.A2(n_278),
.B1(n_280),
.B2(n_212),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_183),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_273),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_270),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_276),
.B1(n_207),
.B2(n_204),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_209),
.B(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_221),
.B(n_166),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_213),
.A2(n_151),
.B1(n_160),
.B2(n_165),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_241),
.B(n_11),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_282),
.B(n_245),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_203),
.A2(n_167),
.B1(n_154),
.B2(n_180),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_180),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_283),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_240),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_203),
.B(n_210),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_284),
.A2(n_292),
.B(n_316),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_244),
.C(n_232),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_287),
.C(n_304),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_240),
.C(n_220),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_288),
.A2(n_299),
.B1(n_249),
.B2(n_253),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_255),
.A2(n_218),
.B1(n_216),
.B2(n_240),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g293 ( 
.A1(n_255),
.A2(n_220),
.B1(n_223),
.B2(n_236),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_274),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_296),
.A2(n_303),
.B1(n_313),
.B2(n_314),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g344 ( 
.A1(n_300),
.A2(n_302),
.B(n_231),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_271),
.A2(n_217),
.B1(n_236),
.B2(n_233),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_228),
.C(n_219),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_282),
.A2(n_245),
.B(n_207),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_258),
.B(n_280),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_217),
.B1(n_228),
.B2(n_219),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_259),
.A2(n_238),
.B1(n_235),
.B2(n_229),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_247),
.B(n_235),
.C(n_229),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_258),
.C(n_266),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_269),
.B(n_273),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_319),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_340),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_254),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_325),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_257),
.Y(n_323)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_277),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_329),
.C(n_332),
.Y(n_349)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_246),
.C(n_262),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_297),
.Y(n_330)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_287),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_334),
.A2(n_303),
.B1(n_299),
.B2(n_317),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_292),
.A2(n_270),
.B1(n_260),
.B2(n_231),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_335),
.A2(n_343),
.B1(n_344),
.B2(n_324),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_270),
.Y(n_336)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_231),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_338),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_295),
.B(n_293),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_342),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_231),
.Y(n_342)
);

AOI22x1_ASAP7_75t_L g343 ( 
.A1(n_291),
.A2(n_290),
.B1(n_295),
.B2(n_288),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_12),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_304),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_318),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_284),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_351),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_291),
.B1(n_290),
.B2(n_296),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_356),
.A2(n_362),
.B1(n_335),
.B2(n_333),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_315),
.C(n_312),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_358),
.C(n_367),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_312),
.C(n_285),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_317),
.Y(n_364)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_365),
.A2(n_371),
.B1(n_340),
.B2(n_326),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_316),
.C(n_310),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_324),
.A2(n_314),
.B1(n_311),
.B2(n_286),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_379),
.B1(n_385),
.B2(n_371),
.Y(n_393)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_318),
.C(n_323),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_373),
.B(n_387),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_357),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_355),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_384),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_343),
.C(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_380),
.C(n_367),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_319),
.B1(n_343),
.B2(n_334),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_349),
.B(n_320),
.C(n_339),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_328),
.B1(n_331),
.B2(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_381),
.Y(n_401)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_382),
.Y(n_398)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_388),
.Y(n_394)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_311),
.B1(n_338),
.B2(n_330),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_369),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_286),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_308),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_391),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_340),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_390),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_308),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_362),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_393),
.A2(n_352),
.B1(n_370),
.B2(n_382),
.Y(n_421)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_405),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_375),
.B(n_354),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_403),
.B(n_404),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_379),
.A2(n_355),
.B(n_368),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_359),
.C(n_361),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_374),
.C(n_387),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_361),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_407),
.B(n_409),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_408),
.A2(n_383),
.B1(n_363),
.B2(n_370),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_391),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_402),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_408),
.A2(n_372),
.B1(n_377),
.B2(n_378),
.Y(n_412)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_380),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_415),
.C(n_417),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_389),
.C(n_388),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_392),
.C(n_385),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_419),
.A2(n_407),
.B1(n_394),
.B2(n_399),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_401),
.A2(n_364),
.B1(n_350),
.B2(n_352),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_360),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_421),
.A2(n_422),
.B1(n_398),
.B2(n_394),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_348),
.B1(n_360),
.B2(n_326),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_405),
.B1(n_396),
.B2(n_399),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_424),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_427),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_406),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_428),
.B(n_431),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_419),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_410),
.A2(n_402),
.B(n_300),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_297),
.C(n_12),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_422),
.C(n_417),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_434),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_430),
.B(n_418),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_436),
.B(n_437),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_430),
.B(n_415),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_432),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_425),
.C(n_414),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_442),
.B(n_444),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_435),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_427),
.C(n_416),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_446),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_441),
.B(n_429),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_447),
.B(n_440),
.Y(n_449)
);

O2A1O1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_449),
.A2(n_433),
.B(n_442),
.C(n_426),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

AO21x1_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_448),
.B(n_431),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_421),
.C(n_416),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_13),
.Y(n_454)
);


endmodule