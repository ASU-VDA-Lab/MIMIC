module fake_aes_3449_n_269 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_269);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_269;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_214;
wire n_267;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_244;
wire n_102;
wire n_119;
wire n_141;
wire n_115;
wire n_97;
wire n_167;
wire n_107;
wire n_158;
wire n_114;
wire n_121;
wire n_171;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_262;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_180;
wire n_137;
wire n_104;
wire n_160;
wire n_98;
wire n_154;
wire n_195;
wire n_165;
wire n_146;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_215;
wire n_108;
wire n_155;
wire n_116;
wire n_209;
wire n_217;
wire n_139;
wire n_230;
wire n_229;
wire n_198;
wire n_169;
wire n_193;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_156;
wire n_124;
wire n_238;
wire n_128;
wire n_120;
wire n_129;
wire n_206;
wire n_135;
wire n_188;
wire n_201;
wire n_197;
wire n_247;
wire n_242;
wire n_260;
wire n_127;
wire n_170;
wire n_157;
wire n_111;
wire n_210;
wire n_202;
wire n_142;
wire n_184;
wire n_245;
wire n_265;
wire n_191;
wire n_264;
wire n_232;
wire n_200;
wire n_208;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_178;
wire n_118;
wire n_258;
wire n_253;
wire n_179;
wire n_266;
wire n_131;
wire n_112;
wire n_205;
wire n_143;
wire n_213;
wire n_235;
wire n_243;
wire n_182;
wire n_263;
wire n_166;
wire n_186;
wire n_162;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_248;
wire n_268;
wire n_231;
wire n_136;
wire n_176;
wire n_144;
wire n_183;
wire n_256;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_223;
wire n_251;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_261;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_246;
wire n_153;
wire n_259;
wire n_99;
wire n_132;
wire n_109;
wire n_151;
wire n_140;
wire n_207;
wire n_257;
wire n_224;
wire n_225;
HB1xp67_ASAP7_75t_L g97 ( .A(n_34), .Y(n_97) );
CKINVDCx14_ASAP7_75t_R g98 ( .A(n_18), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_57), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_35), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_53), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_14), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_78), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_65), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_60), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_27), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_45), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_38), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_61), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_88), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_26), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_28), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_43), .Y(n_115) );
CKINVDCx14_ASAP7_75t_R g116 ( .A(n_67), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_87), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_7), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_31), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_42), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_72), .Y(n_122) );
BUFx5_ASAP7_75t_L g123 ( .A(n_56), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_90), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_91), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_92), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_51), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_70), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_23), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_64), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_15), .Y(n_133) );
INVxp67_ASAP7_75t_SL g134 ( .A(n_52), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_69), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_93), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_94), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_55), .Y(n_138) );
BUFx10_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_58), .Y(n_140) );
BUFx10_ASAP7_75t_L g141 ( .A(n_6), .Y(n_141) );
INVxp67_ASAP7_75t_SL g142 ( .A(n_75), .Y(n_142) );
BUFx5_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_22), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_9), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_37), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_17), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_44), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_50), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_46), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_33), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_101), .B(n_0), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_100), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_97), .B(n_1), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_102), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_111), .B(n_1), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_108), .B(n_2), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_112), .A2(n_114), .B1(n_149), .B2(n_118), .Y(n_159) );
INVx2_ASAP7_75t_SL g160 ( .A(n_141), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_117), .B(n_2), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_99), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_104), .B(n_10), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_157), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_154), .B(n_103), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_164), .Y(n_169) );
NAND2xp33_ASAP7_75t_L g170 ( .A(n_163), .B(n_152), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_154), .B(n_143), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_156), .B(n_109), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_165), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_173), .B(n_153), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_168), .B(n_155), .Y(n_177) );
AOI221xp5_ASAP7_75t_L g178 ( .A1(n_166), .A2(n_156), .B1(n_158), .B2(n_105), .C(n_119), .Y(n_178) );
BUFx8_ASAP7_75t_L g179 ( .A(n_174), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_167), .B(n_98), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_172), .B(n_116), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_171), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_170), .B(n_139), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_169), .B(n_106), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_175), .B(n_107), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_177), .A2(n_142), .B(n_134), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_182), .A2(n_121), .B(n_120), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_176), .A2(n_124), .B1(n_128), .B2(n_122), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_180), .B(n_110), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_185), .Y(n_190) );
AO21x1_ASAP7_75t_L g191 ( .A1(n_181), .A2(n_131), .B(n_129), .Y(n_191) );
NOR2xp33_ASAP7_75t_SL g192 ( .A(n_179), .B(n_113), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_178), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_183), .A2(n_137), .B(n_132), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_193), .B(n_184), .Y(n_195) );
OAI21x1_ASAP7_75t_L g196 ( .A1(n_187), .A2(n_145), .B(n_144), .Y(n_196) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_191), .A2(n_147), .A3(n_148), .B(n_146), .Y(n_197) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_188), .A2(n_151), .A3(n_150), .B(n_115), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_190), .Y(n_199) );
AOI21x1_ASAP7_75t_L g200 ( .A1(n_189), .A2(n_140), .B(n_138), .Y(n_200) );
AOI21x1_ASAP7_75t_L g201 ( .A1(n_194), .A2(n_143), .B(n_127), .Y(n_201) );
AO31x2_ASAP7_75t_L g202 ( .A1(n_186), .A2(n_143), .A3(n_127), .B(n_135), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_192), .B(n_3), .Y(n_203) );
AOI21x1_ASAP7_75t_L g204 ( .A1(n_200), .A2(n_162), .B(n_135), .Y(n_204) );
INVx8_ASAP7_75t_L g205 ( .A(n_203), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_196), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_202), .Y(n_207) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_201), .A2(n_126), .B(n_125), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_195), .B(n_4), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_198), .Y(n_210) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_197), .A2(n_16), .B(n_13), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_197), .B(n_5), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_199), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_210), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_205), .A2(n_133), .B1(n_136), .B2(n_130), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_206), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_212), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_209), .B(n_8), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_211), .Y(n_219) );
AOI21x1_ASAP7_75t_L g220 ( .A1(n_204), .A2(n_20), .B(n_21), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_208), .B(n_24), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_213), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_207), .A2(n_96), .B(n_25), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_210), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_210), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_213), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_217), .A2(n_29), .B1(n_30), .B2(n_32), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_214), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_222), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_223), .B(n_36), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_225), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_218), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_226), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_216), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_219), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_221), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_215), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_220), .B(n_95), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_230), .B(n_59), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_233), .B(n_62), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_240), .A2(n_63), .B1(n_66), .B2(n_68), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_229), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_235), .B(n_71), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_236), .B(n_73), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_237), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_245), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_249), .B(n_239), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_247), .B(n_231), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_250), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_253), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_254), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_255), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_256), .Y(n_257) );
XNOR2xp5_ASAP7_75t_SL g258 ( .A(n_257), .B(n_244), .Y(n_258) );
NOR3xp33_ASAP7_75t_SL g259 ( .A(n_258), .B(n_243), .C(n_242), .Y(n_259) );
AND4x1_ASAP7_75t_L g260 ( .A(n_259), .B(n_234), .C(n_228), .D(n_238), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_260), .B(n_251), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_261), .B(n_252), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_262), .Y(n_263) );
AO22x2_ASAP7_75t_L g264 ( .A1(n_263), .A2(n_248), .B1(n_241), .B2(n_246), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_264), .B(n_74), .Y(n_265) );
NAND3xp33_ASAP7_75t_SL g266 ( .A(n_265), .B(n_77), .C(n_79), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_266), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_267), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_268) );
AOI211xp5_ASAP7_75t_L g269 ( .A1(n_268), .A2(n_84), .B(n_85), .C(n_86), .Y(n_269) );
endmodule