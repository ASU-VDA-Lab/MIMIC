module fake_jpeg_9852_n_38 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_7),
.B(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

HAxp5_ASAP7_75t_SL g17 ( 
.A(n_0),
.B(n_4),
.CON(n_17),
.SN(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_12),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_12),
.C(n_21),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_15),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_26),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_14),
.B1(n_16),
.B2(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_17),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule