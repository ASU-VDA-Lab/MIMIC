module fake_jpeg_241_n_148 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_19),
.A2(n_1),
.B(n_2),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_20),
.B(n_21),
.C(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_29),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_19),
.B(n_25),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_57),
.B(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_73),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_22),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_26),
.B(n_5),
.C(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_5),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_86),
.B(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_4),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_6),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_7),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_79),
.Y(n_105)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_56),
.Y(n_95)
);

NAND2x1_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_26),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_65),
.B1(n_70),
.B2(n_64),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_70),
.B1(n_71),
.B2(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_109),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_66),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_93),
.C(n_91),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_58),
.B1(n_66),
.B2(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_68),
.B1(n_71),
.B2(n_59),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_97),
.B1(n_88),
.B2(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_115),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_85),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_118),
.C(n_77),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_99),
.B(n_82),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_83),
.C(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_96),
.C(n_108),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_88),
.B(n_86),
.Y(n_121)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_97),
.B1(n_76),
.B2(n_87),
.C(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_130),
.B(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_116),
.B1(n_114),
.B2(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_96),
.C(n_62),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_89),
.C(n_107),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_89),
.C(n_107),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_122),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_121),
.B(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_131),
.B(n_133),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_119),
.B1(n_130),
.B2(n_112),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_117),
.B1(n_53),
.B2(n_52),
.Y(n_143)
);

XOR2x1_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_78),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_133),
.B(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_142),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_134),
.A3(n_117),
.B1(n_80),
.B2(n_84),
.C1(n_52),
.C2(n_53),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_140),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_144),
.B1(n_141),
.B2(n_139),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_117),
.Y(n_148)
);


endmodule