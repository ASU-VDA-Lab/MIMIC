module fake_jpeg_30113_n_527 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_61),
.B(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_16),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_80),
.Y(n_138)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_87),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_0),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_30),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_30),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_97),
.Y(n_153)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_35),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_101),
.B(n_44),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_33),
.B(n_0),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_41),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_36),
.B1(n_51),
.B2(n_46),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_128),
.B1(n_39),
.B2(n_31),
.Y(n_170)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_144),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_36),
.B1(n_51),
.B2(n_46),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_48),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_139),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_48),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_82),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_71),
.B(n_20),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_71),
.C(n_43),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_164),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_65),
.A2(n_20),
.B(n_42),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_158),
.C(n_43),
.Y(n_171)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_79),
.B(n_19),
.C(n_42),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_165),
.Y(n_174)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_60),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_53),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_75),
.B(n_44),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_28),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_215),
.Y(n_222)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_167),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_103),
.B1(n_94),
.B2(n_58),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_168),
.A2(n_186),
.B1(n_208),
.B2(n_211),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_171),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_170),
.A2(n_175),
.B1(n_216),
.B2(n_81),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_99),
.B1(n_98),
.B2(n_73),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_182),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_180),
.Y(n_241)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_143),
.Y(n_184)
);

BUFx8_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_193),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_77),
.B1(n_45),
.B2(n_41),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_18),
.B(n_19),
.C(n_45),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_189),
.Y(n_218)
);

INVx6_ASAP7_75t_SL g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_188),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_105),
.B(n_26),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_26),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_196),
.B(n_201),
.Y(n_248)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_113),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_198),
.Y(n_219)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_200),
.Y(n_236)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_31),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_118),
.B(n_69),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_35),
.Y(n_247)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_204),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_138),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g205 ( 
.A(n_114),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_209),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_80),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_69),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_114),
.B(n_39),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_141),
.A2(n_70),
.B1(n_74),
.B2(n_85),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_120),
.C(n_132),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_220),
.B(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_174),
.C(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_141),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_126),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_145),
.C(n_156),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_247),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_224),
.B1(n_238),
.B2(n_255),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_117),
.B1(n_116),
.B2(n_126),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_249),
.B1(n_255),
.B2(n_130),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_129),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_129),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_252),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_191),
.A2(n_117),
.B1(n_116),
.B2(n_161),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_179),
.B(n_145),
.C(n_134),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_190),
.A2(n_72),
.B1(n_142),
.B2(n_107),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_107),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_226),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_267),
.B1(n_277),
.B2(n_288),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_218),
.A2(n_187),
.B(n_202),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_259),
.A2(n_266),
.B(n_246),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_262),
.Y(n_294)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_261),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_245),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_198),
.B1(n_173),
.B2(n_130),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_264),
.A2(n_269),
.B1(n_284),
.B2(n_285),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_218),
.B(n_25),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_265),
.B(n_245),
.Y(n_321)
);

O2A1O1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_225),
.A2(n_182),
.B(n_207),
.C(n_173),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_121),
.B1(n_142),
.B2(n_211),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_231),
.A2(n_188),
.B1(n_212),
.B2(n_200),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_167),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_241),
.A2(n_207),
.B1(n_192),
.B2(n_214),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_247),
.B(n_181),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_252),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_220),
.A2(n_121),
.B1(n_119),
.B2(n_131),
.Y(n_277)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_219),
.Y(n_278)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_286),
.Y(n_295)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_122),
.B1(n_177),
.B2(n_176),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_241),
.A2(n_208),
.B1(n_106),
.B2(n_110),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_237),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_222),
.A2(n_119),
.B1(n_131),
.B2(n_36),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_245),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_222),
.A2(n_25),
.B1(n_28),
.B2(n_106),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_236),
.B1(n_228),
.B2(n_244),
.Y(n_322)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_291),
.A2(n_237),
.B1(n_203),
.B2(n_199),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_217),
.B1(n_249),
.B2(n_223),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_298),
.B1(n_325),
.B2(n_274),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_263),
.A2(n_217),
.B1(n_256),
.B2(n_229),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_299),
.B(n_310),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_250),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_301),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_303),
.A2(n_268),
.B(n_274),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_243),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_309),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_235),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_260),
.B(n_248),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_242),
.C(n_248),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_324),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_265),
.B(n_221),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_312),
.B(n_321),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_275),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_263),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_276),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_258),
.B1(n_278),
.B2(n_283),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_266),
.A2(n_206),
.B(n_253),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_SL g343 ( 
.A(n_323),
.B(n_273),
.C(n_277),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_268),
.B(n_254),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_276),
.A2(n_228),
.B1(n_242),
.B2(n_235),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_289),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_326),
.Y(n_390)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_331),
.Y(n_359)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_261),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_294),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_336),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_306),
.B(n_262),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_341),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_268),
.B(n_287),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_302),
.B(n_315),
.Y(n_361)
);

AO22x1_ASAP7_75t_L g339 ( 
.A1(n_303),
.A2(n_266),
.B1(n_259),
.B2(n_267),
.Y(n_339)
);

AO22x1_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_298),
.B1(n_324),
.B2(n_301),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_296),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_309),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_342),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_343),
.A2(n_346),
.B(n_291),
.Y(n_377)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_345),
.A2(n_352),
.B1(n_358),
.B2(n_291),
.Y(n_376)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_288),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_316),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_23),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_268),
.B1(n_274),
.B2(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_325),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_319),
.A2(n_278),
.B1(n_286),
.B2(n_281),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_302),
.B(n_304),
.Y(n_370)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_320),
.A2(n_283),
.B1(n_280),
.B2(n_275),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_346),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_356),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_371),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_L g364 ( 
.A1(n_336),
.A2(n_293),
.B(n_300),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_367),
.A2(n_376),
.B1(n_343),
.B2(n_331),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_369),
.B(n_377),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_370),
.A2(n_332),
.B1(n_347),
.B2(n_328),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_339),
.A2(n_313),
.B1(n_304),
.B2(n_305),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_305),
.C(n_317),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_355),
.C(n_349),
.Y(n_391)
);

NOR3xp33_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_308),
.C(n_318),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_338),
.A2(n_317),
.B(n_280),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_381),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_342),
.B(n_253),
.Y(n_382)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_339),
.A2(n_134),
.B(n_2),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_384),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_327),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_1),
.Y(n_387)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_1),
.Y(n_388)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_392),
.C(n_404),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_349),
.C(n_354),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_360),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_412),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_397),
.B(n_384),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_340),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_402),
.Y(n_424)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_400),
.Y(n_423)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_411),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_362),
.B(n_340),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_352),
.C(n_334),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_333),
.C(n_348),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_406),
.C(n_408),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_353),
.C(n_335),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_335),
.C(n_357),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_332),
.B1(n_358),
.B2(n_91),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_86),
.C(n_159),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_417),
.C(n_370),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_361),
.B(n_86),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_378),
.Y(n_419)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_414),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_425),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_407),
.B(n_362),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_393),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_426),
.B(n_427),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_408),
.B(n_409),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_440),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_403),
.A2(n_376),
.B1(n_365),
.B2(n_363),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_430),
.A2(n_410),
.B1(n_413),
.B2(n_403),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_365),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_371),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_434),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_375),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_407),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_436),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_395),
.A2(n_373),
.B1(n_366),
.B2(n_359),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_404),
.B(n_381),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_438),
.B(n_35),
.Y(n_463)
);

XNOR2x1_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_416),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_401),
.B(n_388),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_359),
.B1(n_366),
.B2(n_379),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_442),
.B1(n_443),
.B2(n_389),
.Y(n_455)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_397),
.A2(n_382),
.B1(n_385),
.B2(n_379),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_406),
.C(n_405),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_451),
.C(n_452),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_447),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_431),
.A2(n_396),
.B(n_419),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_446),
.A2(n_429),
.B(n_3),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_399),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_450),
.B(n_440),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_399),
.C(n_417),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_385),
.C(n_418),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_432),
.A2(n_400),
.B(n_394),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_457),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_443),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_380),
.C(n_387),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_461),
.C(n_437),
.Y(n_474)
);

INVx13_ASAP7_75t_L g457 ( 
.A(n_424),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_460),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_380),
.C(n_360),
.Y(n_461)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_474),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_465),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_462),
.A2(n_428),
.B(n_420),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_468),
.A2(n_445),
.B(n_447),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_479),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_439),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_450),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_452),
.B(n_430),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_473),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_444),
.A2(n_437),
.B(n_423),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_475),
.A2(n_477),
.B(n_453),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_429),
.C(n_159),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_480),
.C(n_451),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_2),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_460),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_456),
.B(n_3),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_23),
.C(n_6),
.Y(n_480)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_482),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_486),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_494),
.C(n_495),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_5),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_492),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_467),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_472),
.A2(n_449),
.B(n_457),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_493),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_469),
.C(n_449),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_471),
.C(n_480),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_5),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_496),
.B(n_9),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_488),
.A2(n_466),
.B1(n_468),
.B2(n_481),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_506),
.C(n_484),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_491),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_503),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_23),
.C(n_9),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_504),
.A2(n_9),
.B(n_11),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_507),
.B(n_495),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_23),
.C(n_10),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_R g507 ( 
.A(n_489),
.B(n_487),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_511),
.B(n_514),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_508),
.A2(n_486),
.B(n_485),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_512),
.B(n_513),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_485),
.B(n_12),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_23),
.C(n_13),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_504),
.Y(n_517)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_500),
.C(n_501),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_14),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_11),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_519),
.A2(n_497),
.B1(n_506),
.B2(n_503),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_520),
.A2(n_521),
.B(n_522),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_518),
.B(n_13),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_11),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_11),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_14),
.Y(n_527)
);


endmodule