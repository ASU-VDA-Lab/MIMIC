module real_jpeg_4705_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_0),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_0),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_0),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_0),
.B(n_408),
.Y(n_407)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_1),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_1),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_1),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_3),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_3),
.B(n_157),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_3),
.B(n_340),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_3),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_3),
.B(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_4),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_4),
.Y(n_406)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_4),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_5),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_5),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_5),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_5),
.B(n_169),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_5),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_5),
.B(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_6),
.Y(n_381)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_6),
.Y(n_483)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_8),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_8),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_8),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_8),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_8),
.B(n_353),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_8),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_8),
.B(n_494),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_9),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_9),
.Y(n_396)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_12),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_12),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_12),
.B(n_141),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_12),
.B(n_165),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_12),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_12),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_12),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_13),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_13),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_13),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_13),
.B(n_396),
.Y(n_440)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_15),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_15),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_15),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_15),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_15),
.B(n_120),
.Y(n_289)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_17),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_17),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_17),
.B(n_42),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_17),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_17),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_18),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_18),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_18),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_18),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_18),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_18),
.B(n_320),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_19),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_19),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_19),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_19),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_19),
.B(n_141),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_19),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_19),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_35),
.B(n_78),
.C(n_535),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_48),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_28),
.B(n_48),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_30),
.A2(n_31),
.B1(n_41),
.B2(n_61),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_41),
.C(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_32),
.B(n_385),
.Y(n_384)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_52),
.C(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_43),
.Y(n_320)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_44),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_74),
.C(n_76),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_49),
.B(n_525),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_62),
.C(n_64),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_50),
.A2(n_51),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_65),
.C(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_55),
.A2(n_56),
.B1(n_70),
.B2(n_484),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_58),
.Y(n_157)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_60),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_60),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_62),
.B(n_64),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_65),
.A2(n_66),
.B1(n_486),
.B2(n_487),
.Y(n_485)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_70),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_70),
.A2(n_439),
.B1(n_440),
.B2(n_484),
.Y(n_500)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_71),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_72),
.Y(n_250)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_73),
.Y(n_348)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_73),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_526),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_76),
.Y(n_526)
);

AO21x1_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_454),
.B(n_528),
.Y(n_78)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_415),
.B(n_453),
.Y(n_79)
);

AOI21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_371),
.B(n_414),
.Y(n_80)
);

OAI21x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_324),
.B(n_370),
.Y(n_81)
);

AOI21x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_282),
.B(n_323),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_201),
.B(n_281),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_186),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_85),
.B(n_186),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_129),
.B2(n_185),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_86),
.B(n_130),
.C(n_166),
.Y(n_322)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_106),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_88),
.B(n_107),
.C(n_128),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_101),
.C(n_104),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_89),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_191)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_94),
.Y(n_208)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_94),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_94),
.Y(n_386)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_100),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_104),
.Y(n_200)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_103),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_103),
.Y(n_437)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_103),
.Y(n_474)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_105),
.Y(n_351)
);

INVx3_ASAP7_75t_SL g445 ( 
.A(n_105),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_116),
.B1(n_127),
.B2(n_128),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_115),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_111),
.Y(n_115)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_115),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_115),
.B(n_287),
.C(n_300),
.Y(n_331)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_117),
.B(n_122),
.C(n_125),
.Y(n_321)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_166),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_146),
.C(n_158),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_143),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_138),
.C(n_143),
.Y(n_184)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_136),
.Y(n_353)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_142),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_144),
.Y(n_450)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_147),
.B1(n_158),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_155),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_148),
.A2(n_149),
.B1(n_155),
.B2(n_156),
.Y(n_274)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_150),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_153),
.Y(n_309)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_160),
.B(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_160),
.B(n_463),
.Y(n_462)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g360 ( 
.A(n_163),
.Y(n_360)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_165),
.Y(n_238)
);

XOR2x1_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_182),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_167),
.B(n_183),
.C(n_184),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_168),
.B(n_176),
.C(n_180),
.Y(n_300)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_175),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_199),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_187),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_199),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_191),
.B(n_192),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_197),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_276),
.B(n_280),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_261),
.B(n_275),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_241),
.B(n_260),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_228),
.B(n_240),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_212),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_222),
.B2(n_223),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_219),
.C(n_222),
.Y(n_259)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_218),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_227),
.Y(n_245)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_235),
.B(n_239),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_259),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_259),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.C(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_256),
.C(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_271),
.C(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_322),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_322),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_302),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_286),
.C(n_302),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_299),
.B2(n_301),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_292),
.C(n_294),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_305),
.C(n_315),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_315),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_319),
.C(n_321),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_326),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_327),
.B(n_344),
.C(n_368),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_344),
.B1(n_368),
.B2(n_369),
.Y(n_328)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_332),
.B2(n_343),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_333),
.C(n_334),
.Y(n_373)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_332),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_342),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_336),
.B(n_339),
.C(n_342),
.Y(n_402)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx6_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_354),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_345),
.B(n_355),
.C(n_356),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_345),
.Y(n_538)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_349),
.CI(n_352),
.CON(n_345),
.SN(n_345)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_349),
.C(n_352),
.Y(n_411)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_365),
.B2(n_366),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_361),
.B1(n_363),
.B2(n_364),
.Y(n_358)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_359),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_364),
.C(n_365),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_361),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_361),
.A2(n_364),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_364),
.B(n_378),
.C(n_384),
.Y(n_427)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_413),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_413),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_373),
.B(n_375),
.C(n_398),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_398),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_387),
.B2(n_397),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_376),
.B(n_388),
.C(n_389),
.Y(n_421)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_382),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_383),
.A2(n_384),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_383),
.B(n_435),
.C(n_439),
.Y(n_501)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_395),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_392),
.C(n_395),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_401),
.B2(n_412),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_402),
.C(n_403),
.Y(n_417)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_411),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_407),
.B1(n_409),
.B2(n_410),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_407),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_409),
.C(n_425),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_407),
.A2(n_410),
.B1(n_429),
.B2(n_432),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_427),
.C(n_432),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_452),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_452),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_417),
.B(n_419),
.C(n_433),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_433),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_420),
.B(n_424),
.C(n_426),
.Y(n_509)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_441),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_442),
.C(n_443),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.Y(n_434)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_481),
.C(n_484),
.Y(n_480)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_448),
.C(n_451),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_449),
.B2(n_451),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_447),
.Y(n_451)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_513),
.C(n_523),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_510),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_457),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_503),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_503),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_477),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_459),
.B(n_478),
.C(n_498),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.C(n_475),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_460),
.B(n_505),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_461),
.A2(n_475),
.B1(n_476),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_461),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_466),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_467),
.C(n_470),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_464),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_498),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_490),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_485),
.B1(n_488),
.B2(n_489),
.Y(n_479)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_489),
.C(n_490),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_500),
.Y(n_499)
);

INVx6_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_483),
.Y(n_494)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_485),
.Y(n_489)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_495),
.C(n_497),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_493),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.C(n_502),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_508),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_502),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_507),
.C(n_509),
.Y(n_503)
);

FAx1_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_507),
.CI(n_509),
.CON(n_511),
.SN(n_511)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_512),
.Y(n_532)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_511),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_514),
.B(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_516),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_519),
.C(n_520),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_529),
.B(n_530),
.C(n_534),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_527),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_527),
.Y(n_534)
);


endmodule