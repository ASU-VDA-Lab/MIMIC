module fake_aes_7913_n_1408 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1408);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1408;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_659;
wire n_432;
wire n_386;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g308 ( .A(n_172), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_22), .Y(n_309) );
INVxp33_ASAP7_75t_L g310 ( .A(n_3), .Y(n_310) );
INVxp33_ASAP7_75t_SL g311 ( .A(n_267), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_195), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_47), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_20), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_219), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_264), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_168), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_60), .Y(n_318) );
CKINVDCx16_ASAP7_75t_R g319 ( .A(n_194), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_111), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_34), .Y(n_321) );
INVxp33_ASAP7_75t_SL g322 ( .A(n_88), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_68), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_205), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_17), .Y(n_325) );
CKINVDCx14_ASAP7_75t_R g326 ( .A(n_237), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_299), .B(n_236), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_35), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_112), .Y(n_329) );
INVxp33_ASAP7_75t_SL g330 ( .A(n_43), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_255), .Y(n_331) );
INVxp33_ASAP7_75t_SL g332 ( .A(n_188), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_146), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_161), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_117), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_285), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_215), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_110), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_276), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_33), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_102), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_254), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_54), .Y(n_344) );
INVxp33_ASAP7_75t_L g345 ( .A(n_270), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_42), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_70), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_49), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_222), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_93), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_247), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_9), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_54), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_204), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_31), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_75), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_176), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_259), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_63), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_304), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_34), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_115), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_178), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_166), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_274), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_235), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_217), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_289), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_288), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_293), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_31), .Y(n_371) );
INVxp33_ASAP7_75t_SL g372 ( .A(n_82), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_0), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_240), .Y(n_375) );
CKINVDCx16_ASAP7_75t_R g376 ( .A(n_257), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_163), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_173), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_182), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_287), .Y(n_380) );
CKINVDCx14_ASAP7_75t_R g381 ( .A(n_246), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_151), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_3), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_300), .Y(n_384) );
INVxp33_ASAP7_75t_SL g385 ( .A(n_12), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_191), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_105), .Y(n_387) );
INVxp33_ASAP7_75t_SL g388 ( .A(n_291), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_273), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_280), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_7), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_262), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_67), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_218), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_123), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_55), .Y(n_396) );
INVxp33_ASAP7_75t_L g397 ( .A(n_129), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_128), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_180), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_89), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_127), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_181), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_157), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_113), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g405 ( .A(n_227), .Y(n_405) );
INVxp33_ASAP7_75t_L g406 ( .A(n_106), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_171), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_98), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_121), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_252), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_71), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_29), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_6), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_51), .Y(n_414) );
INVxp33_ASAP7_75t_L g415 ( .A(n_45), .Y(n_415) );
INVxp33_ASAP7_75t_SL g416 ( .A(n_292), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_67), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_224), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_62), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_0), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_263), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_65), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_68), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_120), .Y(n_424) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_268), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_167), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_216), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_211), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_37), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_143), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_202), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_20), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_290), .Y(n_433) );
INVxp33_ASAP7_75t_SL g434 ( .A(n_141), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_82), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_70), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_49), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_15), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_203), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_30), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_272), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_103), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_44), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_130), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_17), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_269), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_52), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_156), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_233), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_198), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_208), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_126), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_85), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_30), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_243), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_78), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_14), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_86), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_169), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_321), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_364), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_334), .B(n_1), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_334), .B(n_1), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_364), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_364), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_321), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_401), .B(n_2), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_401), .B(n_2), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_347), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_364), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_407), .B(n_4), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_310), .B(n_415), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_407), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_314), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_347), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_314), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_310), .B(n_4), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g478 ( .A(n_346), .B(n_5), .C(n_6), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_314), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_345), .B(n_5), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_364), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_308), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_314), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_314), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_373), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_367), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_404), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_415), .B(n_7), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_367), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_430), .B(n_8), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_414), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_414), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_414), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
AND2x6_ASAP7_75t_L g496 ( .A(n_467), .B(n_459), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_474), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_467), .B(n_452), .Y(n_498) );
NOR2xp33_ASAP7_75t_R g499 ( .A(n_472), .B(n_326), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_474), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_472), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_472), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_474), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_467), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_486), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_485), .B(n_345), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_467), .B(n_441), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_485), .B(n_397), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_487), .B(n_397), .Y(n_510) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_489), .A2(n_315), .B(n_312), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_467), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_467), .B(n_441), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_486), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_477), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_468), .B(n_309), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_468), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_477), .Y(n_518) );
AO22x2_ASAP7_75t_L g519 ( .A1(n_478), .A2(n_327), .B1(n_313), .B2(n_318), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_474), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_487), .B(n_406), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_495), .B(n_406), .Y(n_522) );
AO22x2_ASAP7_75t_L g523 ( .A1(n_478), .A2(n_327), .B1(n_340), .B2(n_328), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_486), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_468), .B(n_348), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_486), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_474), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_495), .B(n_319), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_476), .Y(n_530) );
NAND2xp33_ASAP7_75t_R g531 ( .A(n_463), .B(n_322), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_476), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_477), .A2(n_350), .B1(n_356), .B2(n_353), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_468), .B(n_316), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_463), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_473), .B(n_426), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_486), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_463), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_468), .B(n_354), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_468), .B(n_471), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_512), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_515), .B(n_471), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_515), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_507), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_536), .Y(n_547) );
INVx4_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_496), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_518), .B(n_471), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_499), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_501), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_505), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_537), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_509), .B(n_482), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g557 ( .A(n_536), .B(n_336), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_505), .B(n_471), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_505), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_507), .Y(n_560) );
BUFx3_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_510), .B(n_480), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_516), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_531), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_517), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_521), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_521), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_516), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_522), .B(n_480), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_498), .B(n_482), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_516), .Y(n_573) );
INVx3_ASAP7_75t_SL g574 ( .A(n_502), .Y(n_574) );
INVxp33_ASAP7_75t_L g575 ( .A(n_528), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_540), .Y(n_576) );
OAI22xp5_ASAP7_75t_SL g577 ( .A1(n_502), .A2(n_323), .B1(n_456), .B2(n_420), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_540), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_542), .B(n_489), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_536), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_538), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_498), .B(n_541), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_542), .A2(n_491), .B1(n_420), .B2(n_456), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_525), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_517), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_498), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_517), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_525), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_498), .B(n_473), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
BUFx12f_ASAP7_75t_L g593 ( .A(n_525), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_533), .B(n_462), .C(n_491), .Y(n_594) );
INVx5_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_512), .A2(n_462), .B(n_471), .C(n_469), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_496), .B(n_473), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_508), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_511), .Y(n_600) );
AND2x6_ASAP7_75t_L g601 ( .A(n_508), .B(n_471), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_508), .B(n_466), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_496), .B(n_376), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_496), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_508), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_513), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_513), .B(n_399), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_513), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_513), .B(n_405), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_511), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_511), .B(n_336), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_497), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_519), .B(n_325), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_519), .B(n_466), .Y(n_614) );
INVx4_ASAP7_75t_L g615 ( .A(n_519), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_519), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_497), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_523), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_523), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_523), .Y(n_620) );
INVx4_ASAP7_75t_L g621 ( .A(n_523), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_500), .A2(n_322), .B1(n_372), .B2(n_330), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_500), .Y(n_623) );
INVx5_ASAP7_75t_L g624 ( .A(n_503), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_504), .B(n_460), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_504), .B(n_344), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_527), .B(n_311), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_527), .B(n_460), .Y(n_628) );
INVx5_ASAP7_75t_L g629 ( .A(n_503), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_529), .B(n_358), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_529), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_600), .A2(n_317), .B1(n_418), .B2(n_362), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_614), .B(n_344), .Y(n_633) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_554), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_555), .B(n_352), .Y(n_635) );
BUFx8_ASAP7_75t_SL g636 ( .A(n_565), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_547), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_547), .B(n_311), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_544), .B(n_550), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_553), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_576), .Y(n_641) );
BUFx12f_ASAP7_75t_L g642 ( .A(n_568), .Y(n_642) );
NAND2x2_ASAP7_75t_L g643 ( .A(n_577), .B(n_459), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_580), .Y(n_644) );
BUFx4f_ASAP7_75t_SL g645 ( .A(n_593), .Y(n_645) );
INVx4_ASAP7_75t_L g646 ( .A(n_593), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_552), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_580), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_546), .A2(n_422), .B1(n_393), .B2(n_361), .C(n_355), .Y(n_649) );
AO21x2_ASAP7_75t_L g650 ( .A1(n_597), .A2(n_329), .B(n_324), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_581), .B(n_355), .C(n_352), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_578), .Y(n_652) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_548), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_600), .A2(n_362), .B1(n_418), .B2(n_317), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_553), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_583), .A2(n_330), .B1(n_385), .B2(n_372), .C(n_323), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_569), .B(n_361), .Y(n_657) );
BUFx12f_ASAP7_75t_L g658 ( .A(n_568), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_579), .A2(n_588), .B1(n_596), .B2(n_572), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_575), .B(n_385), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_559), .Y(n_661) );
O2A1O1Ixp5_ASAP7_75t_L g662 ( .A1(n_571), .A2(n_331), .B(n_349), .C(n_320), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_574), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_544), .B(n_419), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_597), .A2(n_359), .B(n_374), .C(n_371), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_544), .B(n_419), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_574), .Y(n_667) );
BUFx12f_ASAP7_75t_L g668 ( .A(n_565), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_602), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_602), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_579), .A2(n_428), .B1(n_388), .B2(n_416), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_602), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_548), .B(n_332), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_550), .B(n_437), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_564), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_579), .Y(n_676) );
NAND2xp33_ASAP7_75t_L g677 ( .A(n_601), .B(n_428), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_620), .A2(n_388), .B1(n_416), .B2(n_332), .Y(n_678) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_616), .A2(n_437), .B1(n_434), .B2(n_368), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_559), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_543), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
INVx1_ASAP7_75t_SL g683 ( .A(n_626), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_562), .Y(n_684) );
AND2x6_ASAP7_75t_L g685 ( .A(n_549), .B(n_333), .Y(n_685) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_548), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_562), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_543), .Y(n_688) );
INVx4_ASAP7_75t_L g689 ( .A(n_595), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_587), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_573), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_595), .B(n_434), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_615), .A2(n_383), .B1(n_396), .B2(n_391), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_560), .B(n_460), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_575), .B(n_469), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_614), .B(n_358), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_579), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_584), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_613), .B(n_469), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_549), .Y(n_700) );
BUFx12f_ASAP7_75t_L g701 ( .A(n_614), .Y(n_701) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_561), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_626), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_561), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_587), .Y(n_705) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_595), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_615), .A2(n_400), .B1(n_412), .B2(n_411), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_616), .A2(n_381), .B1(n_384), .B2(n_368), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_589), .Y(n_709) );
BUFx2_ASAP7_75t_L g710 ( .A(n_615), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_589), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_585), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_595), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_550), .B(n_384), .Y(n_714) );
AOI21x1_ASAP7_75t_L g715 ( .A1(n_558), .A2(n_534), .B(n_532), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_621), .A2(n_417), .B1(n_423), .B2(n_413), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_586), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_594), .B(n_429), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_592), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_595), .B(n_475), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_563), .B(n_582), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_543), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_558), .A2(n_534), .B(n_532), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_619), .A2(n_403), .B1(n_435), .B2(n_432), .Y(n_725) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_604), .B(n_475), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_590), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_621), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_567), .Y(n_729) );
BUFx4f_ASAP7_75t_L g730 ( .A(n_545), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_591), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_621), .A2(n_436), .B1(n_440), .B2(n_438), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_599), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_606), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_608), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_SL g736 ( .A1(n_610), .A2(n_337), .B(n_338), .C(n_335), .Y(n_736) );
INVx2_ASAP7_75t_SL g737 ( .A(n_556), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_625), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_601), .A2(n_443), .B1(n_447), .B2(n_445), .Y(n_739) );
CKINVDCx8_ASAP7_75t_R g740 ( .A(n_551), .Y(n_740) );
BUFx3_ASAP7_75t_L g741 ( .A(n_567), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_592), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_613), .B(n_475), .Y(n_743) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_607), .B(n_453), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_622), .B(n_454), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_612), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_619), .Y(n_747) );
INVx5_ASAP7_75t_L g748 ( .A(n_567), .Y(n_748) );
INVxp33_ASAP7_75t_L g749 ( .A(n_607), .Y(n_749) );
NOR2xp67_ASAP7_75t_L g750 ( .A(n_609), .B(n_403), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_612), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_557), .A2(n_458), .B1(n_421), .B2(n_425), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_612), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_618), .Y(n_754) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_567), .Y(n_755) );
BUFx2_ASAP7_75t_L g756 ( .A(n_601), .Y(n_756) );
OR2x6_ASAP7_75t_SL g757 ( .A(n_603), .B(n_339), .Y(n_757) );
OAI21xp33_ASAP7_75t_L g758 ( .A1(n_605), .A2(n_392), .B(n_343), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_625), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_566), .Y(n_760) );
INVx4_ASAP7_75t_L g761 ( .A(n_566), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_640), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_695), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_722), .A2(n_605), .B(n_598), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_640), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_718), .B(n_557), .C(n_609), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_641), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_659), .A2(n_611), .B1(n_628), .B2(n_625), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_632), .A2(n_601), .B1(n_627), .B2(n_566), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_655), .Y(n_770) );
INVx2_ASAP7_75t_SL g771 ( .A(n_667), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_652), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_697), .A2(n_628), .B1(n_457), .B2(n_414), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_731), .B(n_601), .Y(n_774) );
O2A1O1Ixp33_ASAP7_75t_SL g775 ( .A1(n_692), .A2(n_623), .B(n_631), .C(n_630), .Y(n_775) );
AO31x2_ASAP7_75t_L g776 ( .A1(n_718), .A2(n_464), .A3(n_465), .B(n_461), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_655), .Y(n_777) );
NAND2x1p5_ASAP7_75t_L g778 ( .A(n_676), .B(n_628), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_683), .B(n_601), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_656), .B(n_457), .C(n_351), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_703), .A2(n_357), .B1(n_363), .B2(n_360), .C(n_342), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_663), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_677), .A2(n_617), .B1(n_457), .B2(n_369), .Y(n_783) );
AOI21xp33_ASAP7_75t_L g784 ( .A1(n_665), .A2(n_370), .B(n_366), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_749), .B(n_617), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_663), .B(n_457), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_662), .A2(n_629), .B(n_624), .Y(n_787) );
BUFx3_ASAP7_75t_L g788 ( .A(n_634), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_745), .A2(n_649), .B1(n_694), .B2(n_660), .C(n_635), .Y(n_789) );
AND2x6_ASAP7_75t_L g790 ( .A(n_637), .B(n_341), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_647), .Y(n_791) );
OAI21xp5_ASAP7_75t_L g792 ( .A1(n_724), .A2(n_734), .B(n_733), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_737), .Y(n_793) );
BUFx8_ASAP7_75t_SL g794 ( .A(n_634), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_657), .B(n_457), .Y(n_795) );
NOR2xp67_ASAP7_75t_L g796 ( .A(n_654), .B(n_8), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_660), .B(n_9), .Y(n_797) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_693), .B(n_377), .C(n_375), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_661), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_645), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_677), .A2(n_380), .B1(n_382), .B2(n_379), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_661), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_671), .A2(n_387), .B1(n_389), .B2(n_386), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_735), .B(n_390), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_680), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_639), .B(n_394), .Y(n_806) );
INVx1_ASAP7_75t_SL g807 ( .A(n_648), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_675), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_680), .Y(n_809) );
AOI21xp5_ASAP7_75t_SL g810 ( .A1(n_637), .A2(n_644), .B(n_653), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_684), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_746), .A2(n_629), .B(n_624), .Y(n_812) );
AOI211xp5_ASAP7_75t_L g813 ( .A1(n_725), .A2(n_402), .B(n_408), .C(n_398), .Y(n_813) );
NAND2x1p5_ASAP7_75t_L g814 ( .A(n_637), .B(n_624), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g815 ( .A1(n_645), .A2(n_424), .B1(n_431), .B2(n_410), .Y(n_815) );
INVx3_ASAP7_75t_L g816 ( .A(n_637), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_746), .A2(n_629), .B(n_624), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_679), .A2(n_442), .B1(n_444), .B2(n_439), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_684), .Y(n_819) );
O2A1O1Ixp33_ASAP7_75t_SL g820 ( .A1(n_692), .A2(n_448), .B(n_450), .C(n_446), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_699), .B(n_10), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_743), .B(n_10), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_682), .B(n_451), .Y(n_823) );
AO32x2_ASAP7_75t_L g824 ( .A1(n_721), .A2(n_486), .A3(n_490), .B1(n_461), .B2(n_464), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_697), .A2(n_455), .B1(n_365), .B2(n_378), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_740), .Y(n_826) );
INVx5_ASAP7_75t_L g827 ( .A(n_644), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_669), .B(n_624), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_648), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_687), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_687), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_691), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_754), .A2(n_365), .B1(n_378), .B2(n_341), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_690), .Y(n_834) );
BUFx4_ASAP7_75t_R g835 ( .A(n_636), .Y(n_835) );
OAI21x1_ASAP7_75t_L g836 ( .A1(n_715), .A2(n_427), .B(n_395), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_646), .B(n_11), .Y(n_837) );
AND2x6_ASAP7_75t_L g838 ( .A(n_644), .B(n_395), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_642), .Y(n_839) );
AO21x1_ASAP7_75t_SL g840 ( .A1(n_739), .A2(n_629), .B(n_96), .Y(n_840) );
OR2x2_ASAP7_75t_L g841 ( .A(n_646), .B(n_11), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_642), .A2(n_449), .B1(n_427), .B2(n_409), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_664), .B(n_12), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_749), .A2(n_449), .B1(n_494), .B2(n_484), .C(n_479), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_693), .A2(n_483), .B1(n_484), .B2(n_479), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_701), .A2(n_409), .B1(n_367), .B2(n_629), .Y(n_846) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_701), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_698), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_712), .Y(n_849) );
AOI22xp33_ASAP7_75t_SL g850 ( .A1(n_643), .A2(n_409), .B1(n_367), .B2(n_488), .Y(n_850) );
A2O1A1Ixp33_ASAP7_75t_L g851 ( .A1(n_758), .A2(n_483), .B(n_484), .C(n_479), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_717), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_727), .B(n_488), .Y(n_853) );
OR2x2_ASAP7_75t_L g854 ( .A(n_666), .B(n_13), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_690), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_674), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_633), .A2(n_492), .B(n_493), .C(n_483), .Y(n_857) );
AND2x4_ASAP7_75t_L g858 ( .A(n_670), .B(n_13), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_738), .B(n_488), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_672), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_707), .A2(n_732), .B1(n_716), .B2(n_739), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_759), .B(n_488), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_730), .B(n_14), .Y(n_863) );
AOI21xp33_ASAP7_75t_L g864 ( .A1(n_650), .A2(n_409), .B(n_367), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_658), .A2(n_409), .B1(n_488), .B2(n_492), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_658), .A2(n_493), .B1(n_494), .B2(n_492), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_705), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_678), .A2(n_494), .B1(n_493), .B2(n_461), .C(n_470), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_730), .B(n_15), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_650), .B(n_16), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_757), .B(n_16), .Y(n_871) );
AND2x2_ASAP7_75t_SL g872 ( .A(n_747), .B(n_18), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_736), .A2(n_530), .B(n_520), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_756), .B(n_18), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_643), .A2(n_530), .B1(n_535), .B2(n_520), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_678), .A2(n_490), .B1(n_464), .B2(n_465), .C(n_470), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_644), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_708), .B(n_19), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_744), .A2(n_535), .B1(n_464), .B2(n_465), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_707), .B(n_19), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_716), .B(n_21), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_710), .A2(n_23), .B1(n_21), .B2(n_22), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_SL g883 ( .A1(n_732), .A2(n_490), .B(n_465), .C(n_470), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_714), .B(n_23), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_705), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_709), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_709), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_651), .A2(n_461), .B1(n_470), .B2(n_481), .Y(n_888) );
AND2x6_ASAP7_75t_L g889 ( .A(n_653), .B(n_481), .Y(n_889) );
BUFx6f_ASAP7_75t_L g890 ( .A(n_729), .Y(n_890) );
INVx8_ASAP7_75t_L g891 ( .A(n_685), .Y(n_891) );
CKINVDCx6p67_ASAP7_75t_R g892 ( .A(n_668), .Y(n_892) );
INVx4_ASAP7_75t_SL g893 ( .A(n_685), .Y(n_893) );
INVx3_ASAP7_75t_L g894 ( .A(n_761), .Y(n_894) );
INVx3_ASAP7_75t_L g895 ( .A(n_761), .Y(n_895) );
OA21x2_ASAP7_75t_L g896 ( .A1(n_751), .A2(n_490), .B(n_481), .Y(n_896) );
BUFx8_ASAP7_75t_L g897 ( .A(n_668), .Y(n_897) );
AO31x2_ASAP7_75t_L g898 ( .A1(n_751), .A2(n_481), .A3(n_486), .B(n_26), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_761), .A2(n_486), .B1(n_503), .B2(n_524), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_711), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_711), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_719), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_719), .Y(n_903) );
INVx2_ASAP7_75t_SL g904 ( .A(n_748), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_775), .A2(n_673), .B(n_736), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_789), .A2(n_752), .B1(n_750), .B2(n_638), .C(n_696), .Y(n_906) );
BUFx2_ASAP7_75t_L g907 ( .A(n_800), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_768), .A2(n_728), .B1(n_726), .B2(n_638), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_861), .A2(n_673), .B1(n_685), .B2(n_742), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_861), .A2(n_685), .B1(n_742), .B2(n_636), .Y(n_910) );
AOI21xp33_ASAP7_75t_SL g911 ( .A1(n_872), .A2(n_24), .B(n_25), .Y(n_911) );
BUFx2_ASAP7_75t_L g912 ( .A(n_788), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_782), .B(n_726), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_789), .A2(n_685), .B1(n_753), .B2(n_720), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_768), .A2(n_753), .B1(n_700), .B2(n_748), .Y(n_915) );
OAI21x1_ASAP7_75t_L g916 ( .A1(n_836), .A2(n_688), .B(n_681), .Y(n_916) );
AND2x2_ASAP7_75t_SL g917 ( .A(n_874), .B(n_653), .Y(n_917) );
OAI22xp5_ASAP7_75t_SL g918 ( .A1(n_850), .A2(n_748), .B1(n_721), .B2(n_720), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_762), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_767), .Y(n_920) );
AOI21xp33_ASAP7_75t_L g921 ( .A1(n_766), .A2(n_720), .B(n_700), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_794), .Y(n_922) );
BUFx4f_ASAP7_75t_SL g923 ( .A(n_897), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_765), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_763), .B(n_748), .Y(n_925) );
OAI211xp5_ASAP7_75t_SL g926 ( .A1(n_813), .A2(n_688), .B(n_723), .C(n_681), .Y(n_926) );
AND2x4_ASAP7_75t_L g927 ( .A(n_893), .B(n_741), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_770), .Y(n_928) );
BUFx2_ASAP7_75t_L g929 ( .A(n_791), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_796), .A2(n_755), .B1(n_729), .B2(n_741), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_856), .B(n_760), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_880), .A2(n_760), .B1(n_723), .B2(n_755), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_764), .A2(n_755), .B(n_729), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_777), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_881), .A2(n_760), .B1(n_755), .B2(n_729), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_821), .B(n_760), .Y(n_936) );
OAI211xp5_ASAP7_75t_L g937 ( .A1(n_850), .A2(n_689), .B(n_704), .C(n_702), .Y(n_937) );
AOI21x1_ASAP7_75t_L g938 ( .A1(n_870), .A2(n_704), .B(n_702), .Y(n_938) );
AOI332xp33_ASAP7_75t_L g939 ( .A1(n_871), .A2(n_24), .A3(n_25), .B1(n_26), .B2(n_27), .B3(n_28), .C1(n_29), .C2(n_32), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_807), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_822), .B(n_27), .Y(n_941) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_864), .A2(n_503), .B(n_506), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_772), .Y(n_943) );
OA21x2_ASAP7_75t_L g944 ( .A1(n_864), .A2(n_503), .B(n_506), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_803), .B(n_28), .Y(n_945) );
BUFx2_ASAP7_75t_L g946 ( .A(n_771), .Y(n_946) );
OA21x2_ASAP7_75t_L g947 ( .A1(n_870), .A2(n_514), .B(n_506), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_797), .A2(n_704), .B1(n_702), .B2(n_686), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_808), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g950 ( .A1(n_780), .A2(n_704), .B1(n_702), .B2(n_689), .C1(n_686), .C2(n_653), .Y(n_950) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_807), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_799), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_803), .B(n_32), .Y(n_953) );
A2O1A1Ixp33_ASAP7_75t_L g954 ( .A1(n_792), .A2(n_686), .B(n_706), .C(n_713), .Y(n_954) );
OAI21x1_ASAP7_75t_L g955 ( .A1(n_792), .A2(n_686), .B(n_706), .Y(n_955) );
AOI21xp33_ASAP7_75t_SL g956 ( .A1(n_826), .A2(n_33), .B(n_35), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_781), .A2(n_713), .B1(n_706), .B2(n_526), .C(n_524), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_863), .B(n_36), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_769), .B(n_706), .Y(n_959) );
BUFx2_ASAP7_75t_L g960 ( .A(n_874), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_837), .B(n_36), .Y(n_961) );
AOI33xp33_ASAP7_75t_L g962 ( .A1(n_882), .A2(n_37), .A3(n_38), .B1(n_39), .B2(n_40), .B3(n_41), .Y(n_962) );
OAI211xp5_ASAP7_75t_SL g963 ( .A1(n_818), .A2(n_38), .B(n_39), .C(n_40), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_891), .A2(n_713), .B1(n_42), .B2(n_43), .Y(n_964) );
INVx3_ASAP7_75t_L g965 ( .A(n_891), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_802), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_801), .A2(n_713), .B1(n_44), .B2(n_45), .Y(n_967) );
OR2x2_ASAP7_75t_L g968 ( .A(n_841), .B(n_41), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g969 ( .A1(n_781), .A2(n_526), .B1(n_524), .B2(n_514), .C(n_506), .Y(n_969) );
OAI22xp33_ASAP7_75t_SL g970 ( .A1(n_858), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_869), .B(n_46), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_778), .B(n_48), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_832), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_784), .A2(n_526), .B1(n_524), .B2(n_514), .C(n_506), .Y(n_974) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_875), .A2(n_526), .B1(n_524), .B2(n_514), .C(n_506), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_829), .B(n_847), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_773), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_977) );
INVx4_ASAP7_75t_L g978 ( .A(n_891), .Y(n_978) );
AND2x4_ASAP7_75t_L g979 ( .A(n_893), .B(n_50), .Y(n_979) );
INVx8_ASAP7_75t_L g980 ( .A(n_827), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_784), .A2(n_514), .B1(n_524), .B2(n_526), .Y(n_981) );
AND2x6_ASAP7_75t_L g982 ( .A(n_893), .B(n_95), .Y(n_982) );
AND2x4_ASAP7_75t_L g983 ( .A(n_827), .B(n_53), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_858), .A2(n_514), .B1(n_526), .B2(n_56), .Y(n_984) );
O2A1O1Ixp33_ASAP7_75t_L g985 ( .A1(n_815), .A2(n_53), .B(n_55), .C(n_56), .Y(n_985) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_778), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_848), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_878), .B(n_57), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_805), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_849), .B(n_57), .Y(n_990) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_773), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_809), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_811), .Y(n_993) );
OAI21x1_ASAP7_75t_L g994 ( .A1(n_810), .A2(n_99), .B(n_97), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_827), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_852), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_795), .A2(n_58), .B1(n_59), .B2(n_61), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g998 ( .A1(n_833), .A2(n_539), .B1(n_62), .B2(n_63), .C(n_64), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_785), .A2(n_539), .B1(n_64), .B2(n_65), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_819), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_884), .A2(n_876), .B1(n_854), .B2(n_843), .Y(n_1001) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_897), .A2(n_61), .B1(n_66), .B2(n_69), .C1(n_71), .C2(n_72), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_783), .A2(n_539), .B1(n_69), .B2(n_72), .C(n_73), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_793), .B(n_66), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_825), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_1005) );
NAND2xp33_ASAP7_75t_L g1006 ( .A(n_790), .B(n_539), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_825), .A2(n_74), .B1(n_76), .B2(n_77), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_830), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_876), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_1009) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_806), .A2(n_79), .B1(n_80), .B2(n_81), .C1(n_83), .C2(n_84), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g1011 ( .A1(n_779), .A2(n_539), .B1(n_80), .B2(n_81), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_798), .A2(n_79), .B1(n_83), .B2(n_84), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_831), .Y(n_1013) );
INVx1_ASAP7_75t_SL g1014 ( .A(n_839), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_868), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_1015) );
OAI22xp5_ASAP7_75t_SL g1016 ( .A1(n_882), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_860), .B(n_90), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_827), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_786), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_868), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_1020) );
NAND2x1_ASAP7_75t_L g1021 ( .A(n_889), .B(n_100), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_834), .Y(n_1022) );
OAI21x1_ASAP7_75t_L g1023 ( .A1(n_899), .A2(n_197), .B(n_307), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_790), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_859), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_806), .B(n_94), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_779), .A2(n_94), .B1(n_539), .B2(n_104), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_774), .A2(n_101), .B1(n_107), .B2(n_108), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_774), .B(n_109), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g1030 ( .A1(n_790), .A2(n_114), .B1(n_116), .B2(n_118), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_859), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_886), .B(n_119), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_804), .A2(n_122), .B1(n_124), .B2(n_125), .Y(n_1033) );
AOI222xp33_ASAP7_75t_L g1034 ( .A1(n_804), .A2(n_131), .B1(n_132), .B2(n_133), .C1(n_134), .C2(n_135), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_823), .B(n_306), .Y(n_1035) );
OAI211xp5_ASAP7_75t_L g1036 ( .A1(n_842), .A2(n_136), .B(n_137), .C(n_138), .Y(n_1036) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_980), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_917), .A2(n_903), .B1(n_902), .B2(n_901), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_920), .Y(n_1039) );
INVxp67_ASAP7_75t_L g1040 ( .A(n_940), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_943), .Y(n_1041) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_960), .A2(n_823), .B1(n_846), .B2(n_895), .Y(n_1042) );
NOR3xp33_ASAP7_75t_L g1043 ( .A(n_906), .B(n_857), .C(n_845), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_945), .B(n_904), .Y(n_1044) );
AO22x1_ASAP7_75t_L g1045 ( .A1(n_979), .A2(n_835), .B1(n_838), .B2(n_790), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_911), .A2(n_820), .B1(n_845), .B2(n_844), .C(n_888), .Y(n_1046) );
AND2x4_ASAP7_75t_L g1047 ( .A(n_978), .B(n_894), .Y(n_1047) );
NAND5xp2_ASAP7_75t_L g1048 ( .A(n_1002), .B(n_865), .C(n_866), .D(n_844), .E(n_892), .Y(n_1048) );
OAI31xp33_ASAP7_75t_L g1049 ( .A1(n_963), .A2(n_883), .A3(n_851), .B(n_894), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_941), .B(n_900), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_949), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_953), .A2(n_840), .B1(n_838), .B2(n_764), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_919), .Y(n_1053) );
AOI21xp5_ASAP7_75t_L g1054 ( .A1(n_954), .A2(n_1006), .B(n_944), .Y(n_1054) );
OAI33xp33_ASAP7_75t_L g1055 ( .A1(n_970), .A2(n_853), .A3(n_862), .B1(n_855), .B2(n_867), .B3(n_887), .Y(n_1055) );
AOI222xp33_ASAP7_75t_L g1056 ( .A1(n_923), .A2(n_838), .B1(n_862), .B2(n_853), .C1(n_787), .C2(n_885), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_919), .Y(n_1057) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_923), .Y(n_1058) );
O2A1O1Ixp5_ASAP7_75t_SL g1059 ( .A1(n_937), .A2(n_816), .B(n_877), .C(n_787), .Y(n_1059) );
NAND2xp5_ASAP7_75t_SL g1060 ( .A(n_917), .B(n_816), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_973), .Y(n_1061) );
NAND3xp33_ASAP7_75t_L g1062 ( .A(n_956), .B(n_879), .C(n_873), .Y(n_1062) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_910), .A2(n_838), .B1(n_895), .B2(n_828), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_980), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_987), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_1016), .A2(n_828), .B1(n_889), .B2(n_873), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_961), .B(n_776), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g1068 ( .A1(n_914), .A2(n_814), .B1(n_890), .B2(n_812), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_924), .Y(n_1069) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_912), .Y(n_1070) );
OR2x2_ASAP7_75t_SL g1071 ( .A(n_968), .B(n_896), .Y(n_1071) );
OAI31xp33_ASAP7_75t_L g1072 ( .A1(n_991), .A2(n_814), .A3(n_889), .B(n_776), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_996), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_1014), .B(n_812), .Y(n_1074) );
AOI321xp33_ASAP7_75t_L g1075 ( .A1(n_1005), .A2(n_898), .A3(n_776), .B1(n_824), .B2(n_889), .C(n_145), .Y(n_1075) );
INVx2_ASAP7_75t_L g1076 ( .A(n_924), .Y(n_1076) );
NAND4xp25_ASAP7_75t_SL g1077 ( .A(n_939), .B(n_817), .C(n_898), .D(n_142), .Y(n_1077) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_991), .A2(n_890), .B1(n_817), .B2(n_896), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_1001), .A2(n_890), .B1(n_898), .B2(n_824), .C(n_147), .Y(n_1079) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_1001), .A2(n_824), .B1(n_140), .B2(n_144), .C(n_148), .Y(n_1080) );
INVx3_ASAP7_75t_L g1081 ( .A(n_980), .Y(n_1081) );
NOR2x1p5_ASAP7_75t_L g1082 ( .A(n_922), .B(n_139), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_1007), .A2(n_149), .B1(n_150), .B2(n_152), .C(n_153), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_990), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_976), .B(n_154), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_946), .B(n_155), .Y(n_1086) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_910), .A2(n_158), .B1(n_159), .B2(n_160), .C(n_162), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_1010), .A2(n_164), .B1(n_165), .B2(n_170), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_913), .B(n_305), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_929), .B(n_174), .Y(n_1090) );
OAI321xp33_ASAP7_75t_L g1091 ( .A1(n_977), .A2(n_175), .A3(n_177), .B1(n_179), .B2(n_183), .C(n_184), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_984), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_988), .A2(n_189), .B1(n_190), .B2(n_192), .Y(n_1093) );
INVx2_ASAP7_75t_L g1094 ( .A(n_928), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_940), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_951), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_926), .A2(n_193), .B1(n_196), .B2(n_199), .Y(n_1097) );
OA21x2_ASAP7_75t_L g1098 ( .A1(n_954), .A2(n_200), .B(n_201), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_928), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_985), .A2(n_206), .B1(n_207), .B2(n_209), .C(n_210), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_952), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_951), .Y(n_1102) );
OAI211xp5_ASAP7_75t_L g1103 ( .A1(n_1024), .A2(n_212), .B(n_213), .C(n_214), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_984), .A2(n_220), .B1(n_221), .B2(n_223), .Y(n_1104) );
OAI21xp5_ASAP7_75t_L g1105 ( .A1(n_909), .A2(n_225), .B(n_226), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1017), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_1026), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_1107) );
INVx3_ASAP7_75t_L g1108 ( .A(n_978), .Y(n_1108) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_909), .A2(n_231), .B1(n_232), .B2(n_234), .C(n_238), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_947), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_998), .A2(n_239), .B1(n_241), .B2(n_242), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1004), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_907), .B(n_244), .Y(n_1113) );
OAI21xp5_ASAP7_75t_L g1114 ( .A1(n_905), .A2(n_245), .B(n_248), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_958), .A2(n_249), .B1(n_250), .B2(n_251), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_971), .B(n_253), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_942), .A2(n_256), .B(n_258), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_952), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_983), .Y(n_1119) );
AOI221xp5_ASAP7_75t_L g1120 ( .A1(n_1015), .A2(n_260), .B1(n_261), .B2(n_265), .C(n_266), .Y(n_1120) );
OAI21xp33_ASAP7_75t_SL g1121 ( .A1(n_962), .A2(n_271), .B(n_275), .Y(n_1121) );
INVx1_ASAP7_75t_SL g1122 ( .A(n_995), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_1025), .A2(n_277), .B1(n_278), .B2(n_279), .Y(n_1123) );
AOI22xp33_ASAP7_75t_SL g1124 ( .A1(n_908), .A2(n_281), .B1(n_282), .B2(n_283), .Y(n_1124) );
OAI31xp33_ASAP7_75t_L g1125 ( .A1(n_1003), .A2(n_284), .A3(n_286), .B(n_294), .Y(n_1125) );
OAI211xp5_ASAP7_75t_SL g1126 ( .A1(n_962), .A2(n_295), .B(n_296), .C(n_297), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_986), .B(n_298), .Y(n_1127) );
OR2x6_ASAP7_75t_L g1128 ( .A(n_979), .B(n_301), .Y(n_1128) );
AOI33xp33_ASAP7_75t_L g1129 ( .A1(n_1015), .A2(n_1020), .A3(n_1009), .B1(n_997), .B2(n_1012), .B3(n_964), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_966), .Y(n_1130) );
OR2x6_ASAP7_75t_L g1131 ( .A(n_983), .B(n_986), .Y(n_1131) );
INVx4_ASAP7_75t_L g1132 ( .A(n_982), .Y(n_1132) );
NAND4xp75_ASAP7_75t_L g1133 ( .A(n_972), .B(n_999), .C(n_1011), .D(n_925), .Y(n_1133) );
AO21x2_ASAP7_75t_L g1134 ( .A1(n_930), .A2(n_938), .B(n_955), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_915), .A2(n_957), .B1(n_997), .B2(n_1020), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_934), .Y(n_1136) );
OA21x2_ASAP7_75t_L g1137 ( .A1(n_933), .A2(n_974), .B(n_916), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_1031), .A2(n_1009), .B1(n_1019), .B2(n_1012), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_993), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1008), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1013), .Y(n_1141) );
BUFx6f_ASAP7_75t_L g1142 ( .A(n_927), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1022), .Y(n_1143) );
OAI31xp33_ASAP7_75t_L g1144 ( .A1(n_1048), .A2(n_1077), .A3(n_1082), .B(n_1126), .Y(n_1144) );
OAI31xp33_ASAP7_75t_L g1145 ( .A1(n_1126), .A2(n_967), .A3(n_930), .B(n_918), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_1037), .Y(n_1146) );
OAI221xp5_ASAP7_75t_SL g1147 ( .A1(n_1129), .A2(n_1033), .B1(n_936), .B2(n_1034), .C(n_969), .Y(n_1147) );
AO21x2_ASAP7_75t_L g1148 ( .A1(n_1078), .A2(n_959), .B(n_921), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1053), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_1135), .A2(n_959), .B1(n_982), .B2(n_1029), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1095), .B(n_995), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1039), .B(n_1018), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1110), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1110), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1057), .B(n_989), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1069), .Y(n_1156) );
INVx3_ASAP7_75t_L g1157 ( .A(n_1132), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1041), .B(n_1018), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1076), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1094), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1099), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1101), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1118), .B(n_989), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1130), .Y(n_1164) );
OAI31xp33_ASAP7_75t_L g1165 ( .A1(n_1042), .A2(n_1027), .A3(n_1036), .B(n_965), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1096), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1132), .B(n_1131), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_1088), .A2(n_1043), .B1(n_1044), .B2(n_1074), .Y(n_1168) );
OAI33xp33_ASAP7_75t_L g1169 ( .A1(n_1102), .A2(n_931), .A3(n_1035), .B1(n_1000), .B2(n_966), .B3(n_992), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1051), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1040), .B(n_992), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1134), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1061), .B(n_1000), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1065), .Y(n_1174) );
AOI33xp33_ASAP7_75t_L g1175 ( .A1(n_1112), .A2(n_1033), .A3(n_1030), .B1(n_932), .B2(n_935), .B3(n_1028), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1073), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1177 ( .A1(n_1088), .A2(n_932), .B1(n_935), .B2(n_1028), .C(n_948), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1136), .B(n_947), .Y(n_1178) );
BUFx3_ASAP7_75t_L g1179 ( .A(n_1081), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1040), .B(n_947), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1122), .B(n_948), .Y(n_1181) );
OAI31xp33_ASAP7_75t_L g1182 ( .A1(n_1042), .A2(n_965), .A3(n_1029), .B(n_1032), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_1131), .A2(n_981), .B1(n_1021), .B2(n_975), .Y(n_1183) );
OAI21xp33_ASAP7_75t_L g1184 ( .A1(n_1121), .A2(n_981), .B(n_950), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1084), .B(n_927), .Y(n_1185) );
INVxp67_ASAP7_75t_SL g1186 ( .A(n_1038), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1070), .Y(n_1187) );
INVx5_ASAP7_75t_SL g1188 ( .A(n_1131), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1139), .B(n_942), .Y(n_1189) );
BUFx2_ASAP7_75t_L g1190 ( .A(n_1128), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1106), .B(n_982), .Y(n_1191) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1134), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1140), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_1066), .A2(n_942), .B1(n_944), .B2(n_982), .C(n_994), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1137), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1141), .B(n_944), .Y(n_1196) );
BUFx3_ASAP7_75t_L g1197 ( .A(n_1081), .Y(n_1197) );
OAI321xp33_ASAP7_75t_L g1198 ( .A1(n_1075), .A2(n_982), .A3(n_1023), .B1(n_1066), .B2(n_1128), .C(n_1087), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1143), .B(n_1067), .Y(n_1199) );
INVx1_ASAP7_75t_SL g1200 ( .A(n_1058), .Y(n_1200) );
BUFx2_ASAP7_75t_L g1201 ( .A(n_1128), .Y(n_1201) );
OAI211xp5_ASAP7_75t_L g1202 ( .A1(n_1113), .A2(n_1056), .B(n_1063), .C(n_1052), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_1043), .A2(n_1068), .B1(n_1055), .B2(n_1138), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1119), .B(n_1050), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1138), .B(n_1142), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1071), .Y(n_1206) );
NAND4xp25_ASAP7_75t_L g1207 ( .A(n_1072), .B(n_1052), .C(n_1086), .D(n_1085), .Y(n_1207) );
AOI211xp5_ASAP7_75t_L g1208 ( .A1(n_1045), .A2(n_1068), .B(n_1090), .C(n_1078), .Y(n_1208) );
AOI211xp5_ASAP7_75t_L g1209 ( .A1(n_1064), .A2(n_1116), .B(n_1089), .C(n_1092), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1098), .Y(n_1210) );
AND2x4_ASAP7_75t_L g1211 ( .A(n_1142), .B(n_1108), .Y(n_1211) );
AOI322xp5_ASAP7_75t_L g1212 ( .A1(n_1124), .A2(n_1108), .A3(n_1093), .B1(n_1111), .B2(n_1046), .C1(n_1097), .C2(n_1100), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1098), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1137), .Y(n_1214) );
INVx2_ASAP7_75t_SL g1215 ( .A(n_1142), .Y(n_1215) );
OAI211xp5_ASAP7_75t_L g1216 ( .A1(n_1124), .A2(n_1093), .B(n_1107), .C(n_1097), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1142), .Y(n_1217) );
OAI33xp33_ASAP7_75t_L g1218 ( .A1(n_1104), .A2(n_1060), .A3(n_1062), .B1(n_1127), .B2(n_1055), .B3(n_1133), .Y(n_1218) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_1047), .Y(n_1219) );
AOI222xp33_ASAP7_75t_L g1220 ( .A1(n_1105), .A2(n_1120), .B1(n_1083), .B2(n_1080), .C1(n_1109), .C2(n_1111), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1054), .B(n_1047), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1054), .B(n_1114), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1123), .B(n_1117), .Y(n_1223) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1079), .Y(n_1224) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_1117), .Y(n_1225) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_1059), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1091), .Y(n_1227) );
NAND3xp33_ASAP7_75t_L g1228 ( .A(n_1049), .B(n_1125), .C(n_1107), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1103), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1178), .B(n_1123), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1153), .B(n_1103), .Y(n_1231) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1149), .Y(n_1232) );
BUFx2_ASAP7_75t_L g1233 ( .A(n_1190), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1149), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1235 ( .A(n_1187), .B(n_1115), .Y(n_1235) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1159), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1237 ( .A(n_1218), .B(n_1202), .C(n_1228), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1170), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_1146), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1178), .B(n_1199), .Y(n_1240) );
NAND4xp25_ASAP7_75t_L g1241 ( .A(n_1144), .B(n_1168), .C(n_1203), .D(n_1208), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1199), .B(n_1189), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1170), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1153), .B(n_1154), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1174), .Y(n_1245) );
NAND4xp25_ASAP7_75t_SL g1246 ( .A(n_1200), .B(n_1209), .C(n_1216), .D(n_1212), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1154), .B(n_1206), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1206), .B(n_1166), .Y(n_1248) );
NAND2xp5_ASAP7_75t_SL g1249 ( .A(n_1190), .B(n_1201), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1176), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1159), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1189), .B(n_1196), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1253 ( .A(n_1201), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1204), .B(n_1193), .Y(n_1254) );
BUFx2_ASAP7_75t_L g1255 ( .A(n_1219), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1196), .B(n_1176), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1221), .B(n_1205), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1156), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1221), .B(n_1205), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1166), .B(n_1164), .Y(n_1260) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_1146), .Y(n_1261) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1156), .Y(n_1262) );
BUFx2_ASAP7_75t_L g1263 ( .A(n_1219), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1173), .B(n_1193), .Y(n_1264) );
AOI322xp5_ASAP7_75t_L g1265 ( .A1(n_1186), .A2(n_1204), .A3(n_1150), .B1(n_1167), .B2(n_1158), .C1(n_1152), .C2(n_1227), .Y(n_1265) );
AND2x4_ASAP7_75t_L g1266 ( .A(n_1157), .B(n_1167), .Y(n_1266) );
HB1xp67_ASAP7_75t_L g1267 ( .A(n_1151), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1173), .B(n_1151), .Y(n_1268) );
NOR3xp33_ASAP7_75t_SL g1269 ( .A(n_1207), .B(n_1198), .C(n_1147), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1160), .B(n_1162), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1157), .Y(n_1271) );
NAND4xp25_ASAP7_75t_L g1272 ( .A(n_1182), .B(n_1185), .C(n_1191), .D(n_1145), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1157), .B(n_1167), .Y(n_1273) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1179), .B(n_1197), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1160), .Y(n_1275) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1180), .B(n_1171), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1161), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_1177), .A2(n_1184), .B1(n_1223), .B2(n_1229), .Y(n_1278) );
OAI211xp5_ASAP7_75t_SL g1279 ( .A1(n_1175), .A2(n_1165), .B(n_1220), .C(n_1184), .Y(n_1279) );
AND2x4_ASAP7_75t_SL g1280 ( .A(n_1211), .B(n_1155), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1163), .B(n_1161), .Y(n_1281) );
NOR2x1p5_ASAP7_75t_L g1282 ( .A(n_1180), .B(n_1181), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1171), .B(n_1181), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_1162), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1217), .B(n_1148), .Y(n_1285) );
NAND2xp33_ASAP7_75t_L g1286 ( .A(n_1183), .B(n_1215), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1172), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1172), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1222), .B(n_1214), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1222), .B(n_1214), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1192), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1217), .B(n_1148), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1238), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1252), .B(n_1192), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1252), .B(n_1195), .Y(n_1295) );
CKINVDCx20_ASAP7_75t_R g1296 ( .A(n_1280), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1248), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1242), .B(n_1195), .Y(n_1298) );
NOR2xp67_ASAP7_75t_L g1299 ( .A(n_1246), .B(n_1194), .Y(n_1299) );
INVxp67_ASAP7_75t_L g1300 ( .A(n_1239), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1242), .B(n_1148), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1264), .B(n_1223), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1238), .Y(n_1303) );
AND2x4_ASAP7_75t_L g1304 ( .A(n_1289), .B(n_1211), .Y(n_1304) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1262), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1243), .Y(n_1306) );
NAND3xp33_ASAP7_75t_L g1307 ( .A(n_1269), .B(n_1226), .C(n_1229), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1267), .B(n_1215), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1243), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1248), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1256), .B(n_1188), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1257), .B(n_1225), .Y(n_1312) );
INVx2_ASAP7_75t_SL g1313 ( .A(n_1280), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1256), .B(n_1188), .Y(n_1314) );
INVx2_ASAP7_75t_L g1315 ( .A(n_1262), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1279), .B(n_1179), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1257), .B(n_1213), .Y(n_1317) );
AOI211x1_ASAP7_75t_SL g1318 ( .A1(n_1241), .A2(n_1227), .B(n_1224), .C(n_1169), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1283), .B(n_1210), .Y(n_1319) );
NAND2xp5_ASAP7_75t_SL g1320 ( .A(n_1274), .B(n_1197), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1283), .B(n_1210), .Y(n_1321) );
NOR4xp25_ASAP7_75t_L g1322 ( .A(n_1278), .B(n_1224), .C(n_1213), .D(n_1226), .Y(n_1322) );
AOI32xp33_ASAP7_75t_L g1323 ( .A1(n_1237), .A2(n_1188), .A3(n_1286), .B1(n_1233), .B2(n_1255), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1245), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1240), .B(n_1188), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1259), .B(n_1240), .Y(n_1326) );
INVx3_ASAP7_75t_L g1327 ( .A(n_1266), .Y(n_1327) );
AND2x4_ASAP7_75t_SL g1328 ( .A(n_1266), .B(n_1273), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1254), .B(n_1268), .Y(n_1329) );
NAND2xp5_ASAP7_75t_SL g1330 ( .A(n_1271), .B(n_1265), .Y(n_1330) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_1282), .A2(n_1261), .B1(n_1271), .B2(n_1233), .Y(n_1331) );
INVx1_ASAP7_75t_SL g1332 ( .A(n_1255), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1250), .B(n_1270), .Y(n_1333) );
OAI21xp5_ASAP7_75t_L g1334 ( .A1(n_1299), .A2(n_1249), .B(n_1253), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1297), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1336 ( .A1(n_1296), .A2(n_1282), .B1(n_1263), .B2(n_1273), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1337 ( .A(n_1326), .B(n_1276), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1293), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1303), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1310), .Y(n_1340) );
OAI221xp5_ASAP7_75t_L g1341 ( .A1(n_1316), .A2(n_1272), .B1(n_1235), .B2(n_1247), .C(n_1263), .Y(n_1341) );
HB1xp67_ASAP7_75t_L g1342 ( .A(n_1332), .Y(n_1342) );
NOR3xp33_ASAP7_75t_L g1343 ( .A(n_1307), .B(n_1330), .C(n_1331), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1302), .B(n_1290), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_1296), .A2(n_1266), .B1(n_1273), .B2(n_1276), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1333), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1303), .Y(n_1347) );
OAI21xp5_ASAP7_75t_SL g1348 ( .A1(n_1323), .A2(n_1318), .B(n_1328), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1306), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1301), .B(n_1290), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1301), .B(n_1289), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1306), .Y(n_1352) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1326), .B(n_1247), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1294), .B(n_1259), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1317), .B(n_1270), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1309), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1324), .Y(n_1357) );
NOR2xp33_ASAP7_75t_L g1358 ( .A(n_1300), .B(n_1244), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1317), .B(n_1260), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1305), .Y(n_1360) );
OAI21xp5_ASAP7_75t_SL g1361 ( .A1(n_1328), .A2(n_1313), .B(n_1320), .Y(n_1361) );
XNOR2x2_ASAP7_75t_L g1362 ( .A(n_1308), .B(n_1231), .Y(n_1362) );
NOR2xp33_ASAP7_75t_R g1363 ( .A(n_1327), .B(n_1231), .Y(n_1363) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1305), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1329), .B(n_1244), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1319), .B(n_1284), .Y(n_1366) );
AOI21xp33_ASAP7_75t_L g1367 ( .A1(n_1319), .A2(n_1292), .B(n_1285), .Y(n_1367) );
AOI221xp5_ASAP7_75t_L g1368 ( .A1(n_1322), .A2(n_1281), .B1(n_1277), .B2(n_1275), .C(n_1258), .Y(n_1368) );
INVx1_ASAP7_75t_SL g1369 ( .A(n_1304), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1304), .B(n_1266), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1294), .Y(n_1371) );
OAI22xp5_ASAP7_75t_SL g1372 ( .A1(n_1327), .A2(n_1273), .B1(n_1275), .B2(n_1258), .Y(n_1372) );
OA22x2_ASAP7_75t_L g1373 ( .A1(n_1327), .A2(n_1230), .B1(n_1232), .B2(n_1234), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1374 ( .A(n_1304), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g1375 ( .A(n_1342), .Y(n_1375) );
OAI21xp5_ASAP7_75t_L g1376 ( .A1(n_1343), .A2(n_1348), .B(n_1361), .Y(n_1376) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1366), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1341), .B(n_1346), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_1365), .A2(n_1358), .B1(n_1368), .B2(n_1345), .C(n_1367), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g1380 ( .A1(n_1334), .A2(n_1336), .B1(n_1374), .B2(n_1373), .C(n_1372), .Y(n_1380) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_1365), .A2(n_1358), .B1(n_1340), .B2(n_1335), .C(n_1363), .Y(n_1381) );
O2A1O1Ixp33_ASAP7_75t_L g1382 ( .A1(n_1362), .A2(n_1353), .B(n_1369), .C(n_1337), .Y(n_1382) );
AOI22xp5_ASAP7_75t_L g1383 ( .A1(n_1373), .A2(n_1312), .B1(n_1371), .B2(n_1344), .Y(n_1383) );
AOI22xp5_ASAP7_75t_L g1384 ( .A1(n_1312), .A2(n_1350), .B1(n_1351), .B2(n_1295), .Y(n_1384) );
A2O1A1Ixp33_ASAP7_75t_L g1385 ( .A1(n_1337), .A2(n_1353), .B(n_1370), .C(n_1354), .Y(n_1385) );
A2O1A1Ixp33_ASAP7_75t_L g1386 ( .A1(n_1354), .A2(n_1355), .B(n_1359), .C(n_1325), .Y(n_1386) );
AOI211x1_ASAP7_75t_SL g1387 ( .A1(n_1376), .A2(n_1311), .B(n_1314), .C(n_1360), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1380), .B(n_1378), .Y(n_1388) );
OAI21xp5_ASAP7_75t_SL g1389 ( .A1(n_1382), .A2(n_1230), .B(n_1321), .Y(n_1389) );
CKINVDCx20_ASAP7_75t_R g1390 ( .A(n_1375), .Y(n_1390) );
OAI21xp5_ASAP7_75t_SL g1391 ( .A1(n_1379), .A2(n_1321), .B(n_1295), .Y(n_1391) );
NAND5xp2_ASAP7_75t_L g1392 ( .A(n_1381), .B(n_1288), .C(n_1291), .D(n_1287), .E(n_1298), .Y(n_1392) );
NOR3xp33_ASAP7_75t_L g1393 ( .A(n_1388), .B(n_1385), .C(n_1386), .Y(n_1393) );
NOR3xp33_ASAP7_75t_L g1394 ( .A(n_1389), .B(n_1383), .C(n_1377), .Y(n_1394) );
OAI221xp5_ASAP7_75t_L g1395 ( .A1(n_1391), .A2(n_1384), .B1(n_1357), .B2(n_1356), .C(n_1352), .Y(n_1395) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_1390), .A2(n_1349), .B1(n_1347), .B2(n_1339), .Y(n_1396) );
XNOR2xp5_ASAP7_75t_L g1397 ( .A(n_1393), .B(n_1387), .Y(n_1397) );
NOR3xp33_ASAP7_75t_SL g1398 ( .A(n_1395), .B(n_1392), .C(n_1338), .Y(n_1398) );
NOR3xp33_ASAP7_75t_L g1399 ( .A(n_1394), .B(n_1360), .C(n_1364), .Y(n_1399) );
AOI21xp5_ASAP7_75t_L g1400 ( .A1(n_1397), .A2(n_1396), .B(n_1364), .Y(n_1400) );
XNOR2xp5_ASAP7_75t_L g1401 ( .A(n_1398), .B(n_1298), .Y(n_1401) );
AOI22x1_ASAP7_75t_SL g1402 ( .A1(n_1399), .A2(n_1315), .B1(n_1291), .B2(n_1287), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1401), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1401), .Y(n_1404) );
AOI222xp33_ASAP7_75t_L g1405 ( .A1(n_1403), .A2(n_1400), .B1(n_1402), .B2(n_1315), .C1(n_1251), .C2(n_1232), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1404), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1406), .Y(n_1407) );
AOI21xp33_ASAP7_75t_L g1408 ( .A1(n_1407), .A2(n_1405), .B(n_1236), .Y(n_1408) );
endmodule