module real_jpeg_13710_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_310, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_310;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_45),
.B1(n_50),
.B2(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_33),
.B1(n_36),
.B2(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_93),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_93),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_45),
.B1(n_50),
.B2(n_93),
.Y(n_218)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_33),
.B1(n_36),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_45),
.B1(n_50),
.B2(n_60),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_33),
.B1(n_36),
.B2(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_158),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_45),
.B1(n_50),
.B2(n_158),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_10),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_33),
.B1(n_36),
.B2(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_185),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_10),
.A2(n_45),
.B1(n_50),
.B2(n_185),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_11),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_11),
.A2(n_30),
.B1(n_53),
.B2(n_54),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_11),
.A2(n_30),
.B1(n_45),
.B2(n_50),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_12),
.A2(n_33),
.B1(n_36),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_12),
.A2(n_45),
.B1(n_50),
.B2(n_69),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_14),
.A2(n_33),
.B1(n_36),
.B2(n_134),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_134),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_14),
.A2(n_45),
.B1(n_50),
.B2(n_134),
.Y(n_252)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_15),
.B(n_188),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_15),
.B(n_36),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_15),
.A2(n_27),
.B(n_224),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_177),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_15),
.A2(n_49),
.B(n_53),
.C(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_15),
.B(n_70),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_15),
.B(n_86),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_15),
.B(n_43),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_15),
.A2(n_36),
.B(n_215),
.Y(n_278)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_17),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_17),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_17),
.A2(n_39),
.B1(n_45),
.B2(n_50),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_94),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_94),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_72),
.C(n_79),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_72),
.B1(n_73),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_24),
.A2(n_25),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_42),
.C(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_27),
.A2(n_33),
.A3(n_35),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_28),
.B(n_177),
.Y(n_176)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_31),
.A2(n_32),
.B1(n_38),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_31),
.A2(n_32),
.B1(n_92),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_31),
.A2(n_32),
.B1(n_133),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_31),
.A2(n_32),
.B1(n_184),
.B2(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_32),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_34),
.B(n_36),
.Y(n_175)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_36),
.A2(n_54),
.A3(n_64),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_57),
.B1(n_58),
.B2(n_71),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_71),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_55),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_51),
.B1(n_55),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_43),
.A2(n_51),
.B1(n_78),
.B2(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_43),
.A2(n_51),
.B1(n_90),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_43),
.A2(n_51),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_43),
.A2(n_51),
.B1(n_152),
.B2(n_209),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_43),
.A2(n_51),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_43),
.A2(n_51),
.B1(n_243),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_44),
.A2(n_129),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_44),
.A2(n_153),
.B1(n_208),
.B2(n_280),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_44)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_45),
.B(n_266),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_48),
.A2(n_50),
.B(n_177),
.Y(n_245)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_51),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_53),
.B(n_65),
.Y(n_216)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_67),
.B2(n_70),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_61),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_61),
.A2(n_70),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_61),
.A2(n_70),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_66),
.B1(n_68),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_62),
.A2(n_66),
.B1(n_76),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_62),
.A2(n_66),
.B1(n_131),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_62),
.A2(n_66),
.B1(n_180),
.B2(n_201),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_62),
.A2(n_66),
.B1(n_199),
.B2(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_91),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_81),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_87),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_84),
.A2(n_86),
.B1(n_149),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_84),
.A2(n_86),
.B1(n_173),
.B2(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_84),
.A2(n_86),
.B1(n_205),
.B2(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_84),
.A2(n_86),
.B1(n_218),
.B2(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_84),
.A2(n_86),
.B1(n_177),
.B2(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_84),
.A2(n_86),
.B1(n_257),
.B2(n_264),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_85),
.A2(n_125),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_85),
.A2(n_147),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_135),
.B(n_308),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_108),
.B(n_111),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_119),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.C(n_132),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_121),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_161),
.B(n_307),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_159),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_138),
.B(n_159),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_143),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.C(n_156),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_145),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_146),
.B(n_150),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_191),
.B(n_306),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_189),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_163),
.B(n_189),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.C(n_169),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_164),
.A2(n_165),
.B1(n_168),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_168),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_169),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.C(n_182),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_170),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_176),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_178),
.B(n_182),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_299),
.B1(n_304),
.B2(n_305),
.C(n_310),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_291),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_235),
.B(n_290),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_219),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_195),
.B(n_219),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.C(n_210),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_196),
.B(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_206),
.A2(n_210),
.B1(n_211),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_217),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_230),
.B2(n_234),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_220),
.B(n_231),
.C(n_233),
.Y(n_292)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_226),
.C(n_229),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_284),
.B(n_289),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_273),
.B(n_283),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_253),
.B(n_272),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_239),
.B(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_249),
.C(n_251),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_261),
.B(n_271),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_259),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_267),
.B(n_270),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_274),
.B(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.C(n_281),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_296),
.C(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);


endmodule