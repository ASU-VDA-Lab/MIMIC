module fake_jpeg_20412_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_20),
.Y(n_57)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_45),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_23),
.B1(n_30),
.B2(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_17),
.B(n_29),
.C(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_48),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_57),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_62),
.B1(n_70),
.B2(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_36),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_39),
.Y(n_110)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_22),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_39),
.B1(n_34),
.B2(n_37),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_39),
.B1(n_34),
.B2(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_85),
.Y(n_109)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_36),
.B(n_59),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_36),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_115),
.B(n_69),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_70),
.B1(n_86),
.B2(n_79),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_77),
.C(n_24),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_127),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_139),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_69),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_17),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_49),
.B(n_85),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_97),
.B(n_100),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_34),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_30),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_31),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_31),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_114),
.B1(n_92),
.B2(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_94),
.B1(n_97),
.B2(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_124),
.B(n_126),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_147),
.B(n_137),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_141),
.B1(n_118),
.B2(n_121),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_161),
.B1(n_165),
.B2(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_156),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_1),
.B1(n_6),
.B2(n_32),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_95),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_163),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_102),
.B1(n_112),
.B2(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_25),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_0),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_27),
.B1(n_29),
.B2(n_3),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_168),
.Y(n_178)
);

OAI322xp33_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_127),
.A3(n_134),
.B1(n_140),
.B2(n_125),
.C1(n_139),
.C2(n_136),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_144),
.C(n_153),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_181),
.B1(n_185),
.B2(n_162),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_189),
.C(n_147),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_130),
.C(n_117),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_179),
.C(n_161),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_25),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_176),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_18),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_143),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_87),
.C(n_33),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_33),
.B1(n_32),
.B2(n_5),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_33),
.B1(n_32),
.B2(n_5),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_152),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_155),
.Y(n_193)
);

NOR2x1_ASAP7_75t_R g189 ( 
.A(n_151),
.B(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_195),
.B1(n_206),
.B2(n_188),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_160),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_197),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_1),
.B(n_6),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_173),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_179),
.C(n_172),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_150),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_214),
.C(n_191),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_178),
.B1(n_182),
.B2(n_186),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_212),
.B1(n_218),
.B2(n_6),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_184),
.B(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_158),
.B1(n_149),
.B2(n_168),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_158),
.C(n_149),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_222),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_197),
.C(n_194),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_229),
.C(n_9),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_191),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_12),
.B(n_13),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_214),
.C(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_217),
.C(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_229),
.B(n_8),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_13),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_9),
.B(n_10),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_14),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_235),
.B(n_238),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_15),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_222),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

NAND2x1p5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_236),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_223),
.B(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_16),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule