module real_aes_8254_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g243 ( .A1(n_0), .A2(n_244), .B(n_245), .C(n_249), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_1), .B(n_185), .Y(n_250) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_3), .B(n_157), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_4), .A2(n_143), .B(n_148), .C(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_5), .A2(n_138), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_6), .A2(n_138), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_7), .B(n_185), .Y(n_555) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_8), .A2(n_173), .B(n_189), .Y(n_188) );
AND2x6_ASAP7_75t_L g143 ( .A(n_9), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_10), .A2(n_143), .B(n_148), .C(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g493 ( .A(n_11), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_12), .B(n_41), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_13), .B(n_248), .Y(n_513) );
INVx1_ASAP7_75t_L g167 ( .A(n_14), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_15), .B(n_157), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_16), .A2(n_158), .B(n_501), .C(n_503), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_17), .B(n_185), .Y(n_504) );
AOI22xp5_ASAP7_75t_SL g468 ( .A1(n_18), .A2(n_112), .B1(n_469), .B2(n_750), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_19), .A2(n_47), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_19), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_19), .B(n_222), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_20), .A2(n_148), .B(n_199), .C(n_218), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_21), .A2(n_197), .B(n_247), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_22), .B(n_248), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_23), .B(n_248), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_24), .Y(n_540) );
INVx1_ASAP7_75t_L g532 ( .A(n_25), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_26), .A2(n_148), .B(n_192), .C(n_199), .Y(n_191) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_28), .Y(n_509) );
INVx1_ASAP7_75t_L g589 ( .A(n_29), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_30), .A2(n_138), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g141 ( .A(n_31), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_32), .A2(n_146), .B(n_161), .C(n_207), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_33), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_34), .A2(n_247), .B(n_552), .C(n_554), .Y(n_551) );
INVxp67_ASAP7_75t_L g590 ( .A(n_35), .Y(n_590) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_36), .A2(n_46), .B1(n_129), .B2(n_130), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_36), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_37), .B(n_194), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_38), .A2(n_148), .B(n_199), .C(n_531), .Y(n_530) );
CKINVDCx14_ASAP7_75t_R g550 ( .A(n_39), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_40), .A2(n_45), .B1(n_476), .B2(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_40), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_42), .A2(n_249), .B(n_491), .C(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_43), .B(n_216), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_44), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_45), .Y(n_476) );
INVx1_ASAP7_75t_L g130 ( .A(n_46), .Y(n_130) );
INVx1_ASAP7_75t_L g126 ( .A(n_47), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_48), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_49), .B(n_138), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_50), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_51), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_52), .A2(n_146), .B(n_151), .C(n_161), .Y(n_145) );
INVx1_ASAP7_75t_L g246 ( .A(n_53), .Y(n_246) );
INVx1_ASAP7_75t_L g152 ( .A(n_54), .Y(n_152) );
INVx1_ASAP7_75t_L g521 ( .A(n_55), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_56), .B(n_138), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_57), .Y(n_225) );
CKINVDCx14_ASAP7_75t_R g489 ( .A(n_58), .Y(n_489) );
INVx1_ASAP7_75t_L g144 ( .A(n_59), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_60), .B(n_138), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_61), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_62), .A2(n_179), .B(n_181), .C(n_183), .Y(n_178) );
INVx1_ASAP7_75t_L g166 ( .A(n_63), .Y(n_166) );
INVx1_ASAP7_75t_SL g553 ( .A(n_64), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_66), .B(n_157), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_67), .B(n_185), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_68), .B(n_158), .Y(n_260) );
INVx1_ASAP7_75t_L g543 ( .A(n_69), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_70), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_71), .B(n_154), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_72), .A2(n_148), .B(n_161), .C(n_231), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_73), .Y(n_177) );
INVx1_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_75), .A2(n_105), .B1(n_116), .B2(n_754), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_76), .A2(n_138), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_77), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_78), .A2(n_138), .B(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_79), .A2(n_471), .B1(n_472), .B2(n_478), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_79), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_80), .A2(n_216), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g499 ( .A(n_81), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_82), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_83), .B(n_153), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_84), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_84), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_85), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_86), .A2(n_138), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g502 ( .A(n_87), .Y(n_502) );
INVx2_ASAP7_75t_L g164 ( .A(n_88), .Y(n_164) );
INVx1_ASAP7_75t_L g512 ( .A(n_89), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_90), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_91), .B(n_248), .Y(n_261) );
INVx2_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
OR2x2_ASAP7_75t_L g464 ( .A(n_92), .B(n_112), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_93), .A2(n_148), .B(n_161), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_94), .B(n_138), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_95), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g208 ( .A(n_96), .Y(n_208) );
INVxp67_ASAP7_75t_L g182 ( .A(n_97), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_98), .B(n_173), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_99), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g232 ( .A(n_100), .Y(n_232) );
INVx1_ASAP7_75t_L g256 ( .A(n_101), .Y(n_256) );
INVx2_ASAP7_75t_L g524 ( .A(n_102), .Y(n_524) );
AND2x2_ASAP7_75t_L g168 ( .A(n_103), .B(n_163), .Y(n_168) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g754 ( .A(n_106), .Y(n_754) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g751 ( .A(n_110), .Y(n_751) );
NOR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx2_ASAP7_75t_L g480 ( .A(n_111), .Y(n_480) );
INVx1_ASAP7_75t_L g749 ( .A(n_111), .Y(n_749) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_467), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g753 ( .A(n_120), .Y(n_753) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_461), .B(n_465), .Y(n_122) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
XOR2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_131), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_131), .A2(n_480), .B1(n_481), .B2(n_748), .Y(n_479) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR5x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_334), .C(n_412), .D(n_436), .E(n_453), .Y(n_132) );
OAI211xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_200), .B(n_251), .C(n_311), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
AND2x2_ASAP7_75t_L g265 ( .A(n_135), .B(n_171), .Y(n_265) );
INVx5_ASAP7_75t_SL g293 ( .A(n_135), .Y(n_293) );
AND2x2_ASAP7_75t_L g329 ( .A(n_135), .B(n_314), .Y(n_329) );
OR2x2_ASAP7_75t_L g368 ( .A(n_135), .B(n_170), .Y(n_368) );
OR2x2_ASAP7_75t_L g399 ( .A(n_135), .B(n_290), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_135), .B(n_303), .Y(n_435) );
AND2x2_ASAP7_75t_L g447 ( .A(n_135), .B(n_290), .Y(n_447) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_168), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_145), .B(n_163), .Y(n_136) );
BUFx2_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_139), .B(n_143), .Y(n_257) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
INVx1_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
INVx1_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
INVx3_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
INVx1_ASAP7_75t_L g194 ( .A(n_142), .Y(n_194) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_142), .Y(n_248) );
INVx4_ASAP7_75t_SL g162 ( .A(n_143), .Y(n_162) );
BUFx3_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_147), .A2(n_162), .B(n_177), .C(n_178), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_147), .A2(n_162), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_147), .A2(n_162), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_147), .A2(n_162), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g520 ( .A1(n_147), .A2(n_162), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_147), .A2(n_162), .B(n_550), .C(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_SL g585 ( .A1(n_147), .A2(n_162), .B(n_586), .C(n_587), .Y(n_585) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx3_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_149), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_156), .C(n_159), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_153), .A2(n_159), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_153), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_153), .A2(n_514), .B(n_543), .C(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_157), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g244 ( .A(n_157), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_157), .A2(n_221), .B(n_532), .C(n_533), .Y(n_531) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_157), .A2(n_180), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_158), .B(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g249 ( .A(n_160), .Y(n_249) );
INVx1_ASAP7_75t_L g503 ( .A(n_160), .Y(n_503) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_163), .A2(n_205), .B(n_206), .Y(n_204) );
INVx2_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_163), .Y(n_226) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_163), .A2(n_487), .B(n_494), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_163), .A2(n_257), .B(n_529), .C(n_530), .Y(n_528) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AND2x2_ASAP7_75t_L g174 ( .A(n_164), .B(n_165), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AND2x2_ASAP7_75t_L g446 ( .A(n_169), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g309 ( .A(n_170), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_187), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_171), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_171), .Y(n_302) );
INVx3_ASAP7_75t_L g317 ( .A(n_171), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_171), .B(n_187), .Y(n_341) );
OR2x2_ASAP7_75t_L g350 ( .A(n_171), .B(n_293), .Y(n_350) );
AND2x2_ASAP7_75t_L g354 ( .A(n_171), .B(n_314), .Y(n_354) );
AND2x2_ASAP7_75t_L g360 ( .A(n_171), .B(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g397 ( .A(n_171), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_171), .B(n_254), .Y(n_411) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_184), .Y(n_171) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_172), .A2(n_497), .B(n_504), .Y(n_496) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_172), .A2(n_519), .B(n_525), .Y(n_518) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_172), .A2(n_548), .B(n_555), .Y(n_547) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g186 ( .A(n_173), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_190), .B(n_191), .Y(n_189) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g264 ( .A(n_174), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_179), .A2(n_232), .B(n_233), .C(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_180), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_180), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g221 ( .A(n_183), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_183), .B(n_588), .Y(n_587) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_185), .A2(n_240), .B(n_250), .Y(n_239) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_186), .B(n_211), .Y(n_210) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_186), .A2(n_229), .B(n_237), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_186), .B(n_238), .Y(n_237) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_255), .B(n_262), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_186), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_186), .B(n_535), .Y(n_534) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_186), .A2(n_539), .B(n_545), .Y(n_538) );
OR2x2_ASAP7_75t_L g303 ( .A(n_187), .B(n_254), .Y(n_303) );
AND2x2_ASAP7_75t_L g314 ( .A(n_187), .B(n_290), .Y(n_314) );
AND2x2_ASAP7_75t_L g326 ( .A(n_187), .B(n_317), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_187), .B(n_254), .Y(n_349) );
INVx1_ASAP7_75t_SL g361 ( .A(n_187), .Y(n_361) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g253 ( .A(n_188), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_188), .B(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_195), .B(n_196), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_196), .A2(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
AND2x2_ASAP7_75t_L g274 ( .A(n_202), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_202), .B(n_227), .Y(n_278) );
AND2x2_ASAP7_75t_L g281 ( .A(n_202), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_202), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g306 ( .A(n_202), .B(n_297), .Y(n_306) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_202), .Y(n_325) );
AND2x2_ASAP7_75t_L g346 ( .A(n_202), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g356 ( .A(n_202), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g402 ( .A(n_202), .B(n_285), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_202), .B(n_308), .Y(n_429) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g299 ( .A(n_203), .Y(n_299) );
AND2x2_ASAP7_75t_L g365 ( .A(n_203), .B(n_297), .Y(n_365) );
AND2x2_ASAP7_75t_L g449 ( .A(n_203), .B(n_317), .Y(n_449) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_210), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_212), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_212), .Y(n_438) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_227), .Y(n_212) );
AND2x2_ASAP7_75t_L g268 ( .A(n_213), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g277 ( .A(n_213), .B(n_275), .Y(n_277) );
INVx5_ASAP7_75t_L g285 ( .A(n_213), .Y(n_285) );
AND2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_239), .Y(n_308) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_213), .Y(n_345) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_217), .B(n_222), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_223), .B(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_226), .A2(n_508), .B(n_515), .Y(n_507) );
INVx1_ASAP7_75t_L g386 ( .A(n_227), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_227), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g419 ( .A(n_227), .B(n_285), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_227), .A2(n_342), .B(n_449), .C(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_239), .Y(n_227) );
BUFx2_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
INVx2_ASAP7_75t_L g273 ( .A(n_228), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g554 ( .A(n_235), .Y(n_554) );
INVx2_ASAP7_75t_L g275 ( .A(n_239), .Y(n_275) );
AND2x2_ASAP7_75t_L g282 ( .A(n_239), .B(n_273), .Y(n_282) );
AND2x2_ASAP7_75t_L g373 ( .A(n_239), .B(n_285), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_247), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g491 ( .A(n_248), .Y(n_491) );
INVx2_ASAP7_75t_L g514 ( .A(n_249), .Y(n_514) );
AOI211x1_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_266), .B(n_279), .C(n_304), .Y(n_251) );
INVx1_ASAP7_75t_L g370 ( .A(n_252), .Y(n_370) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_265), .Y(n_252) );
INVx5_ASAP7_75t_SL g290 ( .A(n_254), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_254), .B(n_360), .Y(n_359) );
AOI311xp33_ASAP7_75t_L g378 ( .A1(n_254), .A2(n_379), .A3(n_381), .B(n_382), .C(n_388), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g413 ( .A1(n_254), .A2(n_326), .B(n_414), .C(n_417), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_258), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_257), .A2(n_509), .B(n_510), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_257), .A2(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g582 ( .A(n_264), .Y(n_582) );
INVxp67_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
NAND4xp25_ASAP7_75t_SL g266 ( .A(n_267), .B(n_270), .C(n_276), .D(n_278), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_267), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g324 ( .A(n_268), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_271), .B(n_277), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_271), .B(n_284), .Y(n_404) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_272), .B(n_285), .Y(n_422) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
INVxp67_ASAP7_75t_L g332 ( .A(n_274), .Y(n_332) );
AND2x4_ASAP7_75t_L g284 ( .A(n_275), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g358 ( .A(n_275), .B(n_297), .Y(n_358) );
INVx1_ASAP7_75t_L g385 ( .A(n_275), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_275), .B(n_372), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_276), .B(n_346), .Y(n_366) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_277), .B(n_299), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_277), .B(n_346), .Y(n_445) );
INVx1_ASAP7_75t_L g456 ( .A(n_278), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_283), .B(n_286), .C(n_294), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g336 ( .A(n_282), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g318 ( .A(n_283), .Y(n_318) );
AND2x2_ASAP7_75t_L g295 ( .A(n_284), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_284), .B(n_346), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_284), .B(n_365), .Y(n_389) );
OR2x2_ASAP7_75t_L g305 ( .A(n_285), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_285), .B(n_297), .Y(n_352) );
AND2x2_ASAP7_75t_L g409 ( .A(n_285), .B(n_365), .Y(n_409) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_285), .Y(n_416) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_287), .A2(n_299), .B1(n_421), .B2(n_423), .C(n_426), .Y(n_420) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g310 ( .A(n_290), .B(n_293), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_290), .B(n_360), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_290), .B(n_317), .Y(n_425) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g410 ( .A(n_292), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g424 ( .A(n_292), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_293), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g321 ( .A(n_293), .B(n_314), .Y(n_321) );
AND2x2_ASAP7_75t_L g391 ( .A(n_293), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_293), .B(n_340), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_293), .B(n_441), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_298), .B(n_300), .Y(n_294) );
INVx2_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
OR2x2_ASAP7_75t_L g351 ( .A(n_299), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g454 ( .A(n_299), .B(n_422), .Y(n_454) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI21xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_307), .B(n_309), .Y(n_304) );
INVx1_ASAP7_75t_L g458 ( .A(n_305), .Y(n_458) );
INVx2_ASAP7_75t_SL g372 ( .A(n_306), .Y(n_372) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_309), .A2(n_390), .B(n_454), .C(n_455), .Y(n_453) );
OAI322xp33_ASAP7_75t_SL g322 ( .A1(n_310), .A2(n_323), .A3(n_326), .B1(n_327), .B2(n_328), .C1(n_330), .C2(n_333), .Y(n_322) );
INVx2_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_318), .B1(n_319), .B2(n_321), .C(n_322), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp33_ASAP7_75t_SL g388 ( .A1(n_313), .A2(n_389), .B1(n_390), .B2(n_393), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_314), .B(n_317), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_314), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g387 ( .A(n_316), .B(n_349), .Y(n_387) );
INVx1_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_321), .A2(n_431), .B(n_433), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_323), .A2(n_356), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g384 ( .A(n_325), .B(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_325), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g441 ( .A(n_326), .Y(n_441) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND4xp25_ASAP7_75t_L g334 ( .A(n_335), .B(n_362), .C(n_378), .D(n_394), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B(n_343), .C(n_355), .Y(n_335) );
INVx1_ASAP7_75t_L g427 ( .A(n_336), .Y(n_427) );
AND2x2_ASAP7_75t_L g375 ( .A(n_337), .B(n_358), .Y(n_375) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_342), .B(n_377), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_351), .B2(n_353), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_345), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g407 ( .A1(n_346), .A2(n_385), .B(n_408), .C(n_410), .Y(n_407) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx1_ASAP7_75t_L g452 ( .A(n_350), .Y(n_452) );
NAND2xp33_ASAP7_75t_SL g442 ( .A(n_351), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g381 ( .A(n_360), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B(n_367), .C(n_369), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_374), .B2(n_376), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_372), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_377), .B(n_398), .Y(n_460) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_386), .B(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_400), .B1(n_403), .B2(n_405), .C(n_407), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_410), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_426) );
NAND3xp33_ASAP7_75t_SL g412 ( .A(n_413), .B(n_420), .C(n_430), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_439), .C(n_448), .Y(n_436) );
INVx1_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_444), .B2(n_446), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g466 ( .A(n_464), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_465), .B(n_468), .C(n_752), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_678), .Y(n_481) );
NAND5xp2_ASAP7_75t_L g482 ( .A(n_483), .B(n_593), .C(n_625), .D(n_642), .E(n_665), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_526), .B1(n_556), .B2(n_560), .C(n_564), .Y(n_483) );
INVx1_ASAP7_75t_L g705 ( .A(n_484), .Y(n_705) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_505), .Y(n_484) );
AND3x2_ASAP7_75t_L g680 ( .A(n_485), .B(n_507), .C(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_486), .B(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g571 ( .A(n_486), .Y(n_571) );
AND2x2_ASAP7_75t_L g575 ( .A(n_486), .B(n_517), .Y(n_575) );
INVx2_ASAP7_75t_L g602 ( .A(n_486), .Y(n_602) );
OR2x2_ASAP7_75t_L g613 ( .A(n_486), .B(n_518), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_486), .B(n_506), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_486), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g692 ( .A(n_486), .B(n_518), .Y(n_692) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_495), .Y(n_574) );
AND2x2_ASAP7_75t_L g633 ( .A(n_495), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_495), .B(n_506), .Y(n_652) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g563 ( .A(n_496), .B(n_506), .Y(n_563) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
AND2x2_ASAP7_75t_L g619 ( .A(n_496), .B(n_518), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_496), .B(n_505), .C(n_602), .Y(n_644) );
AND2x2_ASAP7_75t_L g709 ( .A(n_496), .B(n_507), .Y(n_709) );
AND2x2_ASAP7_75t_L g743 ( .A(n_496), .B(n_506), .Y(n_743) );
INVxp67_ASAP7_75t_L g572 ( .A(n_505), .Y(n_572) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_506), .B(n_602), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_506), .B(n_633), .Y(n_641) );
AND2x2_ASAP7_75t_L g691 ( .A(n_506), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g719 ( .A(n_506), .Y(n_719) );
INVx4_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g626 ( .A(n_507), .B(n_619), .Y(n_626) );
BUFx3_ASAP7_75t_L g658 ( .A(n_507), .Y(n_658) );
INVx2_ASAP7_75t_L g634 ( .A(n_517), .Y(n_634) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_518), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_526), .A2(n_694), .B1(n_696), .B2(n_697), .Y(n_693) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
AND2x2_ASAP7_75t_L g556 ( .A(n_527), .B(n_557), .Y(n_556) );
INVx3_ASAP7_75t_SL g567 ( .A(n_527), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_527), .B(n_597), .Y(n_629) );
OR2x2_ASAP7_75t_L g648 ( .A(n_527), .B(n_537), .Y(n_648) );
AND2x2_ASAP7_75t_L g653 ( .A(n_527), .B(n_605), .Y(n_653) );
AND2x2_ASAP7_75t_L g656 ( .A(n_527), .B(n_598), .Y(n_656) );
AND2x2_ASAP7_75t_L g668 ( .A(n_527), .B(n_547), .Y(n_668) );
AND2x2_ASAP7_75t_L g684 ( .A(n_527), .B(n_538), .Y(n_684) );
AND2x4_ASAP7_75t_L g687 ( .A(n_527), .B(n_558), .Y(n_687) );
OR2x2_ASAP7_75t_L g704 ( .A(n_527), .B(n_640), .Y(n_704) );
OR2x2_ASAP7_75t_L g735 ( .A(n_527), .B(n_580), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_527), .B(n_663), .Y(n_737) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
AND2x2_ASAP7_75t_L g611 ( .A(n_536), .B(n_578), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_536), .B(n_598), .Y(n_730) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_547), .Y(n_536) );
AND2x2_ASAP7_75t_L g566 ( .A(n_537), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g605 ( .A(n_537), .B(n_580), .Y(n_605) );
AND2x2_ASAP7_75t_L g623 ( .A(n_537), .B(n_558), .Y(n_623) );
OR2x2_ASAP7_75t_L g640 ( .A(n_537), .B(n_598), .Y(n_640) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g559 ( .A(n_538), .Y(n_559) );
AND2x2_ASAP7_75t_L g663 ( .A(n_538), .B(n_547), .Y(n_663) );
INVx2_ASAP7_75t_L g558 ( .A(n_547), .Y(n_558) );
INVx1_ASAP7_75t_L g675 ( .A(n_547), .Y(n_675) );
AND2x2_ASAP7_75t_L g725 ( .A(n_547), .B(n_567), .Y(n_725) );
AND2x2_ASAP7_75t_L g577 ( .A(n_557), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g609 ( .A(n_557), .B(n_567), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_557), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g596 ( .A(n_558), .B(n_567), .Y(n_596) );
OR2x2_ASAP7_75t_L g712 ( .A(n_559), .B(n_686), .Y(n_712) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_562), .B(n_692), .Y(n_698) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OAI32xp33_ASAP7_75t_L g654 ( .A1(n_563), .A2(n_655), .A3(n_657), .B1(n_659), .B2(n_660), .Y(n_654) );
OR2x2_ASAP7_75t_L g671 ( .A(n_563), .B(n_613), .Y(n_671) );
OAI21xp33_ASAP7_75t_SL g696 ( .A1(n_563), .A2(n_573), .B(n_601), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B1(n_573), .B2(n_576), .Y(n_564) );
INVxp33_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_566), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_567), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g622 ( .A(n_567), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g722 ( .A(n_567), .B(n_663), .Y(n_722) );
OR2x2_ASAP7_75t_L g746 ( .A(n_567), .B(n_640), .Y(n_746) );
AOI21xp33_ASAP7_75t_L g729 ( .A1(n_568), .A2(n_628), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_570), .B(n_575), .Y(n_624) );
AND2x2_ASAP7_75t_L g646 ( .A(n_571), .B(n_619), .Y(n_646) );
INVx1_ASAP7_75t_L g659 ( .A(n_571), .Y(n_659) );
OR2x2_ASAP7_75t_L g664 ( .A(n_571), .B(n_598), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_574), .B(n_613), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_575), .A2(n_595), .B1(n_600), .B2(n_604), .Y(n_594) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_578), .A2(n_637), .B1(n_644), .B2(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g721 ( .A(n_578), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_580), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g740 ( .A(n_580), .B(n_623), .Y(n_740) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .B(n_591), .Y(n_580) );
INVx1_ASAP7_75t_L g599 ( .A(n_581), .Y(n_599) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_584), .A2(n_592), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_606), .B1(n_607), .B2(n_612), .C(n_614), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_598), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_596), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g615 ( .A(n_597), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_597), .A2(n_703), .B(n_704), .C(n_705), .Y(n_702) );
AND2x2_ASAP7_75t_L g707 ( .A(n_597), .B(n_687), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_SL g745 ( .A1(n_597), .A2(n_686), .B(n_746), .C(n_747), .Y(n_745) );
BUFx3_ASAP7_75t_L g637 ( .A(n_598), .Y(n_637) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_601), .B(n_658), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g720 ( .A1(n_601), .A2(n_721), .B(n_723), .C(n_729), .Y(n_720) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVxp67_ASAP7_75t_L g681 ( .A(n_603), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_605), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_609), .A2(n_626), .B(n_627), .C(n_635), .Y(n_625) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g710 ( .A(n_613), .Y(n_710) );
OR2x2_ASAP7_75t_L g727 ( .A(n_613), .B(n_657), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_621), .B2(n_624), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_616), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
OR2x2_ASAP7_75t_L g714 ( .A(n_618), .B(n_658), .Y(n_714) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g669 ( .A(n_619), .B(n_659), .Y(n_669) );
INVx1_ASAP7_75t_L g677 ( .A(n_620), .Y(n_677) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_623), .B(n_637), .Y(n_685) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_633), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g742 ( .A(n_634), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g672 ( .A(n_636), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_637), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_637), .B(n_668), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_637), .B(n_663), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_637), .B(n_684), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_637), .A2(n_647), .B(n_687), .C(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AOI221xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_647), .B1(n_649), .B2(n_653), .C(n_654), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_651), .B(n_659), .Y(n_733) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_653), .A2(n_668), .B(n_670), .C(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_656), .B(n_663), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_657), .B(n_710), .Y(n_747) );
CKINVDCx16_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
INVxp33_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
AOI21xp33_ASAP7_75t_SL g673 ( .A1(n_662), .A2(n_674), .B(n_676), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_662), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_663), .B(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B1(n_670), .B2(n_672), .C(n_673), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_669), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g703 ( .A(n_675), .Y(n_703) );
NAND5xp2_ASAP7_75t_L g678 ( .A(n_679), .B(n_706), .C(n_720), .D(n_731), .E(n_744), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B(n_689), .C(n_702), .Y(n_679) );
INVx2_ASAP7_75t_SL g726 ( .A(n_680), .Y(n_726) );
NAND4xp25_ASAP7_75t_SL g682 ( .A(n_683), .B(n_685), .C(n_686), .D(n_688), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_688), .A2(n_690), .B(n_693), .C(n_699), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_691), .A2(n_732), .B1(n_734), .B2(n_736), .C(n_738), .Y(n_731) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI221xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_708), .B1(n_711), .B2(n_713), .C(n_715), .Y(n_706) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_714), .A2(n_737), .B1(n_739), .B2(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule