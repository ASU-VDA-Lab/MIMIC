module fake_ibex_562_n_713 (n_85, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_63, n_98, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_112, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_123, n_24, n_52, n_99, n_105, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_117, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_713);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_123;
input n_24;
input n_52;
input n_99;
input n_105;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_713;

wire n_151;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_688;
wire n_130;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_652;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_645;
wire n_500;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_383;
wire n_561;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_673;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_127;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_136;
wire n_261;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_636;
wire n_594;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_137;
wire n_679;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_672;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_135;
wire n_520;
wire n_684;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_405;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_639;
wire n_303;
wire n_362;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_668;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_231;
wire n_298;
wire n_202;
wire n_587;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_L g133 ( 
.A(n_9),
.B(n_48),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_81),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_71),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g140 ( 
.A(n_43),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_27),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_16),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_42),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_65),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_54),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_19),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_68),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_39),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_66),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_57),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_88),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_46),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_91),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_73),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_53),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_36),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_94),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_59),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_95),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_41),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_52),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_45),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_99),
.B(n_35),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_49),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_51),
.Y(n_184)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_32),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_64),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_23),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_28),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_61),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_38),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_9),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_110),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_86),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_93),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_92),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_143),
.B(n_0),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_134),
.B(n_33),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

OAI22x1_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

OAI22x1_ASAP7_75t_SL g217 ( 
.A1(n_197),
.A2(n_207),
.B1(n_185),
.B2(n_135),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_2),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_136),
.A2(n_63),
.B(n_124),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx8_ASAP7_75t_R g222 ( 
.A(n_162),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_168),
.A2(n_62),
.B(n_121),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g224 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_5),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_13),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_13),
.Y(n_237)
);

BUFx8_ASAP7_75t_L g238 ( 
.A(n_126),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_128),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_135),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_160),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

OAI22x1_ASAP7_75t_SL g245 ( 
.A1(n_160),
.A2(n_173),
.B1(n_166),
.B2(n_167),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_20),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_127),
.Y(n_249)
);

OAI22x1_ASAP7_75t_SL g250 ( 
.A1(n_166),
.A2(n_172),
.B1(n_167),
.B2(n_173),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_130),
.B(n_34),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx6p67_ASAP7_75t_R g253 ( 
.A(n_172),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_137),
.B(n_20),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_144),
.B(n_21),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_148),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

CKINVDCx6p67_ASAP7_75t_R g260 ( 
.A(n_181),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_151),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_157),
.B(n_25),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_158),
.B(n_25),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_244),
.B(n_184),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_152),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_163),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_214),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_211),
.B(n_189),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_208),
.A2(n_191),
.B1(n_196),
.B2(n_204),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_214),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

OR2x6_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_133),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_212),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_216),
.B(n_26),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_259),
.B(n_139),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

OR2x6_ASAP7_75t_L g301 ( 
.A(n_224),
.B(n_181),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_147),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_149),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_213),
.B(n_161),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_234),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_164),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_222),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_249),
.B(n_155),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_253),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_213),
.B(n_165),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_219),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_251),
.B(n_174),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_219),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_223),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_159),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_223),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_255),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_273),
.B(n_231),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_297),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_253),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_272),
.B(n_257),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_333),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_238),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_309),
.A2(n_256),
.B1(n_264),
.B2(n_254),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_260),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_317),
.B(n_265),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_226),
.Y(n_349)
);

AOI221xp5_ASAP7_75t_L g350 ( 
.A1(n_281),
.A2(n_261),
.B1(n_217),
.B2(n_248),
.C(n_215),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_243),
.C(n_240),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_325),
.A2(n_138),
.B1(n_153),
.B2(n_188),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_179),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_245),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_169),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_171),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_268),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_146),
.Y(n_360)
);

AO22x2_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_250),
.B1(n_322),
.B2(n_301),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_199),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_267),
.B(n_200),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_203),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_288),
.B(n_205),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_274),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_280),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_268),
.B(n_278),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_268),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_277),
.B(n_285),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_278),
.B(n_180),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_291),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_183),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_278),
.B(n_187),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_294),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_295),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_318),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_296),
.Y(n_380)
);

AOI221xp5_ASAP7_75t_SL g381 ( 
.A1(n_329),
.A2(n_202),
.B1(n_201),
.B2(n_198),
.C(n_182),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_302),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_284),
.B(n_195),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_302),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_307),
.B(n_258),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_315),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_316),
.B(n_87),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_291),
.B(n_28),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_29),
.Y(n_390)
);

OR2x6_ASAP7_75t_L g391 ( 
.A(n_291),
.B(n_31),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_316),
.B(n_32),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_299),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_387),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_381),
.A2(n_334),
.B(n_342),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_335),
.A2(n_312),
.B(n_313),
.C(n_311),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_328),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_349),
.A2(n_370),
.B(n_348),
.Y(n_398)
);

AOI21x1_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_312),
.B(n_313),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_328),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

AO21x1_ASAP7_75t_L g403 ( 
.A1(n_390),
.A2(n_308),
.B(n_310),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_344),
.B(n_328),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_344),
.A2(n_311),
.B1(n_327),
.B2(n_331),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_336),
.A2(n_328),
.B1(n_331),
.B2(n_327),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_387),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_353),
.B(n_343),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_385),
.A2(n_376),
.B(n_373),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

A2O1A1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_347),
.A2(n_305),
.B(n_304),
.C(n_300),
.Y(n_414)
);

BUFx8_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_47),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

O2A1O1Ixp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_275),
.B(n_287),
.C(n_286),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_374),
.A2(n_269),
.B1(n_283),
.B2(n_282),
.Y(n_421)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_391),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_367),
.A2(n_269),
.B(n_283),
.Y(n_424)
);

BUFx12f_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_55),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_351),
.B(n_56),
.Y(n_427)
);

INVx11_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

AND2x4_ASAP7_75t_SL g430 ( 
.A(n_374),
.B(n_276),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_374),
.B(n_69),
.Y(n_431)
);

BUFx12f_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_377),
.B(n_378),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_380),
.A2(n_266),
.B(n_290),
.C(n_76),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_382),
.A2(n_70),
.B(n_74),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_80),
.B(n_82),
.Y(n_437)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_350),
.B(n_83),
.C(n_84),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_356),
.A2(n_102),
.B(n_103),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_357),
.A2(n_106),
.B(n_107),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_422),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_413),
.B(n_366),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_395),
.A2(n_363),
.B(n_365),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_361),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_412),
.A2(n_372),
.B(n_364),
.C(n_354),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_111),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_428),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_416),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_393),
.Y(n_454)
);

AO31x2_ASAP7_75t_L g455 ( 
.A1(n_396),
.A2(n_435),
.A3(n_439),
.B(n_406),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_434),
.A2(n_405),
.B1(n_433),
.B2(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_397),
.B(n_427),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_438),
.A2(n_426),
.B1(n_417),
.B2(n_432),
.Y(n_458)
);

CKINVDCx6p67_ASAP7_75t_R g459 ( 
.A(n_431),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

AO31x2_ASAP7_75t_L g461 ( 
.A1(n_414),
.A2(n_443),
.A3(n_441),
.B(n_421),
.Y(n_461)
);

BUFx2_ASAP7_75t_SL g462 ( 
.A(n_394),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_407),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_404),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_400),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_436),
.A2(n_437),
.B(n_424),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_442),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_430),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

AO31x2_ASAP7_75t_L g473 ( 
.A1(n_403),
.A2(n_326),
.A3(n_332),
.B(n_329),
.Y(n_473)
);

OAI21xp33_ASAP7_75t_L g474 ( 
.A1(n_413),
.A2(n_289),
.B(n_342),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_410),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_410),
.B(n_359),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_413),
.A2(n_339),
.B1(n_351),
.B2(n_260),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_410),
.B(n_359),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_395),
.A2(n_386),
.B(n_369),
.Y(n_481)
);

OAI21x1_ASAP7_75t_SL g482 ( 
.A1(n_405),
.A2(n_395),
.B(n_403),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_432),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_410),
.B(n_359),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_410),
.B(n_359),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_395),
.A2(n_386),
.B(n_369),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

AO31x2_ASAP7_75t_L g488 ( 
.A1(n_403),
.A2(n_326),
.A3(n_332),
.B(n_329),
.Y(n_488)
);

AO31x2_ASAP7_75t_L g489 ( 
.A1(n_403),
.A2(n_326),
.A3(n_332),
.B(n_329),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_413),
.B(n_359),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_428),
.Y(n_491)
);

AO31x2_ASAP7_75t_L g492 ( 
.A1(n_403),
.A2(n_326),
.A3(n_332),
.B(n_329),
.Y(n_492)
);

NOR2x1_ASAP7_75t_SL g493 ( 
.A(n_425),
.B(n_432),
.Y(n_493)
);

A2O1A1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_412),
.A2(n_395),
.B(n_335),
.C(n_398),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_395),
.A2(n_386),
.B(n_369),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_422),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_416),
.B(n_411),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_416),
.B(n_411),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

AOI21xp33_ASAP7_75t_L g501 ( 
.A1(n_393),
.A2(n_324),
.B(n_346),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_403),
.A2(n_395),
.B(n_399),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_412),
.A2(n_395),
.B(n_335),
.C(n_398),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_412),
.A2(n_395),
.B(n_335),
.C(n_398),
.Y(n_504)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_410),
.B(n_359),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_410),
.B(n_359),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_410),
.B(n_359),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_433),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_413),
.B(n_339),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_410),
.B(n_359),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_491),
.Y(n_515)
);

AND2x4_ASAP7_75t_SL g516 ( 
.A(n_453),
.B(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_466),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_458),
.A2(n_456),
.B1(n_457),
.B2(n_459),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_444),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_474),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_480),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_487),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_447),
.A2(n_454),
.B1(n_501),
.B2(n_478),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_472),
.B(n_510),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_484),
.B(n_485),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_505),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_507),
.Y(n_528)
);

INVx6_ASAP7_75t_L g529 ( 
.A(n_499),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_513),
.Y(n_530)
);

AO31x2_ASAP7_75t_L g531 ( 
.A1(n_486),
.A2(n_495),
.A3(n_446),
.B(n_471),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_458),
.A2(n_511),
.B1(n_510),
.B2(n_468),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_452),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_476),
.Y(n_534)
);

BUFx2_ASAP7_75t_SL g535 ( 
.A(n_483),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

OR3x4_ASAP7_75t_SL g537 ( 
.A(n_483),
.B(n_464),
.C(n_479),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

OAI21x1_ASAP7_75t_SL g539 ( 
.A1(n_463),
.A2(n_465),
.B(n_468),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_499),
.A2(n_470),
.B1(n_496),
.B2(n_512),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_469),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_473),
.Y(n_542)
);

AOI21xp33_ASAP7_75t_L g543 ( 
.A1(n_502),
.A2(n_467),
.B(n_450),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_460),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_462),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_455),
.B(n_489),
.Y(n_547)
);

BUFx2_ASAP7_75t_R g548 ( 
.A(n_445),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_498),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_455),
.B(n_488),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_455),
.B(n_488),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_488),
.A2(n_489),
.B(n_492),
.Y(n_552)
);

AO21x2_ASAP7_75t_L g553 ( 
.A1(n_461),
.A2(n_482),
.B(n_481),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_451),
.B(n_425),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_494),
.A2(n_504),
.B(n_503),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_483),
.B(n_422),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_493),
.B(n_499),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_478),
.A2(n_324),
.B(n_352),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_472),
.B(n_510),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_494),
.A2(n_504),
.B(n_503),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_490),
.B(n_359),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_478),
.A2(n_260),
.B1(n_253),
.B2(n_352),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_468),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_490),
.B(n_359),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_413),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_472),
.B(n_510),
.Y(n_568)
);

O2A1O1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_448),
.A2(n_503),
.B(n_504),
.C(n_494),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_499),
.B(n_394),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_494),
.A2(n_504),
.B(n_503),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_565),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_565),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_518),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_519),
.A2(n_532),
.B1(n_564),
.B2(n_524),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_554),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_522),
.B(n_526),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_528),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_525),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_567),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_519),
.B(n_539),
.Y(n_582)
);

CKINVDCx8_ASAP7_75t_R g583 ( 
.A(n_535),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_542),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_532),
.A2(n_521),
.B1(n_563),
.B2(n_566),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_560),
.B(n_568),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_558),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_514),
.B(n_517),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_559),
.B(n_523),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_546),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

BUFx2_ASAP7_75t_SL g593 ( 
.A(n_555),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_520),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_547),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_550),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_551),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_551),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_569),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_544),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_548),
.A2(n_549),
.B1(n_540),
.B2(n_529),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_556),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_529),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_571),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_606),
.B(n_552),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_606),
.B(n_553),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_573),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_607),
.B(n_553),
.Y(n_614)
);

BUFx4f_ASAP7_75t_SL g615 ( 
.A(n_587),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_578),
.B(n_545),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_580),
.B(n_573),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_543),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_582),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_610),
.B(n_548),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_586),
.B(n_572),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_584),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_584),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_529),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_596),
.B(n_557),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_590),
.B(n_570),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_579),
.B(n_557),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_597),
.B(n_562),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_597),
.B(n_538),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_598),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_611),
.B(n_601),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_612),
.B(n_595),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_615),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_620),
.A2(n_575),
.B1(n_585),
.B2(n_602),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_620),
.A2(n_601),
.B1(n_602),
.B2(n_589),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_599),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_614),
.B(n_595),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_621),
.B(n_600),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_615),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_628),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_622),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_623),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_630),
.B(n_619),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_640),
.B(n_617),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_631),
.B(n_617),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_633),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_638),
.B(n_621),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_638),
.B(n_613),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_630),
.B(n_632),
.Y(n_649)
);

AND2x4_ASAP7_75t_SL g650 ( 
.A(n_641),
.B(n_629),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_630),
.B(n_618),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_618),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_636),
.B(n_613),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_636),
.B(n_628),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_649),
.B(n_641),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_653),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_649),
.B(n_632),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_652),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_651),
.B(n_635),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_647),
.B(n_642),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_637),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_653),
.B(n_637),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_647),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_646),
.A2(n_639),
.B1(n_633),
.B2(n_634),
.Y(n_664)
);

NOR2x1p5_ASAP7_75t_L g665 ( 
.A(n_648),
.B(n_633),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_661),
.B(n_643),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_656),
.B(n_645),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_665),
.A2(n_643),
.B1(n_639),
.B2(n_654),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_664),
.A2(n_605),
.B(n_592),
.C(n_594),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_660),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_661),
.B(n_643),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_655),
.Y(n_672)
);

AOI32xp33_ASAP7_75t_L g673 ( 
.A1(n_657),
.A2(n_650),
.A3(n_639),
.B1(n_620),
.B2(n_626),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_659),
.B(n_644),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_674),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_663),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_670),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_669),
.A2(n_655),
.B(n_624),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_677),
.B(n_668),
.C(n_673),
.Y(n_679)
);

NOR2x1_ASAP7_75t_L g680 ( 
.A(n_678),
.B(n_668),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_675),
.B(n_666),
.Y(n_681)
);

AOI211xp5_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_591),
.B(n_515),
.C(n_676),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_680),
.B(n_583),
.Y(n_683)
);

NOR2x1_ASAP7_75t_L g684 ( 
.A(n_683),
.B(n_527),
.Y(n_684)
);

NOR2x1_ASAP7_75t_L g685 ( 
.A(n_682),
.B(n_593),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_684),
.B(n_681),
.Y(n_686)
);

NOR2x1_ASAP7_75t_L g687 ( 
.A(n_685),
.B(n_533),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_686),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_687),
.B(n_534),
.C(n_604),
.Y(n_689)
);

XNOR2xp5_ASAP7_75t_L g690 ( 
.A(n_689),
.B(n_593),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_688),
.B(n_667),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_688),
.A2(n_583),
.B1(n_591),
.B2(n_658),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_691),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_692),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_690),
.A2(n_591),
.B1(n_536),
.B2(n_590),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g696 ( 
.A(n_690),
.B(n_603),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_690),
.A2(n_581),
.B(n_608),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_694),
.A2(n_590),
.B1(n_671),
.B2(n_577),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_693),
.B(n_624),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_696),
.B(n_537),
.C(n_608),
.Y(n_700)
);

NAND3xp33_ASAP7_75t_L g701 ( 
.A(n_695),
.B(n_590),
.C(n_627),
.Y(n_701)
);

NAND2xp67_ASAP7_75t_L g702 ( 
.A(n_697),
.B(n_588),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_694),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_694),
.A2(n_590),
.B1(n_627),
.B2(n_625),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_703),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_SL g706 ( 
.A(n_700),
.B(n_616),
.C(n_574),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_698),
.B(n_588),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_699),
.B(n_662),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_705),
.A2(n_704),
.B(n_701),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_707),
.B(n_702),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_709),
.A2(n_706),
.B(n_708),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_711),
.B(n_710),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_712),
.A2(n_576),
.B(n_625),
.C(n_616),
.Y(n_713)
);


endmodule