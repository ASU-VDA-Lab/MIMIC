module fake_jpeg_7908_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_3),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx2_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_16),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_31),
.B1(n_25),
.B2(n_14),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_46),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_28),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_56),
.C(n_1),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_25),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_26),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_34),
.B1(n_28),
.B2(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_0),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_1),
.B(n_2),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_68),
.B(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_32),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_54),
.B1(n_40),
.B2(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_54),
.B1(n_56),
.B2(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_54),
.B1(n_28),
.B2(n_46),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_63),
.B(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_87),
.B(n_70),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_60),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_78),
.C(n_74),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_72),
.C(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_96),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_80),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_83),
.B(n_63),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_76),
.C(n_82),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_100),
.C(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_77),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_61),
.C(n_75),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.A3(n_103),
.B1(n_77),
.B2(n_21),
.C1(n_4),
.C2(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_69),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_104),
.Y(n_105)
);


endmodule