module fake_jpeg_18640_n_91 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_91);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_21),
.A2(n_22),
.B1(n_14),
.B2(n_12),
.Y(n_23)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_18),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_14),
.B1(n_13),
.B2(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_17),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_22),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_17),
.B1(n_9),
.B2(n_13),
.Y(n_38)
);

OAI22x1_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_23),
.B1(n_39),
.B2(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_45),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_29),
.B(n_9),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_47),
.B(n_50),
.Y(n_53)
);

AOI22x1_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_47),
.B1(n_41),
.B2(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_8),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_0),
.B(n_1),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_51),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_16),
.B(n_10),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_30),
.C(n_31),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_60),
.C(n_57),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_57),
.B(n_15),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_55),
.B1(n_22),
.B2(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_11),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_22),
.C(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_70),
.Y(n_75)
);

AOI21x1_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_1),
.B(n_4),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_60),
.C(n_53),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_15),
.C(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_15),
.B2(n_2),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_61),
.B1(n_2),
.B2(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_76),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_64),
.Y(n_80)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_1),
.CI(n_5),
.CON(n_76),
.SN(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_80),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_75),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_76),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.C(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_76),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_71),
.B1(n_81),
.B2(n_7),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_81),
.B(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);


endmodule