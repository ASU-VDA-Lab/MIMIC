module real_aes_7460_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_1), .A2(n_154), .B(n_157), .C(n_160), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_2), .A2(n_180), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g540 ( .A(n_3), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_4), .B(n_203), .Y(n_226) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_5), .A2(n_180), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g154 ( .A(n_6), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g187 ( .A(n_7), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_41), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_8), .B(n_41), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_9), .A2(n_234), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_10), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g472 ( .A(n_11), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_12), .B(n_209), .Y(n_511) );
INVx1_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
INVx1_ASAP7_75t_L g523 ( .A(n_14), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_15), .A2(n_188), .B(n_198), .C(n_201), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_16), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_17), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_18), .B(n_479), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_19), .B(n_180), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_20), .B(n_244), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_21), .A2(n_209), .B(n_210), .C(n_212), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_22), .B(n_203), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_23), .B(n_166), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_24), .A2(n_200), .B(n_201), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_25), .B(n_166), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_26), .Y(n_262) );
INVx1_ASAP7_75t_L g252 ( .A(n_27), .Y(n_252) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_28), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_29), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_30), .B(n_166), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_31), .A2(n_64), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_31), .Y(n_131) );
INVx1_ASAP7_75t_L g239 ( .A(n_32), .Y(n_239) );
INVx1_ASAP7_75t_L g461 ( .A(n_33), .Y(n_461) );
INVx2_ASAP7_75t_L g152 ( .A(n_34), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_35), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_36), .A2(n_209), .B(n_222), .C(n_224), .Y(n_221) );
INVxp67_ASAP7_75t_L g241 ( .A(n_37), .Y(n_241) );
CKINVDCx14_ASAP7_75t_R g220 ( .A(n_38), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_39), .A2(n_157), .B(n_251), .C(n_255), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_40), .A2(n_154), .B(n_157), .C(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g460 ( .A(n_42), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_43), .A2(n_168), .B(n_185), .C(n_186), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_44), .B(n_166), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_45), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_46), .Y(n_236) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_47), .A2(n_449), .B1(n_724), .B2(n_727), .C1(n_728), .C2(n_730), .Y(n_448) );
INVx1_ASAP7_75t_L g207 ( .A(n_48), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_49), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_50), .B(n_180), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_51), .A2(n_157), .B1(n_212), .B2(n_459), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_52), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_53), .Y(n_537) );
CKINVDCx14_ASAP7_75t_R g182 ( .A(n_54), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_55), .A2(n_185), .B(n_224), .C(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_56), .Y(n_503) );
INVx1_ASAP7_75t_L g469 ( .A(n_57), .Y(n_469) );
INVx1_ASAP7_75t_L g155 ( .A(n_58), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_59), .A2(n_77), .B1(n_725), .B2(n_726), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_59), .Y(n_726) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
INVx1_ASAP7_75t_SL g223 ( .A(n_61), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_62), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_63), .B(n_203), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_64), .Y(n_130) );
INVx1_ASAP7_75t_L g265 ( .A(n_65), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_SL g478 ( .A1(n_66), .A2(n_224), .B(n_479), .C(n_480), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_67), .Y(n_481) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_69), .A2(n_180), .B(n_181), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_70), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_71), .A2(n_180), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_72), .Y(n_464) );
INVx1_ASAP7_75t_L g497 ( .A(n_73), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_74), .A2(n_234), .B(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g196 ( .A(n_75), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_76), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_77), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_78), .A2(n_102), .B1(n_115), .B2(n_734), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_79), .A2(n_154), .B(n_157), .C(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_80), .A2(n_180), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g199 ( .A(n_81), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_82), .B(n_240), .Y(n_491) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx1_ASAP7_75t_L g161 ( .A(n_84), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_85), .B(n_479), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_86), .A2(n_154), .B(n_157), .C(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
OR2x2_ASAP7_75t_L g123 ( .A(n_87), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g723 ( .A(n_87), .B(n_125), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_88), .A2(n_157), .B(n_264), .C(n_267), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_89), .B(n_142), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_90), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_91), .A2(n_154), .B(n_157), .C(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_92), .Y(n_515) );
INVx1_ASAP7_75t_L g477 ( .A(n_93), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_94), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_95), .B(n_240), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_96), .B(n_173), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_97), .B(n_173), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g211 ( .A(n_99), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_100), .A2(n_180), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g735 ( .A(n_105), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g125 ( .A(n_110), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g720 ( .A(n_111), .B(n_125), .Y(n_720) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_111), .B(n_124), .Y(n_732) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_447), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g733 ( .A(n_120), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_444), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_123), .Y(n_446) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_132), .B2(n_133), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_132), .A2(n_450), .B1(n_718), .B2(n_721), .Y(n_449) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_133), .A2(n_718), .B1(n_723), .B2(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_399), .Y(n_133) );
NAND5xp2_ASAP7_75t_L g134 ( .A(n_135), .B(n_311), .C(n_349), .D(n_370), .E(n_387), .Y(n_134) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_283), .C(n_304), .Y(n_135) );
OAI221xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_215), .B1(n_246), .B2(n_270), .C(n_274), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_175), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_139), .B(n_272), .Y(n_291) );
OR2x2_ASAP7_75t_L g318 ( .A(n_139), .B(n_192), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_139), .B(n_192), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_139), .B(n_178), .Y(n_346) );
AND2x2_ASAP7_75t_L g384 ( .A(n_139), .B(n_348), .Y(n_384) );
AND2x2_ASAP7_75t_L g413 ( .A(n_139), .B(n_323), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_139), .B(n_295), .Y(n_430) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g310 ( .A(n_140), .B(n_191), .Y(n_310) );
BUFx3_ASAP7_75t_L g335 ( .A(n_140), .Y(n_335) );
AND2x2_ASAP7_75t_L g364 ( .A(n_140), .B(n_192), .Y(n_364) );
AND3x2_ASAP7_75t_L g377 ( .A(n_140), .B(n_378), .C(n_379), .Y(n_377) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_147), .B(n_170), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_141), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_141), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_141), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_142), .A2(n_179), .B(n_190), .Y(n_178) );
INVx2_ASAP7_75t_L g245 ( .A(n_142), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_142), .A2(n_149), .B(n_249), .C(n_250), .Y(n_248) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_142), .A2(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_L g174 ( .A(n_143), .B(n_144), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_156), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_149), .A2(n_262), .B(n_263), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_149), .A2(n_189), .B1(n_458), .B2(n_462), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_149), .A2(n_497), .B(n_498), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_149), .A2(n_537), .B(n_538), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
AND2x4_ASAP7_75t_L g180 ( .A(n_150), .B(n_154), .Y(n_180) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g242 ( .A(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx1_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
INVx1_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
INVx3_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
INVx1_ASAP7_75t_L g479 ( .A(n_153), .Y(n_479) );
INVx4_ASAP7_75t_SL g189 ( .A(n_154), .Y(n_189) );
BUFx3_ASAP7_75t_L g255 ( .A(n_154), .Y(n_255) );
INVx5_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx3_ASAP7_75t_L g169 ( .A(n_158), .Y(n_169) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_165), .C(n_167), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_162), .A2(n_167), .B(n_265), .C(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g459 ( .A1(n_163), .A2(n_164), .B1(n_460), .B2(n_461), .Y(n_459) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx4_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
INVx2_ASAP7_75t_L g185 ( .A(n_166), .Y(n_185) );
INVx4_ASAP7_75t_L g209 ( .A(n_166), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_167), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_167), .A2(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g201 ( .A(n_169), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVx3_ASAP7_75t_L g203 ( .A(n_172), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_172), .B(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_172), .A2(n_261), .B(n_268), .Y(n_260) );
NOR2xp33_ASAP7_75t_SL g493 ( .A(n_172), .B(n_494), .Y(n_493) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_173), .Y(n_193) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_173), .A2(n_475), .B(n_482), .Y(n_474) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
INVx1_ASAP7_75t_L g300 ( .A(n_175), .Y(n_300) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_191), .Y(n_175) );
AOI32xp33_ASAP7_75t_L g355 ( .A1(n_176), .A2(n_307), .A3(n_356), .B1(n_359), .B2(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g282 ( .A(n_177), .B(n_191), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_177), .B(n_310), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_177), .B(n_332), .Y(n_360) );
OR2x2_ASAP7_75t_L g366 ( .A(n_177), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_177), .B(n_321), .Y(n_391) );
OR2x2_ASAP7_75t_L g409 ( .A(n_177), .B(n_228), .Y(n_409) );
BUFx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g273 ( .A(n_178), .B(n_204), .Y(n_273) );
INVx2_ASAP7_75t_L g295 ( .A(n_178), .Y(n_295) );
OR2x2_ASAP7_75t_L g317 ( .A(n_178), .B(n_204), .Y(n_317) );
AND2x2_ASAP7_75t_L g322 ( .A(n_178), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_178), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_178), .B(n_272), .Y(n_378) );
BUFx2_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_189), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_183), .A2(n_189), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_SL g206 ( .A1(n_183), .A2(n_189), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_183), .A2(n_189), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_183), .A2(n_189), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_183), .A2(n_189), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_183), .A2(n_189), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_183), .A2(n_189), .B(n_520), .C(n_521), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx5_ASAP7_75t_L g240 ( .A(n_188), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_188), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_188), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
INVx1_ASAP7_75t_SL g429 ( .A(n_191), .Y(n_429) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_204), .Y(n_191) );
INVx1_ASAP7_75t_SL g272 ( .A(n_192), .Y(n_272) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_192), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_192), .B(n_358), .Y(n_357) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_192), .B(n_295), .C(n_413), .Y(n_424) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_202), .Y(n_192) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_193), .A2(n_205), .B(n_214), .Y(n_204) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_193), .A2(n_218), .B(n_226), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_200), .B(n_211), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_200), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_200), .B(n_523), .Y(n_522) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_203), .A2(n_467), .B(n_473), .Y(n_466) );
INVx2_ASAP7_75t_L g323 ( .A(n_204), .Y(n_323) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_204), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_209), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g542 ( .A(n_212), .Y(n_542) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_227), .Y(n_215) );
INVx1_ASAP7_75t_L g359 ( .A(n_216), .Y(n_359) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g277 ( .A(n_217), .B(n_259), .Y(n_277) );
INVx2_ASAP7_75t_L g294 ( .A(n_217), .Y(n_294) );
AND2x2_ASAP7_75t_L g299 ( .A(n_217), .B(n_260), .Y(n_299) );
AND2x2_ASAP7_75t_L g314 ( .A(n_217), .B(n_247), .Y(n_314) );
AND2x2_ASAP7_75t_L g326 ( .A(n_217), .B(n_298), .Y(n_326) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_225), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_227), .B(n_342), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_227), .B(n_299), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_227), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_227), .B(n_293), .Y(n_421) );
BUFx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g258 ( .A(n_228), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_228), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g303 ( .A(n_228), .B(n_247), .Y(n_303) );
AND2x2_ASAP7_75t_L g329 ( .A(n_228), .B(n_259), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_228), .B(n_369), .Y(n_368) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_233), .B(n_243), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_230), .A2(n_288), .B(n_289), .Y(n_287) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_230), .A2(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI21xp5_ASAP7_75t_SL g487 ( .A1(n_231), .A2(n_488), .B(n_489), .Y(n_487) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_232), .A2(n_457), .B(n_463), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_232), .B(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_232), .A2(n_536), .B(n_543), .Y(n_535) );
INVx1_ASAP7_75t_L g288 ( .A(n_233), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_238), .B(n_242), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_240), .A2(n_252), .B(n_253), .C(n_254), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_240), .A2(n_540), .B(n_541), .C(n_542), .Y(n_539) );
INVx2_ASAP7_75t_L g254 ( .A(n_242), .Y(n_254) );
INVx1_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_245), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_245), .A2(n_507), .B(n_514), .Y(n_506) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_258), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_247), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g293 ( .A(n_247), .B(n_294), .Y(n_293) );
INVx3_ASAP7_75t_SL g298 ( .A(n_247), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_247), .B(n_285), .Y(n_351) );
OR2x2_ASAP7_75t_L g361 ( .A(n_247), .B(n_287), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_247), .B(n_329), .Y(n_389) );
OR2x2_ASAP7_75t_L g419 ( .A(n_247), .B(n_259), .Y(n_419) );
AND2x2_ASAP7_75t_L g423 ( .A(n_247), .B(n_260), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_247), .B(n_299), .Y(n_436) );
AND2x2_ASAP7_75t_L g443 ( .A(n_247), .B(n_325), .Y(n_443) );
OR2x6_ASAP7_75t_L g247 ( .A(n_248), .B(n_256), .Y(n_247) );
INVx1_ASAP7_75t_SL g386 ( .A(n_258), .Y(n_386) );
AND2x2_ASAP7_75t_L g325 ( .A(n_259), .B(n_287), .Y(n_325) );
AND2x2_ASAP7_75t_L g339 ( .A(n_259), .B(n_294), .Y(n_339) );
AND2x2_ASAP7_75t_L g342 ( .A(n_259), .B(n_298), .Y(n_342) );
INVx1_ASAP7_75t_L g369 ( .A(n_259), .Y(n_369) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g281 ( .A(n_260), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_271), .A2(n_317), .B(n_441), .C(n_442), .Y(n_440) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g347 ( .A(n_272), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_273), .B(n_290), .Y(n_305) );
AND2x2_ASAP7_75t_L g331 ( .A(n_273), .B(n_332), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_278), .B(n_282), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_276), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_277), .B(n_298), .Y(n_343) );
AND2x2_ASAP7_75t_L g434 ( .A(n_277), .B(n_285), .Y(n_434) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g307 ( .A(n_281), .B(n_294), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_281), .B(n_292), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_291), .A3(n_292), .B1(n_295), .B2(n_296), .C1(n_300), .C2(n_301), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x2_ASAP7_75t_L g395 ( .A(n_285), .B(n_307), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_285), .B(n_359), .Y(n_441) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g338 ( .A(n_287), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g404 ( .A(n_291), .B(n_317), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_292), .B(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_293), .B(n_325), .Y(n_382) );
AND2x2_ASAP7_75t_L g328 ( .A(n_294), .B(n_298), .Y(n_328) );
AND2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_295), .A2(n_374), .B(n_434), .C(n_435), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_296), .A2(n_309), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_298), .B(n_325), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_298), .B(n_339), .Y(n_371) );
AND2x2_ASAP7_75t_L g405 ( .A(n_298), .B(n_307), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_299), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_SL g415 ( .A(n_299), .Y(n_415) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_303), .A2(n_331), .B1(n_333), .B2(n_338), .Y(n_330) );
OAI22xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_306), .B1(n_308), .B2(n_309), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_305), .A2(n_341), .B1(n_343), .B2(n_344), .Y(n_340) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_310), .A2(n_412), .B1(n_414), .B2(n_416), .C(n_420), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B(n_319), .C(n_340), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OR2x2_ASAP7_75t_L g381 ( .A(n_317), .B(n_334), .Y(n_381) );
INVx1_ASAP7_75t_L g432 ( .A(n_317), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_318), .A2(n_320), .B1(n_324), .B2(n_327), .C(n_330), .Y(n_319) );
INVx2_ASAP7_75t_SL g374 ( .A(n_318), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g439 ( .A(n_321), .Y(n_439) );
AND2x2_ASAP7_75t_L g363 ( .A(n_322), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g410 ( .A(n_326), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_334), .B(n_436), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_338), .A2(n_350), .B(n_352), .C(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g427 ( .A(n_341), .Y(n_427) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_345), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx2_ASAP7_75t_L g358 ( .A(n_348), .Y(n_358) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI222xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_361), .B1(n_362), .B2(n_365), .C1(n_366), .C2(n_368), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g394 ( .A(n_358), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_361), .B(n_415), .Y(n_414) );
NAND2xp33_ASAP7_75t_SL g392 ( .A(n_362), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g367 ( .A(n_364), .Y(n_367) );
AND2x2_ASAP7_75t_L g431 ( .A(n_364), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g397 ( .A(n_367), .B(n_394), .Y(n_397) );
INVx1_ASAP7_75t_L g426 ( .A(n_368), .Y(n_426) );
AOI211xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B(n_375), .C(n_380), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_374), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_377), .A2(n_405), .A3(n_410), .B1(n_426), .B2(n_427), .C1(n_428), .C2(n_431), .Y(n_425) );
AND2x2_ASAP7_75t_L g412 ( .A(n_378), .B(n_413), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_383), .B2(n_385), .Y(n_380) );
INVxp33_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B1(n_392), .B2(n_395), .C(n_396), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND5xp2_ASAP7_75t_L g399 ( .A(n_400), .B(n_411), .C(n_425), .D(n_433), .E(n_437), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_405), .B(n_406), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp33_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_413), .A2(n_438), .B(n_439), .C(n_440), .Y(n_437) );
AOI31xp33_ASAP7_75t_L g420 ( .A1(n_415), .A2(n_421), .A3(n_422), .B(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g438 ( .A(n_436), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_444), .B(n_448), .C(n_733), .Y(n_447) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g729 ( .A(n_450), .Y(n_729) );
AND3x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_643), .C(n_692), .Y(n_450) );
NOR3xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_550), .C(n_588), .Y(n_451) );
OAI222xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_483), .B1(n_525), .B2(n_531), .C1(n_545), .C2(n_548), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_465), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_454), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_454), .B(n_593), .Y(n_684) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g561 ( .A(n_455), .B(n_474), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_455), .B(n_466), .Y(n_569) );
AND2x2_ASAP7_75t_L g604 ( .A(n_455), .B(n_581), .Y(n_604) );
OR2x2_ASAP7_75t_L g628 ( .A(n_455), .B(n_466), .Y(n_628) );
OR2x2_ASAP7_75t_L g636 ( .A(n_455), .B(n_535), .Y(n_636) );
AND2x2_ASAP7_75t_L g639 ( .A(n_455), .B(n_474), .Y(n_639) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g533 ( .A(n_456), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g547 ( .A(n_456), .B(n_474), .Y(n_547) );
AND2x2_ASAP7_75t_L g597 ( .A(n_456), .B(n_535), .Y(n_597) );
AND2x2_ASAP7_75t_L g610 ( .A(n_456), .B(n_466), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_456), .B(n_696), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_465), .A2(n_636), .B(n_637), .C(n_640), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_465), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_465), .B(n_580), .Y(n_702) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_474), .Y(n_465) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_466), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g560 ( .A(n_466), .Y(n_560) );
AND2x2_ASAP7_75t_L g587 ( .A(n_466), .B(n_581), .Y(n_587) );
INVx1_ASAP7_75t_SL g595 ( .A(n_466), .Y(n_595) );
AND2x2_ASAP7_75t_L g618 ( .A(n_466), .B(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g696 ( .A(n_466), .Y(n_696) );
BUFx2_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
INVx1_ASAP7_75t_L g594 ( .A(n_474), .Y(n_594) );
INVx3_ASAP7_75t_L g619 ( .A(n_474), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_483), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_504), .Y(n_483) );
INVx1_ASAP7_75t_L g615 ( .A(n_484), .Y(n_615) );
OAI32xp33_ASAP7_75t_L g621 ( .A1(n_484), .A2(n_560), .A3(n_622), .B1(n_623), .B2(n_624), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_484), .A2(n_626), .B1(n_629), .B2(n_634), .Y(n_625) );
INVx4_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g563 ( .A(n_485), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g641 ( .A(n_485), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g711 ( .A(n_485), .B(n_657), .Y(n_711) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
AND2x2_ASAP7_75t_L g526 ( .A(n_486), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
INVx1_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
OR2x2_ASAP7_75t_L g583 ( .A(n_486), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g590 ( .A(n_486), .B(n_564), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_486), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g611 ( .A(n_486), .B(n_529), .Y(n_611) );
INVx3_ASAP7_75t_L g633 ( .A(n_486), .Y(n_633) );
AND2x2_ASAP7_75t_L g658 ( .A(n_486), .B(n_530), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_486), .B(n_623), .Y(n_706) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx2_ASAP7_75t_L g530 ( .A(n_495), .Y(n_530) );
AND2x2_ASAP7_75t_L g662 ( .A(n_495), .B(n_505), .Y(n_662) );
INVx2_ASAP7_75t_L g704 ( .A(n_504), .Y(n_704) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_516), .Y(n_504) );
INVx1_ASAP7_75t_L g549 ( .A(n_505), .Y(n_549) );
AND2x2_ASAP7_75t_L g576 ( .A(n_505), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_505), .B(n_530), .Y(n_584) );
AND2x2_ASAP7_75t_L g642 ( .A(n_505), .B(n_565), .Y(n_642) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g528 ( .A(n_506), .Y(n_528) );
AND2x2_ASAP7_75t_L g555 ( .A(n_506), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g564 ( .A(n_506), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_506), .B(n_530), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_516), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_516), .B(n_530), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_516), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g657 ( .A(n_516), .Y(n_657) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g529 ( .A(n_517), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_525), .A2(n_535), .B1(n_694), .B2(n_697), .Y(n_693) );
INVx1_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_527), .A2(n_638), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_528), .B(n_633), .Y(n_650) );
INVx1_ASAP7_75t_L g675 ( .A(n_528), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_529), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_555), .Y(n_602) );
INVx2_ASAP7_75t_L g558 ( .A(n_530), .Y(n_558) );
INVx1_ASAP7_75t_L g608 ( .A(n_530), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_531), .A2(n_683), .B1(n_700), .B2(n_703), .C(n_705), .Y(n_699) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g570 ( .A(n_532), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_532), .B(n_581), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_533), .B(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g624 ( .A(n_533), .B(n_570), .Y(n_624) );
INVx3_ASAP7_75t_SL g665 ( .A(n_533), .Y(n_665) );
AND2x2_ASAP7_75t_L g609 ( .A(n_534), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g638 ( .A(n_534), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_534), .B(n_547), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_534), .B(n_593), .Y(n_679) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
OAI322xp33_ASAP7_75t_L g676 ( .A1(n_535), .A2(n_607), .A3(n_629), .B1(n_677), .B2(n_679), .C1(n_680), .C2(n_681), .Y(n_676) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_546), .A2(n_549), .B(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_SL g626 ( .A(n_547), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g648 ( .A(n_547), .B(n_560), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_547), .B(n_587), .Y(n_663) );
INVxp67_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g620 ( .A1(n_549), .A2(n_621), .B(n_625), .C(n_635), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_559), .B1(n_562), .B2(n_566), .C(n_571), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g574 ( .A(n_558), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g691 ( .A(n_558), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_559), .A2(n_708), .B1(n_713), .B2(n_714), .C(n_716), .Y(n_707) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_560), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g607 ( .A(n_560), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_560), .B(n_638), .Y(n_645) );
AND2x2_ASAP7_75t_L g687 ( .A(n_560), .B(n_665), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_561), .B(n_586), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_561), .A2(n_573), .B1(n_683), .B2(n_684), .Y(n_682) );
OR2x2_ASAP7_75t_L g713 ( .A(n_561), .B(n_581), .Y(n_713) );
CKINVDCx16_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g690 ( .A(n_564), .Y(n_690) );
AND2x2_ASAP7_75t_L g715 ( .A(n_564), .B(n_658), .Y(n_715) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_SL g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g579 ( .A(n_569), .B(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_578), .B1(n_582), .B2(n_585), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx1_ASAP7_75t_L g646 ( .A(n_574), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_574), .B(n_614), .Y(n_681) );
AOI322xp5_ASAP7_75t_L g605 ( .A1(n_576), .A2(n_606), .A3(n_608), .B1(n_609), .B2(n_611), .C1(n_612), .C2(n_616), .Y(n_605) );
INVxp67_ASAP7_75t_L g599 ( .A(n_577), .Y(n_599) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_579), .A2(n_584), .B1(n_601), .B2(n_603), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_580), .B(n_593), .Y(n_680) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_581), .B(n_619), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_581), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g677 ( .A(n_583), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g588 ( .A(n_589), .B(n_605), .C(n_620), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_596), .B2(n_598), .C(n_600), .Y(n_589) );
AND2x2_ASAP7_75t_L g596 ( .A(n_592), .B(n_597), .Y(n_596) );
INVx3_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g606 ( .A(n_597), .B(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_599), .Y(n_678) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_604), .B(n_618), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_607), .B(n_665), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_608), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g683 ( .A(n_611), .Y(n_683) );
AND2x2_ASAP7_75t_L g698 ( .A(n_611), .B(n_675), .Y(n_698) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g692 ( .A1(n_622), .A2(n_693), .B(n_699), .C(n_707), .Y(n_692) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g661 ( .A(n_632), .B(n_662), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g703 ( .A(n_633), .B(n_704), .Y(n_703) );
CKINVDCx16_ASAP7_75t_R g673 ( .A(n_636), .Y(n_673) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g668 ( .A(n_642), .Y(n_668) );
AND2x2_ASAP7_75t_L g672 ( .A(n_642), .B(n_658), .Y(n_672) );
NOR5xp2_ASAP7_75t_L g643 ( .A(n_644), .B(n_659), .C(n_676), .D(n_682), .E(n_685), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_649), .C(n_651), .Y(n_644) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_648), .B(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g674 ( .A(n_658), .B(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_663), .B1(n_664), .B2(n_666), .C(n_669), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g712 ( .A(n_672), .Y(n_712) );
AOI211xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_688), .B(n_690), .C(n_691), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx14_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx14_ASAP7_75t_R g727 ( .A(n_724), .Y(n_727) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
endmodule