module fake_jpeg_14469_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_74),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_18),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_101),
.Y(n_110)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_80),
.Y(n_152)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_102),
.Y(n_134)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_88),
.Y(n_116)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_42),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_105),
.B(n_112),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_31),
.B1(n_41),
.B2(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_109),
.A2(n_113),
.B1(n_117),
.B2(n_119),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_43),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_31),
.B1(n_41),
.B2(n_50),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_50),
.B1(n_34),
.B2(n_37),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_65),
.A2(n_50),
.B1(n_34),
.B2(n_37),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_87),
.B1(n_95),
.B2(n_64),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_128),
.A2(n_131),
.B1(n_137),
.B2(n_148),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_55),
.A2(n_50),
.B1(n_34),
.B2(n_37),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_34),
.B1(n_37),
.B2(n_36),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_43),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_144),
.B(n_159),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_29),
.B1(n_32),
.B2(n_40),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_161),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_56),
.A2(n_29),
.B1(n_40),
.B2(n_45),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_93),
.B(n_45),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_62),
.B(n_44),
.C(n_48),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_47),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_98),
.B(n_42),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_166),
.B(n_1),
.Y(n_222)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_167),
.Y(n_269)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_169),
.Y(n_280)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_183),
.Y(n_236)
);

AOI32xp33_ASAP7_75t_L g175 ( 
.A1(n_114),
.A2(n_81),
.A3(n_80),
.B1(n_58),
.B2(n_42),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_175),
.A2(n_189),
.B(n_204),
.Y(n_253)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_185),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_116),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_178),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_51),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_126),
.B(n_51),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_33),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_199),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_139),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_47),
.B1(n_68),
.B2(n_84),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_221),
.B1(n_162),
.B2(n_7),
.Y(n_267)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_206),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_51),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_209),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_48),
.B(n_46),
.C(n_33),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_111),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_48),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_123),
.B(n_115),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_113),
.A2(n_91),
.B1(n_70),
.B2(n_83),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_225),
.B1(n_152),
.B2(n_119),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_106),
.B(n_46),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_227),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_107),
.A2(n_46),
.B1(n_33),
.B2(n_42),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_163),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_219),
.Y(n_265)
);

NOR2x1_ASAP7_75t_R g218 ( 
.A(n_109),
.B(n_42),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_117),
.Y(n_228)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_222),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_131),
.A2(n_82),
.B1(n_77),
.B2(n_3),
.Y(n_221)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_137),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_107),
.A2(n_88),
.B1(n_2),
.B2(n_5),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_228),
.B(n_223),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_179),
.B(n_135),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_229),
.B(n_241),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_231),
.A2(n_248),
.B1(n_264),
.B2(n_275),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_177),
.A2(n_142),
.B1(n_141),
.B2(n_133),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_237),
.A2(n_173),
.B1(n_172),
.B2(n_194),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_204),
.B(n_202),
.C(n_178),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_240),
.A2(n_246),
.B(n_262),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_196),
.B(n_141),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_163),
.B(n_116),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_184),
.B(n_142),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_247),
.B(n_259),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_128),
.B1(n_140),
.B2(n_153),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_180),
.B(n_157),
.C(n_153),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_173),
.C(n_206),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_209),
.B(n_133),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_185),
.A2(n_88),
.B(n_5),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_221),
.A2(n_162),
.B1(n_154),
.B2(n_8),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_169),
.B1(n_191),
.B2(n_195),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_213),
.B(n_181),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_170),
.B(n_1),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_218),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_203),
.B(n_8),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_9),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_207),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_248),
.B1(n_231),
.B2(n_272),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_245),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_281),
.Y(n_366)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_238),
.B(n_190),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_284),
.B(n_312),
.Y(n_338)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_286),
.B(n_307),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_197),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_298),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_288),
.Y(n_343)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_192),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_296),
.Y(n_370)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_299),
.A2(n_301),
.B1(n_317),
.B2(n_324),
.Y(n_356)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_228),
.A2(n_252),
.B1(n_267),
.B2(n_240),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_236),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_314),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_233),
.B(n_187),
.C(n_220),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_304),
.C(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_229),
.C(n_247),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_199),
.B(n_182),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_305),
.A2(n_306),
.B(n_323),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_238),
.A2(n_224),
.B(n_219),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_242),
.B(n_168),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_309),
.B1(n_321),
.B2(n_269),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_258),
.A2(n_241),
.B1(n_259),
.B2(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_315),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_176),
.C(n_171),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_313),
.B(n_296),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_246),
.A2(n_253),
.B(n_262),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_328),
.B(n_255),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_251),
.A2(n_193),
.B1(n_201),
.B2(n_227),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_270),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_319),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_260),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_276),
.A2(n_10),
.B(n_11),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_320),
.A2(n_255),
.B1(n_263),
.B2(n_269),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_234),
.A2(n_188),
.B1(n_167),
.B2(n_12),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_266),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_266),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_326),
.Y(n_344)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_13),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_329),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_257),
.A2(n_13),
.B(n_14),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_254),
.C(n_257),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_349),
.C(n_355),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_301),
.A2(n_280),
.B1(n_250),
.B2(n_261),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_346),
.B1(n_363),
.B2(n_371),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_339),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_313),
.B(n_316),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_340),
.A2(n_342),
.B(n_358),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_290),
.A2(n_313),
.B(n_305),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_280),
.B1(n_261),
.B2(n_273),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_357),
.B1(n_367),
.B2(n_283),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_277),
.C(n_256),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_300),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_282),
.B(n_287),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_359),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_277),
.C(n_256),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_295),
.A2(n_243),
.B1(n_249),
.B2(n_273),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_263),
.B(n_249),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_263),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_314),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_369),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_328),
.A2(n_289),
.B(n_322),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_299),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_14),
.C(n_16),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_323),
.C(n_324),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_295),
.A2(n_14),
.B1(n_16),
.B2(n_309),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_329),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_317),
.A2(n_288),
.B1(n_284),
.B2(n_302),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_347),
.B(n_312),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_375),
.B(n_377),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_394),
.C(n_395),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_366),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_321),
.B(n_319),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_379),
.A2(n_401),
.B(n_403),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_366),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_384),
.Y(n_418)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_298),
.B1(n_293),
.B2(n_285),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_383),
.A2(n_386),
.B1(n_398),
.B2(n_404),
.Y(n_426)
);

OAI22x1_ASAP7_75t_SL g386 ( 
.A1(n_348),
.A2(n_319),
.B1(n_294),
.B2(n_297),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_341),
.B(n_292),
.Y(n_390)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_344),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_393),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_281),
.C(n_310),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_325),
.Y(n_395)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_397),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_338),
.B(n_286),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_409),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_400),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_343),
.A2(n_326),
.B1(n_336),
.B2(n_356),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_343),
.A2(n_360),
.B1(n_334),
.B2(n_346),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_331),
.A2(n_368),
.B1(n_339),
.B2(n_355),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_357),
.B1(n_338),
.B2(n_369),
.Y(n_407)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_331),
.A2(n_368),
.B1(n_370),
.B2(n_362),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_333),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_433),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_342),
.B(n_340),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_413),
.A2(n_420),
.B(n_430),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_390),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_416),
.B(n_388),
.Y(n_448)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_374),
.A2(n_353),
.B(n_345),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_333),
.C(n_349),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_424),
.C(n_431),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_368),
.C(n_354),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_399),
.A2(n_365),
.B(n_332),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_376),
.C(n_409),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_350),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_382),
.B(n_400),
.Y(n_434)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_365),
.Y(n_436)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_436),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_391),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_439),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_427),
.B(n_396),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_442),
.B(n_455),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_441),
.A2(n_379),
.B1(n_386),
.B2(n_387),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_444),
.A2(n_464),
.B1(n_440),
.B2(n_435),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_417),
.Y(n_446)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_441),
.A2(n_401),
.B1(n_404),
.B2(n_373),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_423),
.B1(n_412),
.B2(n_410),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_388),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_461),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_411),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_468),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_431),
.B(n_396),
.Y(n_453)
);

XNOR2x1_ASAP7_75t_L g489 ( 
.A(n_453),
.B(n_330),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_385),
.C(n_383),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_457),
.C(n_460),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_418),
.B(n_384),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_385),
.C(n_389),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_423),
.A2(n_373),
.B1(n_425),
.B2(n_439),
.Y(n_459)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_381),
.C(n_387),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_379),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_426),
.A2(n_408),
.B1(n_406),
.B2(n_337),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_465),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_364),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_434),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_330),
.C(n_332),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_430),
.C(n_438),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_410),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_445),
.A2(n_413),
.B(n_437),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_476),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_471),
.A2(n_464),
.B1(n_463),
.B2(n_445),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_414),
.Y(n_475)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_475),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_467),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_437),
.C(n_412),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_480),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_420),
.C(n_414),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_419),
.C(n_429),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_483),
.C(n_484),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_419),
.C(n_429),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_440),
.C(n_438),
.Y(n_484)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_444),
.A2(n_432),
.B1(n_435),
.B2(n_422),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_361),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_432),
.B(n_363),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_466),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_461),
.Y(n_499)
);

AOI21xp33_ASAP7_75t_L g492 ( 
.A1(n_486),
.A2(n_475),
.B(n_469),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_492),
.B(n_476),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_499),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_460),
.Y(n_495)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_456),
.C(n_453),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_500),
.Y(n_517)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_462),
.B1(n_446),
.B2(n_443),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_501),
.A2(n_472),
.B1(n_470),
.B2(n_488),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_480),
.A2(n_456),
.B(n_452),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_503),
.B(n_504),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_361),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_489),
.B(n_337),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_506),
.B(n_473),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_487),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_474),
.B(n_482),
.C(n_473),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_508),
.B(n_483),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_502),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_510),
.B(n_520),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_494),
.Y(n_529)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_490),
.B(n_471),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g531 ( 
.A1(n_513),
.A2(n_523),
.B(n_507),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_515),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_519),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_493),
.B(n_504),
.C(n_508),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_479),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_491),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_505),
.A2(n_488),
.B(n_472),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_495),
.C(n_517),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_532),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_529),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_497),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_509),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_513),
.C(n_522),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_477),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_516),
.B(n_498),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_533),
.B(n_521),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_530),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_536),
.A2(n_526),
.B(n_528),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_539),
.B(n_541),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_523),
.Y(n_541)
);

O2A1O1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_542),
.A2(n_543),
.B(n_544),
.C(n_515),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_537),
.A2(n_534),
.B(n_529),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_546),
.A2(n_547),
.B(n_531),
.Y(n_548)
);

NAND4xp25_ASAP7_75t_SL g547 ( 
.A(n_545),
.B(n_540),
.C(n_538),
.D(n_536),
.Y(n_547)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_548),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_525),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_485),
.C(n_499),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_506),
.Y(n_552)
);


endmodule