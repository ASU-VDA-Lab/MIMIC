module fake_jpeg_19953_n_309 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_20),
.B1(n_14),
.B2(n_18),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_24),
.B2(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_54),
.B1(n_30),
.B2(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_35),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_47),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_46),
.B1(n_37),
.B2(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_77),
.B1(n_60),
.B2(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_37),
.B1(n_30),
.B2(n_24),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_41),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_85),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_83),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_37),
.B1(n_45),
.B2(n_26),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_38),
.B(n_37),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_57),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_76),
.C(n_73),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_71),
.C(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_52),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_62),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_45),
.B1(n_30),
.B2(n_44),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_38),
.B1(n_61),
.B2(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_103),
.B1(n_109),
.B2(n_82),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_27),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_117),
.C(n_79),
.Y(n_138)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_71),
.B1(n_70),
.B2(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_100),
.C(n_117),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_116),
.B(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_71),
.B1(n_65),
.B2(n_68),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_98),
.Y(n_122)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_67),
.B(n_35),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_83),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_67),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_34),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_26),
.B1(n_41),
.B2(n_29),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_34),
.B(n_14),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_75),
.B1(n_90),
.B2(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_104),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_132),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_139),
.B1(n_44),
.B2(n_78),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_142),
.B(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_86),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_136),
.Y(n_167)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_150),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_32),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_87),
.B1(n_45),
.B2(n_94),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_140),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_105),
.Y(n_142)
);

CKINVDCx10_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_144),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_55),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_148),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_18),
.C(n_16),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_55),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_44),
.C(n_17),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_181),
.B1(n_143),
.B2(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_138),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_12),
.B(n_15),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_175),
.B(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_152),
.C(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_90),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_90),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_81),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_174),
.B1(n_179),
.B2(n_78),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_42),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_4),
.B(n_10),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_32),
.B(n_24),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_42),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_15),
.B(n_16),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_151),
.B1(n_131),
.B2(n_134),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_189),
.B1(n_206),
.B2(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_192),
.C(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_129),
.B1(n_139),
.B2(n_127),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_135),
.B(n_127),
.C(n_146),
.D(n_141),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_154),
.C(n_164),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_147),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_141),
.C(n_134),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_197),
.B1(n_200),
.B2(n_202),
.Y(n_217)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_143),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_78),
.B1(n_41),
.B2(n_20),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_53),
.C(n_31),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_41),
.B1(n_53),
.B2(n_42),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_165),
.C(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_192),
.C(n_204),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_203),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_23),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_161),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_215),
.C(n_219),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_208),
.B(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_167),
.B1(n_155),
.B2(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_160),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_159),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_177),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_225),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_153),
.B1(n_179),
.B2(n_169),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_177),
.B1(n_164),
.B2(n_181),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_206),
.B1(n_174),
.B2(n_178),
.Y(n_234)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_172),
.C(n_171),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_31),
.C(n_28),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_190),
.B(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_232),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_187),
.B(n_196),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_229),
.B1(n_212),
.B2(n_187),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_222),
.B1(n_211),
.B2(n_221),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_31),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_209),
.B(n_9),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_40),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_209),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_219),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_22),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_22),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_22),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_261),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_236),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_31),
.C(n_28),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_260),
.C(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_28),
.C(n_17),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_22),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_260),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_247),
.C(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_271),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_239),
.C(n_238),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_242),
.B(n_231),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_6),
.B(n_7),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_236),
.C(n_242),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_7),
.B1(n_9),
.B2(n_8),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_245),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_23),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_258),
.B1(n_232),
.B2(n_234),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_23),
.A3(n_5),
.B1(n_6),
.B2(n_4),
.C1(n_17),
.C2(n_13),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_28),
.C(n_11),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_286),
.C(n_265),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_285),
.B1(n_4),
.B2(n_1),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_5),
.B(n_6),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_11),
.C(n_17),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_11),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_264),
.C(n_11),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_0),
.C(n_1),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_297),
.A2(n_1),
.B(n_2),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_2),
.A3(n_3),
.B1(n_13),
.B2(n_17),
.C1(n_286),
.C2(n_281),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_290),
.B1(n_291),
.B2(n_296),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.C(n_304),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_289),
.B(n_287),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_298),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_2),
.B(n_3),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_2),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_3),
.C(n_154),
.Y(n_309)
);


endmodule