module fake_jpeg_8719_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_14),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_52),
.B1(n_61),
.B2(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_55),
.B(n_54),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_20),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_60),
.B1(n_45),
.B2(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_45),
.B1(n_48),
.B2(n_57),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_22),
.B1(n_41),
.B2(n_39),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_87),
.B1(n_91),
.B2(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_97),
.C(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_46),
.C(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_46),
.B1(n_8),
.B2(n_7),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_8),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_95),
.B(n_94),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_107),
.B1(n_105),
.B2(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_103),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_83),
.B1(n_104),
.B2(n_86),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_21),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_106),
.B(n_26),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_96),
.C(n_28),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_25),
.C(n_30),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_31),
.C(n_32),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_34),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);


endmodule