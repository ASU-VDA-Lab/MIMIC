module fake_jpeg_26983_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_20),
.B(n_28),
.C(n_32),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_47),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_28),
.B1(n_27),
.B2(n_18),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_17),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_31),
.B1(n_16),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_69),
.B1(n_34),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_16),
.B1(n_26),
.B2(n_31),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_67),
.B1(n_20),
.B2(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_27),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_16),
.B1(n_26),
.B2(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_22),
.B1(n_21),
.B2(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_16),
.B1(n_26),
.B2(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_34),
.B1(n_24),
.B2(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_74),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_73),
.B(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_103),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_55),
.B1(n_47),
.B2(n_48),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_82),
.Y(n_130)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_22),
.B1(n_17),
.B2(n_19),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_86),
.Y(n_131)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_91),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_18),
.B1(n_32),
.B2(n_21),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_39),
.B1(n_17),
.B2(n_30),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_93),
.A2(n_5),
.B(n_6),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_22),
.B1(n_33),
.B2(n_29),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_46),
.B1(n_49),
.B2(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_17),
.B1(n_30),
.B2(n_19),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_23),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_46),
.A2(n_30),
.B1(n_19),
.B2(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_50),
.B(n_10),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_33),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_56),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_61),
.B1(n_29),
.B2(n_35),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_56),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_119),
.B1(n_129),
.B2(n_132),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_35),
.B(n_23),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_93),
.C(n_83),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_23),
.B(n_1),
.C(n_2),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_82),
.B(n_100),
.C(n_7),
.D(n_6),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_93),
.B1(n_96),
.B2(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_138),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_100),
.B1(n_92),
.B2(n_107),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_154),
.B(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_134),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_146),
.B1(n_151),
.B2(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_144),
.B(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_77),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_148),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_110),
.B1(n_138),
.B2(n_137),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_75),
.B1(n_93),
.B2(n_85),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_150),
.B1(n_110),
.B2(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_88),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_153),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_93),
.B1(n_103),
.B2(n_78),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_106),
.B1(n_109),
.B2(n_96),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_70),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_158),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_82),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_91),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_87),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_81),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_100),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_92),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_116),
.B(n_117),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_186),
.B1(n_189),
.B2(n_196),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_130),
.C(n_123),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_201),
.C(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_136),
.B1(n_139),
.B2(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_139),
.B1(n_119),
.B2(n_117),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_202),
.B(n_157),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_139),
.B1(n_116),
.B2(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_145),
.B(n_14),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_148),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_126),
.C(n_8),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_13),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_123),
.C(n_111),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_126),
.B(n_118),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_111),
.C(n_115),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_209),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_141),
.B(n_153),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_179),
.B(n_177),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_154),
.B(n_146),
.C(n_167),
.D(n_168),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_211),
.B(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_140),
.B1(n_150),
.B2(n_169),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_191),
.B1(n_179),
.B2(n_174),
.Y(n_249)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_171),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_178),
.B1(n_189),
.B2(n_151),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_226),
.B1(n_200),
.B2(n_191),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_183),
.B(n_174),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_161),
.B1(n_142),
.B2(n_155),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_176),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_115),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_231),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_121),
.B(n_71),
.C(n_155),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_193),
.B1(n_195),
.B2(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_216),
.B1(n_211),
.B2(n_192),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_173),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_238),
.A2(n_249),
.B1(n_198),
.B2(n_190),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_242),
.B(n_251),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_183),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_173),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_248),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_252),
.B(n_121),
.Y(n_268)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_177),
.B(n_190),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_231),
.B1(n_207),
.B2(n_220),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_234),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_228),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_228),
.C(n_222),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_248),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_266),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_232),
.C(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_230),
.C(n_223),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_213),
.C(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_249),
.C(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_246),
.B1(n_234),
.B2(n_236),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_271),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_216),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_269),
.B1(n_246),
.B2(n_238),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_266),
.B(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_192),
.B1(n_156),
.B2(n_71),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_162),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_241),
.B1(n_244),
.B2(n_249),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_276),
.B1(n_284),
.B2(n_265),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_283),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_281),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_250),
.B(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_235),
.B1(n_245),
.B2(n_237),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_247),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.C(n_259),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_237),
.C(n_243),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_243),
.B1(n_250),
.B2(n_233),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_281),
.B1(n_278),
.B2(n_285),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_86),
.B1(n_9),
.B2(n_11),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_261),
.C(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_247),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_252),
.C(n_233),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_79),
.C(n_94),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_277),
.B(n_294),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_288),
.B1(n_280),
.B2(n_278),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_306),
.B1(n_298),
.B2(n_297),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_277),
.B(n_8),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_291),
.B(n_9),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_299),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_303),
.A2(n_287),
.B(n_292),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_101),
.C(n_9),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_12),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_11),
.B(n_12),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_315),
.B(n_12),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_316),
.B(n_317),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_310),
.B(n_14),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_15),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_15),
.B(n_5),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);


endmodule