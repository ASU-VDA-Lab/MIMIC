module fake_jpeg_30039_n_423 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_423);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_423;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_0),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_64),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_0),
.CON(n_62),
.SN(n_62)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_39),
.B1(n_38),
.B2(n_20),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_73),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_29),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_74),
.B1(n_28),
.B2(n_19),
.Y(n_117)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_16),
.B1(n_15),
.B2(n_3),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_30),
.B(n_15),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_37),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_32),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_19),
.B1(n_28),
.B2(n_30),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_95),
.B1(n_121),
.B2(n_23),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_91),
.B(n_123),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_75),
.B1(n_72),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_93),
.A2(n_128),
.B1(n_35),
.B2(n_22),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_28),
.B1(n_19),
.B2(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_24),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_93),
.B(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_125),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_39),
.B1(n_38),
.B2(n_20),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_49),
.B(n_37),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_129),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_39),
.B1(n_35),
.B2(n_23),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_33),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_63),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_18),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_46),
.B(n_18),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_17),
.Y(n_150)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_68),
.B1(n_74),
.B2(n_65),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_142),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_155),
.B(n_46),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_69),
.B1(n_71),
.B2(n_79),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_35),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_153),
.C(n_168),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_150),
.Y(n_177)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_162),
.B1(n_165),
.B2(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_84),
.B1(n_83),
.B2(n_78),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_98),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_0),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_23),
.B(n_22),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_22),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_98),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_89),
.B(n_96),
.C(n_103),
.Y(n_168)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_94),
.B(n_2),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_153),
.C(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_171),
.B(n_132),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_110),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_166),
.B1(n_139),
.B2(n_163),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_194),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_200),
.B1(n_210),
.B2(n_211),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_155),
.B(n_141),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_189),
.B(n_174),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_142),
.B1(n_151),
.B2(n_145),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_138),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_163),
.B1(n_92),
.B2(n_88),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_165),
.B1(n_160),
.B2(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_205),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_154),
.B1(n_156),
.B2(n_104),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_188),
.B(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_177),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_213),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_140),
.B1(n_168),
.B2(n_149),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_140),
.B1(n_108),
.B2(n_130),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_229),
.B(n_235),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_219),
.B1(n_165),
.B2(n_190),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_175),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_230),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_144),
.C(n_143),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_153),
.B(n_170),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_174),
.B(n_176),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_213),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_189),
.B(n_181),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_201),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_227),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_199),
.B(n_202),
.C(n_195),
.D(n_196),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_229),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_196),
.B1(n_210),
.B2(n_211),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_253),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_211),
.B1(n_200),
.B2(n_197),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_200),
.B1(n_206),
.B2(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_202),
.B1(n_205),
.B2(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_218),
.B(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_250),
.B(n_254),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_170),
.B1(n_186),
.B2(n_190),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_230),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_161),
.A3(n_167),
.B1(n_146),
.B2(n_193),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_224),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_259),
.B(n_265),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_239),
.B1(n_249),
.B2(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_228),
.C(n_218),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_274),
.C(n_275),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_263),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_243),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_217),
.B(n_223),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_268),
.B(n_270),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_254),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_234),
.B1(n_231),
.B2(n_220),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_241),
.B1(n_252),
.B2(n_226),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_226),
.B(n_193),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_209),
.C(n_192),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_182),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_278),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_243),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_279),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_280),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_240),
.B(n_247),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_284),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_272),
.B1(n_266),
.B2(n_273),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_241),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_295),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_270),
.B(n_259),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_180),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_192),
.C(n_158),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_265),
.C(n_275),
.Y(n_304)
);

A2O1A1O1Ixp25_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_231),
.B(n_220),
.C(n_252),
.D(n_180),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_322),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_307),
.C(n_316),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_294),
.B1(n_284),
.B2(n_288),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_273),
.C(n_258),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_272),
.B1(n_271),
.B2(n_268),
.Y(n_312)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_271),
.B1(n_258),
.B2(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_220),
.C(n_191),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_291),
.B(n_180),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_280),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_320),
.Y(n_346)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_291),
.B(n_198),
.CI(n_180),
.CON(n_320),
.SN(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_198),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_191),
.C(n_157),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_289),
.C(n_297),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_295),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_333),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_310),
.B(n_285),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_328),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_303),
.A2(n_299),
.B1(n_292),
.B2(n_290),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_341),
.Y(n_355)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_301),
.B(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_335),
.C(n_337),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_297),
.C(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_186),
.C(n_162),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_186),
.C(n_87),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_342),
.C(n_344),
.Y(n_357)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_SL g340 ( 
.A(n_302),
.B(n_190),
.C(n_159),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_87),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_169),
.C(n_137),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_309),
.A2(n_159),
.B1(n_130),
.B2(n_108),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_346),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_315),
.B1(n_300),
.B2(n_308),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_354),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_327),
.A2(n_305),
.B(n_320),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_358),
.B(n_361),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_333),
.A2(n_323),
.B1(n_320),
.B2(n_317),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_134),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_2),
.B(n_3),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_115),
.C(n_136),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_360),
.B(n_343),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_324),
.A2(n_2),
.B(n_3),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_367),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_355),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_349),
.A2(n_334),
.B1(n_338),
.B2(n_344),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_370),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_343),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_326),
.B1(n_324),
.B2(n_337),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_373),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_359),
.A2(n_342),
.B1(n_325),
.B2(n_92),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_352),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_352),
.C(n_357),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_355),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_361),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_4),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_347),
.B(n_363),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_353),
.A2(n_136),
.B1(n_106),
.B2(n_109),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_109),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_386),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_380),
.B(n_385),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_390),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_368),
.A2(n_358),
.B(n_360),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_4),
.B(n_5),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_364),
.Y(n_385)
);

AOI321xp33_ASAP7_75t_L g388 ( 
.A1(n_372),
.A2(n_364),
.A3(n_357),
.B1(n_122),
.B2(n_134),
.C(n_120),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_388),
.B(n_389),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_371),
.B(n_120),
.CI(n_97),
.CON(n_389),
.SN(n_389)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_387),
.A2(n_370),
.B(n_366),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_400),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_377),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_395),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_384),
.B(n_369),
.Y(n_395)
);

FAx1_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_371),
.CI(n_378),
.CON(n_397),
.SN(n_397)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_398),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_97),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_389),
.A2(n_122),
.B(n_127),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_401),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_106),
.C(n_17),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_407),
.Y(n_412)
);

OAI21x1_ASAP7_75t_SL g406 ( 
.A1(n_393),
.A2(n_4),
.B(n_6),
.Y(n_406)
);

AOI322xp5_ASAP7_75t_L g411 ( 
.A1(n_406),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_6),
.C(n_7),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_397),
.C(n_17),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_9),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_404),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_411),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_403),
.A2(n_6),
.B(n_9),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_414),
.C(n_9),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_412),
.A2(n_408),
.B(n_10),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_11),
.C(n_12),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_419),
.B(n_415),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_418),
.C(n_13),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_13),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_422),
.A2(n_13),
.B(n_17),
.Y(n_423)
);


endmodule