module fake_jpeg_25148_n_251 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_27),
.B1(n_42),
.B2(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_23),
.B1(n_24),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_52),
.B1(n_39),
.B2(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_55),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_26),
.B2(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_14),
.B1(n_31),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_58),
.B1(n_26),
.B2(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_28),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_35),
.C(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_37),
.B1(n_34),
.B2(n_43),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_26),
.B1(n_42),
.B2(n_14),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_43),
.B1(n_40),
.B2(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_43),
.B1(n_30),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_32),
.B1(n_30),
.B2(n_40),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_77),
.B1(n_44),
.B2(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_44),
.B1(n_65),
.B2(n_51),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_88),
.B(n_93),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_16),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_69),
.B1(n_66),
.B2(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_101),
.B1(n_81),
.B2(n_86),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_74),
.C(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_102),
.C(n_97),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_74),
.B1(n_62),
.B2(n_46),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_72),
.C(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_72),
.B1(n_56),
.B2(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_106),
.B1(n_80),
.B2(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_68),
.B1(n_65),
.B2(n_53),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_109),
.B(n_96),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_89),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_124),
.C(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_79),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_94),
.B1(n_78),
.B2(n_81),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_127),
.B1(n_110),
.B2(n_17),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_112),
.B1(n_107),
.B2(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_32),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_16),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_87),
.B1(n_17),
.B2(n_21),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_21),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_11),
.B(n_21),
.Y(n_134)
);

NOR4xp25_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_111),
.C(n_11),
.D(n_104),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_117),
.B1(n_120),
.B2(n_124),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_144),
.C(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_110),
.B1(n_18),
.B2(n_17),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_18),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_18),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_45),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_149),
.B(n_114),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_33),
.C(n_28),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_131),
.C(n_119),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_20),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_153),
.B(n_121),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_15),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_129),
.C(n_125),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_165),
.C(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_147),
.C(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_137),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_20),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_127),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_151),
.B1(n_138),
.B2(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_33),
.C(n_28),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_141),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_149),
.B1(n_140),
.B2(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_33),
.C(n_28),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_45),
.C(n_35),
.Y(n_189)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_164),
.B1(n_176),
.B2(n_175),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_140),
.C(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_193),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_160),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_45),
.C(n_28),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.C(n_173),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_20),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_45),
.C(n_28),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_162),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_206),
.B1(n_181),
.B2(n_191),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_179),
.A2(n_161),
.B(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_200),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_15),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_0),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_168),
.B1(n_167),
.B2(n_159),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_189),
.B1(n_182),
.B2(n_15),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_192),
.C(n_194),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_13),
.C(n_29),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_211),
.B(n_215),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_0),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_15),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_214),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_207),
.B1(n_197),
.B2(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_201),
.C(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_224),
.C(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_202),
.C(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_225),
.B(n_2),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_2),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_29),
.B(n_3),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_2),
.B(n_3),
.Y(n_230)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_216),
.B(n_3),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_2),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_29),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_29),
.C(n_6),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_5),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_237),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_244),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_5),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_247),
.B(n_244),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_7),
.B(n_9),
.Y(n_249)
);

AOI31xp33_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_7),
.A3(n_9),
.B(n_10),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_7),
.C(n_10),
.Y(n_251)
);


endmodule