module fake_jpeg_9299_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_23),
.Y(n_42)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_13),
.B1(n_16),
.B2(n_19),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_36),
.B(n_28),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_35),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_13),
.B1(n_23),
.B2(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_46),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_51),
.B(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_26),
.C(n_33),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_65),
.B(n_51),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_28),
.C(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_74),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_50),
.B1(n_40),
.B2(n_41),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_41),
.B1(n_64),
.B2(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_49),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_40),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_64),
.B1(n_53),
.B2(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_66),
.C(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_57),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_73),
.B(n_71),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_70),
.B(n_75),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_81),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_82),
.A3(n_91),
.B1(n_93),
.B2(n_95),
.C1(n_56),
.C2(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_9),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_21),
.C(n_2),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_106),
.A3(n_105),
.B1(n_29),
.B2(n_6),
.C1(n_3),
.C2(n_5),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_12),
.A3(n_24),
.B1(n_6),
.B2(n_3),
.C1(n_19),
.C2(n_1),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_24),
.Y(n_114)
);


endmodule