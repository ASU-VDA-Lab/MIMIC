module fake_jpeg_2182_n_660 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_660);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_660;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_2),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_13),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_8),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_60),
.B(n_61),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_64),
.Y(n_182)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_65),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_71),
.Y(n_147)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_70),
.B(n_75),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_8),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_72),
.B(n_73),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_74),
.B(n_80),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_26),
.B(n_7),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_26),
.B(n_10),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_87),
.B(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_89),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_90),
.Y(n_217)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_10),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_97),
.B(n_99),
.Y(n_169)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_6),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_100),
.Y(n_164)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_32),
.B(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_104),
.Y(n_173)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_32),
.B(n_5),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_30),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_119),
.Y(n_172)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_48),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_124),
.B(n_127),
.Y(n_192)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_29),
.Y(n_126)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_30),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_27),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_39),
.B1(n_20),
.B2(n_46),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_130),
.A2(n_35),
.B1(n_82),
.B2(n_81),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_60),
.B(n_59),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_137),
.B(n_155),
.Y(n_242)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_67),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_159),
.B(n_160),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_83),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_92),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_170),
.B(n_184),
.Y(n_243)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_64),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_171),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_68),
.B(n_59),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_178),
.B(n_186),
.Y(n_259)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_115),
.B(n_47),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_95),
.B(n_47),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_190),
.B(n_198),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_114),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_193),
.B(n_195),
.Y(n_267)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_65),
.B(n_57),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_129),
.B(n_57),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_199),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_98),
.B(n_48),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_86),
.B(n_51),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_125),
.B(n_49),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_205),
.B(n_206),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_113),
.B(n_51),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_49),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_209),
.A2(n_1),
.B(n_3),
.Y(n_278)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_78),
.B(n_46),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_212),
.B(n_16),
.Y(n_286)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_103),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_12),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_154),
.A2(n_89),
.B1(n_112),
.B2(n_109),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_221),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_332)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_164),
.A2(n_39),
.B1(n_56),
.B2(n_44),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_41),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_224),
.B(n_228),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_225),
.Y(n_344)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_132),
.Y(n_226)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_226),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_227),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_169),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_229),
.B(n_246),
.Y(n_326)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

INVx11_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_164),
.A2(n_44),
.B1(n_27),
.B2(n_85),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_231),
.A2(n_234),
.B1(n_282),
.B2(n_284),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_233),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_27),
.B1(n_44),
.B2(n_107),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_156),
.B(n_34),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_235),
.B(n_240),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_123),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_239),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_145),
.B(n_41),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_152),
.B(n_41),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_244),
.B(n_279),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_245),
.B(n_272),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_187),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_147),
.A2(n_94),
.B1(n_90),
.B2(n_77),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_173),
.A2(n_76),
.B1(n_35),
.B2(n_107),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_158),
.B(n_121),
.C(n_69),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_149),
.C(n_135),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_130),
.A2(n_41),
.B1(n_85),
.B2(n_128),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_146),
.Y(n_251)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_163),
.Y(n_252)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_189),
.B(n_41),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_254),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_168),
.A2(n_128),
.B1(n_54),
.B2(n_29),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_255),
.A2(n_138),
.B1(n_167),
.B2(n_201),
.Y(n_336)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_153),
.A2(n_54),
.B1(n_12),
.B2(n_15),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_187),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_261),
.B(n_149),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_263),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_140),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_148),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_144),
.Y(n_266)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_270),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_177),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_271),
.A2(n_161),
.B1(n_162),
.B2(n_202),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_139),
.Y(n_273)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_131),
.A2(n_15),
.B1(n_17),
.B2(n_4),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_277),
.A2(n_294),
.B1(n_217),
.B2(n_202),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_278),
.A2(n_289),
.B(n_293),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_134),
.B(n_5),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_214),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_188),
.A2(n_16),
.B1(n_18),
.B2(n_143),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_216),
.Y(n_318)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_141),
.A2(n_16),
.B(n_182),
.C(n_208),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_208),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_166),
.B(n_182),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_201),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_174),
.A2(n_166),
.B(n_175),
.C(n_135),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_218),
.A2(n_185),
.B1(n_148),
.B2(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_185),
.B(n_218),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_295),
.B(n_176),
.Y(n_352)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_175),
.Y(n_296)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_342),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_303),
.B(n_307),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_224),
.B(n_217),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_306),
.B(n_313),
.C(n_343),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_257),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_243),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_327),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_310),
.A2(n_315),
.B1(n_328),
.B2(n_276),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_235),
.B(n_138),
.C(n_216),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_318),
.B(n_227),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_142),
.B(n_179),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_233),
.A2(n_177),
.B1(n_200),
.B2(n_180),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_229),
.B(n_167),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_356),
.Y(n_359)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_355),
.B(n_292),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_279),
.A2(n_252),
.B1(n_280),
.B2(n_295),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_337),
.A2(n_265),
.B1(n_264),
.B2(n_246),
.Y(n_369)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_240),
.B(n_142),
.C(n_161),
.Y(n_343)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_293),
.A2(n_200),
.B1(n_176),
.B2(n_162),
.Y(n_345)
);

O2A1O1Ixp33_ASAP7_75t_SL g358 ( 
.A1(n_345),
.A2(n_221),
.B(n_271),
.C(n_294),
.Y(n_358)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_346),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_236),
.Y(n_350)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_352),
.B(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_237),
.Y(n_353)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_237),
.Y(n_354)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_245),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_183),
.Y(n_356)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_SL g430 ( 
.A1(n_358),
.A2(n_367),
.B(n_368),
.C(n_400),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_348),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_364),
.Y(n_405)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_244),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_259),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_383),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_332),
.A2(n_291),
.B1(n_286),
.B2(n_277),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_332),
.A2(n_228),
.B1(n_196),
.B2(n_254),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_369),
.A2(n_370),
.B1(n_397),
.B2(n_298),
.Y(n_435)
);

CKINVDCx12_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_324),
.B(n_242),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_331),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_307),
.B(n_238),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_381),
.Y(n_404)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_342),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_385),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_326),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_382),
.Y(n_426)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_386),
.A2(n_402),
.B1(n_232),
.B2(n_316),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_309),
.B(n_222),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_391),
.Y(n_428)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_297),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_249),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_390),
.Y(n_431)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_305),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_327),
.B(n_292),
.Y(n_391)
);

BUFx24_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_392),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_393),
.B(n_398),
.Y(n_438)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_396),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_283),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_304),
.A2(n_310),
.B1(n_328),
.B2(n_321),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_308),
.B(n_288),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_399),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_351),
.A2(n_196),
.B1(n_254),
.B2(n_183),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_287),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_401),
.Y(n_425)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_313),
.B(n_239),
.C(n_269),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_354),
.C(n_353),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_373),
.A2(n_322),
.B(n_349),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_406),
.A2(n_419),
.B(n_427),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_360),
.B(n_302),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_408),
.B(n_409),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_343),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g411 ( 
.A(n_379),
.B(n_384),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_L g459 ( 
.A1(n_411),
.A2(n_407),
.B(n_428),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_400),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_352),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_416),
.C(n_418),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_350),
.C(n_346),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_373),
.A2(n_322),
.B(n_311),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_364),
.B(n_375),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_424),
.C(n_432),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_397),
.A2(n_345),
.B1(n_329),
.B2(n_253),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_440),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_325),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_325),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_375),
.B(n_317),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_436),
.C(n_437),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_435),
.A2(n_398),
.B1(n_362),
.B2(n_366),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_317),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_239),
.C(n_312),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_384),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_385),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_383),
.A2(n_226),
.B1(n_334),
.B2(n_225),
.Y(n_440)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_379),
.A2(n_320),
.B(n_300),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_442),
.A2(n_392),
.B(n_371),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_404),
.B(n_365),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_444),
.B(n_446),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_414),
.B(n_367),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_414),
.B(n_359),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_447),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_449),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_429),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_454),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_431),
.B(n_396),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_457),
.Y(n_495)
);

OAI21xp33_ASAP7_75t_SL g506 ( 
.A1(n_452),
.A2(n_335),
.B(n_301),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_442),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_368),
.Y(n_457)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_458),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_459),
.B(n_460),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_410),
.B(n_393),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_431),
.A2(n_377),
.B1(n_370),
.B2(n_358),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_467),
.B1(n_422),
.B2(n_440),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_405),
.B(n_363),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_463),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_423),
.A2(n_377),
.B1(n_358),
.B2(n_378),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_464),
.A2(n_476),
.B1(n_478),
.B2(n_407),
.Y(n_487)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_471),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_466),
.B(n_436),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_430),
.A2(n_388),
.B1(n_382),
.B2(n_394),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_438),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_402),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_469),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_361),
.C(n_390),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_473),
.C(n_477),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_361),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_426),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_472),
.B(n_474),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_408),
.B(n_392),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_412),
.B(n_392),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_380),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_475),
.B(n_433),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_430),
.A2(n_357),
.B1(n_380),
.B2(n_376),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_409),
.B(n_376),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_483),
.A2(n_450),
.B1(n_472),
.B2(n_448),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_487),
.A2(n_457),
.B1(n_474),
.B2(n_449),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_488),
.B(n_494),
.Y(n_536)
);

NOR4xp25_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_420),
.C(n_424),
.D(n_419),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_489),
.B(n_497),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_445),
.A2(n_430),
.B(n_415),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_490),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_445),
.A2(n_406),
.B(n_430),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g541 ( 
.A(n_492),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_446),
.A2(n_415),
.B1(n_413),
.B2(n_437),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_493),
.A2(n_508),
.B1(n_512),
.B2(n_448),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_460),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_476),
.A2(n_415),
.B(n_426),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_496),
.B(n_498),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_467),
.A2(n_434),
.B(n_432),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_453),
.B(n_416),
.C(n_362),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_503),
.C(n_513),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_417),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_501),
.B(n_506),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_366),
.C(n_421),
.Y(n_503)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_507),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_447),
.A2(n_433),
.B1(n_344),
.B2(n_339),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_471),
.A2(n_475),
.B1(n_462),
.B2(n_463),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_509),
.A2(n_511),
.B1(n_316),
.B2(n_314),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_461),
.A2(n_232),
.B1(n_320),
.B2(n_300),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_454),
.A2(n_344),
.B1(n_298),
.B2(n_340),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_443),
.B(n_477),
.C(n_456),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_513),
.B(n_443),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_515),
.B(n_521),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_480),
.A2(n_444),
.B1(n_468),
.B2(n_462),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_517),
.A2(n_524),
.B1(n_532),
.B2(n_545),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_470),
.C(n_456),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_522),
.C(n_528),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_502),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_526),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_520),
.A2(n_538),
.B1(n_506),
.B2(n_512),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_482),
.B(n_455),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_455),
.C(n_473),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_466),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_543),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_525),
.A2(n_524),
.B1(n_490),
.B2(n_501),
.Y(n_557)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_500),
.B(n_451),
.C(n_458),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_529),
.Y(n_546)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_504),
.Y(n_531)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_531),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_480),
.A2(n_457),
.B1(n_465),
.B2(n_340),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_499),
.Y(n_533)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_335),
.C(n_323),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_539),
.C(n_503),
.Y(n_556)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_499),
.Y(n_535)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_535),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_484),
.B(n_312),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_537),
.B(n_510),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_501),
.A2(n_334),
.B1(n_251),
.B2(n_262),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_497),
.B(n_323),
.C(n_296),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_486),
.Y(n_540)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_540),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_314),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_542),
.A2(n_487),
.B1(n_479),
.B2(n_495),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_554),
.A2(n_560),
.B1(n_527),
.B2(n_530),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_536),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_555),
.B(n_566),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_556),
.B(n_563),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_557),
.A2(n_559),
.B1(n_274),
.B2(n_266),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_516),
.C(n_534),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_558),
.B(n_564),
.C(n_566),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_525),
.A2(n_483),
.B1(n_495),
.B2(n_510),
.Y(n_559)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_561),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_516),
.B(n_493),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_498),
.C(n_505),
.Y(n_564)
);

INVx6_ASAP7_75t_L g565 ( 
.A(n_526),
.Y(n_565)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_565),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_505),
.C(n_485),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_523),
.B(n_486),
.C(n_496),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_570),
.C(n_301),
.Y(n_588)
);

AOI21x1_ASAP7_75t_SL g569 ( 
.A1(n_527),
.A2(n_479),
.B(n_492),
.Y(n_569)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_569),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_522),
.B(n_507),
.C(n_481),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_514),
.A2(n_484),
.B1(n_509),
.B2(n_511),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_571),
.A2(n_230),
.B1(n_263),
.B2(n_241),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_559),
.A2(n_530),
.B(n_541),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_572),
.A2(n_563),
.B(n_548),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_550),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_573),
.B(n_577),
.Y(n_595)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_574),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_585),
.Y(n_597)
);

AOI322xp5_ASAP7_75t_SL g577 ( 
.A1(n_552),
.A2(n_489),
.A3(n_544),
.B1(n_491),
.B2(n_528),
.C1(n_508),
.C2(n_543),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_554),
.A2(n_491),
.B1(n_520),
.B2(n_544),
.Y(n_579)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_579),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_570),
.B(n_539),
.Y(n_582)
);

CKINVDCx14_ASAP7_75t_R g601 ( 
.A(n_582),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_565),
.B(n_538),
.Y(n_583)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_583),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_586),
.B(n_588),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_553),
.B(n_347),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_589),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_547),
.B(n_283),
.Y(n_589)
);

BUFx24_ASAP7_75t_SL g590 ( 
.A(n_547),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_590),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_546),
.B(n_275),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_592),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_567),
.A2(n_211),
.B1(n_347),
.B2(n_275),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_549),
.B(n_281),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_593),
.B(n_562),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_558),
.C(n_551),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_598),
.B(n_605),
.Y(n_625)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_602),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_572),
.A2(n_569),
.B(n_557),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_603),
.B(n_607),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_584),
.B(n_551),
.C(n_564),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_568),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_556),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_609),
.A2(n_610),
.B1(n_611),
.B2(n_330),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_560),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_576),
.B(n_548),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_612),
.A2(n_585),
.B(n_583),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_598),
.B(n_576),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_616),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_594),
.A2(n_581),
.B1(n_575),
.B2(n_579),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_615),
.A2(n_606),
.B1(n_610),
.B2(n_597),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_596),
.B(n_578),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_578),
.C(n_588),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_617),
.B(n_618),
.C(n_619),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_601),
.B(n_589),
.C(n_581),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_609),
.B(n_612),
.C(n_611),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_595),
.A2(n_607),
.B(n_608),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_620),
.A2(n_599),
.B1(n_606),
.B2(n_604),
.Y(n_633)
);

XOR2x2_ASAP7_75t_L g631 ( 
.A(n_621),
.B(n_597),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_594),
.B(n_281),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_623),
.B(n_602),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_603),
.B(n_290),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_627),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_269),
.Y(n_626)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_626),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_618),
.B(n_604),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_629),
.B(n_636),
.Y(n_640)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_631),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_632),
.A2(n_633),
.B1(n_256),
.B2(n_211),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_600),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_634),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_SL g636 ( 
.A1(n_613),
.A2(n_622),
.B1(n_619),
.B2(n_621),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_617),
.Y(n_639)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_639),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_636),
.A2(n_630),
.B(n_622),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_641),
.A2(n_642),
.B(n_643),
.Y(n_647)
);

NOR2x1_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_624),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_628),
.A2(n_615),
.B(n_600),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_646),
.B(n_635),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_645),
.B(n_628),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_648),
.A2(n_649),
.B(n_644),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_640),
.A2(n_629),
.B(n_637),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_650),
.B(n_640),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_652),
.A2(n_653),
.B(n_272),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_651),
.B(n_646),
.C(n_642),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_647),
.B(n_637),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_655),
.B(n_656),
.C(n_273),
.Y(n_657)
);

AO21x1_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_220),
.B(n_258),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_220),
.C(n_258),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_220),
.C(n_238),
.Y(n_660)
);


endmodule