module fake_jpeg_13891_n_604 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_604);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_604;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_17),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_62),
.Y(n_161)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_63),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_74),
.Y(n_130)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_68),
.Y(n_162)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_76),
.B(n_78),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_79),
.B(n_89),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_21),
.B(n_9),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_87),
.Y(n_136)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_23),
.B(n_7),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_24),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_20),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_90),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_43),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_106),
.Y(n_142)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_57),
.B(n_7),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_10),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_119),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_16),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_32),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_118),
.Y(n_199)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_122),
.Y(n_197)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_121),
.A2(n_34),
.B1(n_71),
.B2(n_93),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_89),
.B1(n_79),
.B2(n_90),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_124),
.A2(n_165),
.B1(n_191),
.B2(n_45),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_69),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_127),
.B(n_137),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_131),
.B(n_154),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_101),
.B1(n_105),
.B2(n_103),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_54),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_51),
.B1(n_53),
.B2(n_20),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_156),
.A2(n_176),
.B1(n_80),
.B2(n_73),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_170),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_54),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_159),
.B(n_167),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_51),
.B1(n_44),
.B2(n_42),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_44),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_42),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_169),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_25),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_111),
.B(n_25),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_182),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_61),
.A2(n_27),
.B1(n_41),
.B2(n_33),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_38),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_121),
.A2(n_45),
.B(n_15),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_52),
.B1(n_41),
.B2(n_33),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_188),
.A2(n_190),
.B1(n_0),
.B2(n_1),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_117),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_70),
.A2(n_38),
.B1(n_35),
.B2(n_30),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_130),
.Y(n_225)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_201),
.A2(n_202),
.B1(n_229),
.B2(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_131),
.A2(n_102),
.B1(n_92),
.B2(n_83),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g284 ( 
.A(n_204),
.Y(n_284)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_205),
.Y(n_317)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_208),
.Y(n_303)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_209),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g279 ( 
.A1(n_210),
.A2(n_239),
.B1(n_262),
.B2(n_128),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_156),
.A2(n_122),
.B1(n_45),
.B2(n_11),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_211),
.A2(n_215),
.B1(n_269),
.B2(n_186),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_216),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_219),
.B(n_242),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_220),
.B(n_227),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_225),
.A2(n_228),
.B(n_246),
.Y(n_305)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_226),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_138),
.B(n_5),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_4),
.B1(n_13),
.B2(n_12),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_232),
.Y(n_301)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_235),
.Y(n_310)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_236),
.Y(n_311)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_237),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_238),
.Y(n_320)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_3),
.B1(n_11),
.B2(n_12),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_241),
.Y(n_298)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_136),
.B(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_244),
.Y(n_304)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_153),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_197),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_245),
.B(n_249),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_142),
.B(n_15),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_259),
.B1(n_195),
.B2(n_149),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_185),
.Y(n_289)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_125),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_190),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_254),
.B(n_255),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_132),
.B(n_1),
.Y(n_255)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_258),
.B1(n_261),
.B2(n_266),
.Y(n_275)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_125),
.Y(n_257)
);

INVx8_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_161),
.A2(n_2),
.B1(n_193),
.B2(n_157),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_145),
.A2(n_181),
.B1(n_188),
.B2(n_129),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_123),
.Y(n_260)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_128),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_142),
.A2(n_176),
.B(n_175),
.C(n_173),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_133),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_263),
.Y(n_272)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_147),
.Y(n_266)
);

BUFx4f_ASAP7_75t_L g267 ( 
.A(n_139),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_267),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_268),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_129),
.A2(n_140),
.B1(n_186),
.B2(n_155),
.Y(n_269)
);

AO22x2_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_123),
.B1(n_126),
.B2(n_179),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_270),
.A2(n_211),
.B(n_268),
.C(n_269),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_126),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_271),
.B(n_296),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_195),
.C(n_185),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_274),
.B(n_293),
.C(n_294),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_276),
.A2(n_283),
.B1(n_222),
.B2(n_266),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_214),
.A2(n_161),
.B1(n_157),
.B2(n_174),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_278),
.A2(n_290),
.B1(n_299),
.B2(n_285),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_279),
.A2(n_208),
.B1(n_236),
.B2(n_234),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_210),
.A2(n_139),
.B1(n_155),
.B2(n_149),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_289),
.B(n_231),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_221),
.B(n_218),
.C(n_224),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_239),
.C(n_214),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_295),
.A2(n_256),
.B1(n_216),
.B2(n_230),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_179),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_151),
.C(n_192),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_323),
.C(n_227),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_262),
.A2(n_228),
.B1(n_235),
.B2(n_257),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_258),
.B(n_253),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_151),
.C(n_252),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_268),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_177),
.Y(n_360)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_271),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_332),
.Y(n_376)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

AO21x1_ASAP7_75t_L g386 ( 
.A1(n_331),
.A2(n_366),
.B(n_273),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_304),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_287),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_339),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_335),
.A2(n_320),
.B1(n_303),
.B2(n_309),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_237),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_351),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_298),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g395 ( 
.A1(n_340),
.A2(n_322),
.B(n_288),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_274),
.B(n_238),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_206),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_343),
.B(n_352),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_358),
.B1(n_359),
.B2(n_368),
.Y(n_373)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_346),
.Y(n_385)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_310),
.A2(n_209),
.B(n_192),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_347),
.A2(n_340),
.B(n_369),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_284),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_349),
.Y(n_396)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_350),
.A2(n_359),
.B1(n_328),
.B2(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_286),
.B(n_233),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_294),
.B(n_296),
.CI(n_289),
.CON(n_352),
.SN(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_284),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_354),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_272),
.B(n_170),
.Y(n_354)
);

INVx13_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_315),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_212),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_295),
.A2(n_310),
.B1(n_291),
.B2(n_270),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_291),
.A2(n_147),
.B1(n_177),
.B2(n_248),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_361),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_326),
.B(n_297),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_270),
.A2(n_204),
.B(n_267),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_309),
.B(n_303),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_292),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_363),
.Y(n_389)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_364),
.A2(n_369),
.B1(n_370),
.B2(n_285),
.Y(n_384)
);

AOI32xp33_ASAP7_75t_L g365 ( 
.A1(n_279),
.A2(n_204),
.A3(n_267),
.B1(n_270),
.B2(n_300),
.Y(n_365)
);

AOI32xp33_ASAP7_75t_L g379 ( 
.A1(n_365),
.A2(n_311),
.A3(n_319),
.B1(n_320),
.B2(n_277),
.Y(n_379)
);

XNOR2x1_ASAP7_75t_SL g366 ( 
.A(n_279),
.B(n_323),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_279),
.B(n_282),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_367),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_275),
.A2(n_313),
.B1(n_302),
.B2(n_318),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_290),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_387),
.B1(n_390),
.B2(n_406),
.Y(n_427)
);

OAI22x1_ASAP7_75t_SL g375 ( 
.A1(n_365),
.A2(n_299),
.B1(n_273),
.B2(n_318),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_375),
.A2(n_342),
.B1(n_329),
.B2(n_330),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_300),
.B(n_311),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_377),
.A2(n_393),
.B(n_398),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_379),
.A2(n_381),
.B(n_386),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_358),
.A2(n_324),
.B1(n_314),
.B2(n_306),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_324),
.B1(n_314),
.B2(n_306),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_391),
.A2(n_395),
.B(n_397),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_331),
.A2(n_307),
.B(n_288),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_307),
.B(n_316),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_356),
.A2(n_317),
.B(n_322),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_347),
.A2(n_316),
.B(n_317),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_401),
.A2(n_402),
.B(n_407),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_366),
.A2(n_281),
.B(n_312),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_312),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_404),
.B(n_357),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_338),
.A2(n_368),
.B1(n_341),
.B2(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_400),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_428),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_406),
.A2(n_350),
.B1(n_335),
.B2(n_333),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_413),
.A2(n_414),
.B1(n_420),
.B2(n_421),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_406),
.A2(n_335),
.B1(n_333),
.B2(n_352),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_332),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_415),
.B(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_339),
.Y(n_416)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_334),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_419),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_373),
.A2(n_352),
.B1(n_337),
.B2(n_351),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_373),
.A2(n_354),
.B1(n_361),
.B2(n_341),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_400),
.Y(n_422)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_422),
.Y(n_472)
);

INVx13_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_425),
.A2(n_438),
.B1(n_386),
.B2(n_381),
.Y(n_455)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_403),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_426),
.Y(n_475)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_431),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_382),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_336),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_394),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_377),
.A2(n_345),
.B(n_349),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_433),
.Y(n_470)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_434),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_377),
.A2(n_364),
.B(n_346),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_398),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_376),
.B(n_327),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_437),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_382),
.B(n_355),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_392),
.A2(n_405),
.B1(n_378),
.B2(n_379),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_404),
.B(n_380),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_439),
.B(n_441),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_389),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_440),
.B(n_380),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_372),
.B(n_392),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_396),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_443),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_409),
.A2(n_378),
.B1(n_375),
.B2(n_386),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_444),
.A2(n_438),
.B(n_401),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_445),
.B(n_453),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_443),
.A2(n_389),
.B1(n_371),
.B2(n_384),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

NOR3xp33_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_436),
.C(n_428),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_449),
.B(n_398),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_432),
.B(n_408),
.Y(n_453)
);

OAI21xp33_ASAP7_75t_SL g454 ( 
.A1(n_416),
.A2(n_407),
.B(n_401),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_R g493 ( 
.A(n_454),
.B(n_471),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_L g498 ( 
.A(n_455),
.B(n_456),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_375),
.B1(n_395),
.B2(n_393),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_456),
.A2(n_474),
.B1(n_423),
.B2(n_429),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_425),
.A2(n_386),
.B1(n_373),
.B2(n_374),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_461),
.A2(n_413),
.B1(n_421),
.B2(n_410),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_415),
.A2(n_388),
.B1(n_387),
.B2(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_437),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_431),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_396),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_440),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_402),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_469),
.B(n_471),
.C(n_441),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_402),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_427),
.A2(n_393),
.B1(n_407),
.B2(n_387),
.Y(n_474)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_477),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g520 ( 
.A(n_478),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_457),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_480),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_457),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_411),
.Y(n_481)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_481),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_498),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_419),
.Y(n_484)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_484),
.Y(n_516)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_487),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_444),
.A2(n_410),
.B(n_423),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_489),
.Y(n_507)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_490),
.A2(n_501),
.B1(n_467),
.B2(n_460),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_492),
.B1(n_458),
.B2(n_451),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_474),
.A2(n_429),
.B1(n_430),
.B2(n_433),
.Y(n_492)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_496),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_470),
.A2(n_391),
.B(n_442),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_494),
.B(n_499),
.Y(n_509)
);

AO21x1_ASAP7_75t_L g495 ( 
.A1(n_448),
.A2(n_435),
.B(n_442),
.Y(n_495)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_495),
.A2(n_461),
.B1(n_451),
.B2(n_458),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_417),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_502),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_459),
.B(n_439),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_500),
.B(n_462),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_460),
.B(n_422),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_412),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_503),
.B(n_450),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_445),
.C(n_448),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_511),
.C(n_512),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_469),
.C(n_453),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_450),
.C(n_467),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_514),
.A2(n_484),
.B(n_481),
.Y(n_532)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_523),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_521),
.Y(n_538)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_522),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_441),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_482),
.A2(n_462),
.B1(n_475),
.B2(n_473),
.Y(n_524)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_524),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_495),
.B(n_475),
.C(n_391),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_491),
.C(n_495),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_482),
.A2(n_472),
.B1(n_412),
.B2(n_452),
.Y(n_526)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_526),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_509),
.A2(n_494),
.B(n_476),
.Y(n_529)
);

OAI21x1_ASAP7_75t_SL g560 ( 
.A1(n_529),
.A2(n_496),
.B(n_501),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_507),
.A2(n_488),
.B(n_496),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_530),
.A2(n_532),
.B(n_483),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_521),
.Y(n_547)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_516),
.Y(n_533)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_533),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_508),
.B(n_492),
.C(n_498),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_541),
.Y(n_556)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_505),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_517),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_544),
.Y(n_551)
);

OAI21xp33_ASAP7_75t_L g543 ( 
.A1(n_520),
.A2(n_497),
.B(n_490),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_543),
.Y(n_549)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_527),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_506),
.A2(n_479),
.B1(n_480),
.B2(n_477),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_545),
.A2(n_513),
.B1(n_538),
.B2(n_539),
.Y(n_548)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_524),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_515),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_547),
.B(n_554),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_548),
.B(n_552),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_525),
.C(n_526),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_535),
.B(n_478),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_553),
.B(n_558),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_557),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_510),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_510),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_529),
.B(n_512),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_559),
.B(n_561),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_560),
.A2(n_536),
.B1(n_539),
.B2(n_540),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_SL g561 ( 
.A(n_537),
.B(n_511),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_538),
.A2(n_487),
.B1(n_485),
.B2(n_518),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_562),
.B(n_518),
.Y(n_574)
);

BUFx24_ASAP7_75t_SL g565 ( 
.A(n_556),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_565),
.B(n_573),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_549),
.B(n_499),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_566),
.B(n_569),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_547),
.B(n_540),
.C(n_528),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_570),
.A2(n_501),
.B(n_504),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_552),
.A2(n_528),
.B(n_536),
.Y(n_571)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_571),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_515),
.C(n_532),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_569),
.C(n_564),
.Y(n_577)
);

FAx1_ASAP7_75t_SL g573 ( 
.A(n_555),
.B(n_530),
.CI(n_545),
.CON(n_573),
.SN(n_573)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_523),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_550),
.B1(n_533),
.B2(n_502),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_576),
.A2(n_579),
.B1(n_581),
.B2(n_582),
.Y(n_590)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_577),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_572),
.A2(n_518),
.B1(n_559),
.B2(n_562),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_564),
.A2(n_489),
.B1(n_472),
.B2(n_412),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_584),
.B(n_426),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_561),
.C(n_558),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_568),
.C(n_563),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_586),
.B(n_587),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_577),
.B(n_573),
.C(n_519),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_580),
.B(n_504),
.C(n_551),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_588),
.B(n_585),
.Y(n_596)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_589),
.Y(n_594)
);

XNOR2x1_ASAP7_75t_L g591 ( 
.A(n_579),
.B(n_424),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_591),
.B(n_581),
.C(n_583),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_593),
.A2(n_596),
.B(n_586),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_597),
.B(n_598),
.C(n_594),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_595),
.A2(n_592),
.B(n_578),
.Y(n_598)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_599),
.Y(n_600)
);

AO21x1_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_590),
.B(n_591),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_601),
.A2(n_397),
.B(n_434),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_602),
.B(n_397),
.C(n_424),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_383),
.B1(n_390),
.B2(n_583),
.Y(n_604)
);


endmodule