module fake_jpeg_23262_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_49),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_56),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_37),
.B(n_17),
.C(n_19),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_75),
.B1(n_78),
.B2(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_37),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_45),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_20),
.B(n_23),
.C(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_0),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_64),
.B1(n_69),
.B2(n_71),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_19),
.B1(n_31),
.B2(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_23),
.B1(n_28),
.B2(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_25),
.B1(n_35),
.B2(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_73),
.Y(n_100)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_49),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_87),
.B1(n_108),
.B2(n_110),
.Y(n_139)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_95),
.Y(n_152)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_93),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_90),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_91),
.B(n_97),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_92),
.Y(n_148)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_39),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_39),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_49),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_48),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_61),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_115),
.B1(n_96),
.B2(n_84),
.Y(n_137)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_45),
.B1(n_43),
.B2(n_48),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_77),
.B1(n_73),
.B2(n_45),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_130),
.B1(n_104),
.B2(n_94),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_89),
.B1(n_116),
.B2(n_95),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_91),
.B1(n_93),
.B2(n_82),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_85),
.B(n_105),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_52),
.C(n_45),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_124),
.C(n_129),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_48),
.C(n_43),
.Y(n_124)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_43),
.C(n_42),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_55),
.B1(n_42),
.B2(n_26),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_143),
.Y(n_176)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_26),
.B(n_22),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_108),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_147),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_86),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_154),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_155),
.A2(n_179),
.B(n_184),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_111),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_180),
.B1(n_182),
.B2(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_130),
.B1(n_124),
.B2(n_139),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_109),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_162),
.B(n_167),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_144),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_36),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_118),
.B(n_0),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_170),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_55),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_3),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_42),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_4),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_181),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_21),
.B(n_18),
.C(n_6),
.D(n_7),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_76),
.B1(n_21),
.B2(n_18),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_4),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_121),
.A2(n_18),
.B1(n_6),
.B2(n_7),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_125),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_5),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_128),
.B(n_5),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_188),
.B(n_200),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_193),
.B1(n_196),
.B2(n_202),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_197),
.B(n_216),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_136),
.B1(n_143),
.B2(n_127),
.Y(n_192)
);

AOI22x1_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_179),
.B1(n_180),
.B2(n_184),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_160),
.B1(n_171),
.B2(n_169),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_125),
.B1(n_150),
.B2(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_120),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_182),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_176),
.A2(n_5),
.B(n_6),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_215),
.B(n_185),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_8),
.B(n_9),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_9),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_218),
.A2(n_233),
.B1(n_241),
.B2(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_226),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_228),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_162),
.B(n_177),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_165),
.C(n_167),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_232),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_184),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_175),
.B(n_170),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_193),
.B(n_10),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_212),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_186),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_209),
.Y(n_251)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_203),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_187),
.A2(n_10),
.B(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_11),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_254),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_197),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_211),
.B1(n_196),
.B2(n_189),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_255),
.A2(n_259),
.B1(n_260),
.B2(n_218),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_244),
.B1(n_252),
.B2(n_250),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_209),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_245),
.B(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_216),
.B1(n_204),
.B2(n_188),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_205),
.B1(n_208),
.B2(n_212),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_208),
.B1(n_198),
.B2(n_215),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_263),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_235),
.C(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_273),
.C(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_221),
.C(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_239),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_276),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_222),
.B1(n_224),
.B2(n_237),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_278),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_226),
.B1(n_227),
.B2(n_225),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_225),
.B(n_223),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_281),
.A2(n_255),
.B1(n_258),
.B2(n_215),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_279),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_291),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_279),
.B1(n_271),
.B2(n_267),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_258),
.B1(n_253),
.B2(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_199),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_264),
.C(n_265),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_214),
.C(n_14),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_214),
.C(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_299),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_283),
.B(n_288),
.C(n_284),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_269),
.C(n_280),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_280),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_293),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_286),
.Y(n_312)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_307),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_312),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_310),
.B(n_301),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_292),
.B(n_266),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_317),
.B1(n_299),
.B2(n_287),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_306),
.B(n_298),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_320),
.A2(n_321),
.B(n_318),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_288),
.B(n_307),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_270),
.B(n_296),
.Y(n_324)
);

AOI321xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_12),
.A3(n_15),
.B1(n_16),
.B2(n_323),
.C(n_319),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_12),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_15),
.Y(n_327)
);


endmodule