module real_jpeg_13658_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_244;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_68),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_70),
.Y(n_203)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_6),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_6),
.A2(n_59),
.B1(n_62),
.B2(n_149),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_149),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_149),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_59),
.B1(n_62),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_7),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_78),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_12),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_12),
.A2(n_59),
.B1(n_62),
.B2(n_101),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_101),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_101),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_13),
.A2(n_52),
.B1(n_59),
.B2(n_62),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_14),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_14),
.A2(n_64),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_14),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_14),
.B(n_62),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_141),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_14),
.A2(n_43),
.B(n_48),
.C(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_14),
.B(n_109),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_14),
.B(n_32),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_14),
.B(n_53),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_14),
.A2(n_62),
.B(n_200),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_16),
.A2(n_45),
.B1(n_59),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_45),
.Y(n_137)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_86),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_23),
.B(n_80),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_28),
.A2(n_32),
.B(n_37),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_28),
.A2(n_32),
.B1(n_92),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_28),
.A2(n_32),
.B1(n_137),
.B2(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_28),
.A2(n_32),
.B1(n_179),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_28),
.A2(n_32),
.B1(n_203),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_28),
.A2(n_32),
.B1(n_141),
.B2(n_236),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_28),
.A2(n_32),
.B1(n_229),
.B2(n_236),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_29),
.B(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_31),
.A2(n_34),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_31),
.A2(n_90),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_35),
.A2(n_49),
.B(n_141),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_50),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_44),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_43),
.B(n_74),
.Y(n_201)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_44),
.A2(n_62),
.A3(n_75),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_46),
.A2(n_53),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_46),
.A2(n_53),
.B1(n_95),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_46),
.A2(n_53),
.B1(n_167),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_46),
.A2(n_53),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_46),
.A2(n_53),
.B1(n_215),
.B2(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_50),
.A2(n_96),
.B1(n_194),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_57),
.A2(n_58),
.B1(n_148),
.B2(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_60),
.B(n_62),
.Y(n_139)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_65),
.B(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_72),
.A2(n_73),
.B1(n_144),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_72),
.A2(n_73),
.B1(n_175),
.B2(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_73),
.Y(n_109)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_82),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_88),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_89),
.B(n_93),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_99),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_123),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B(n_112),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_109),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_107),
.A2(n_109),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_155),
.B(n_270),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_153),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_127),
.B(n_153),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_133),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_132),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_133),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_142),
.C(n_146),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_146),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_186),
.B(n_264),
.C(n_269),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_180),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_157),
.B(n_180),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_170),
.C(n_172),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_159),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_164),
.C(n_169),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_170),
.B(n_172),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.C(n_178),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_183),
.C(n_184),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_263),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_207),
.B(n_262),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_204),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_189),
.B(n_204),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_195),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_190),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_192),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_256),
.B(n_261),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_245),
.B(n_255),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_225),
.B(n_244),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_221),
.C(n_223),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_233),
.B(n_243),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_242),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);


endmodule