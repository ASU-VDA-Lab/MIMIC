module fake_jpeg_9148_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_14),
.Y(n_15)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_16),
.A2(n_6),
.B1(n_9),
.B2(n_7),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_18),
.B1(n_9),
.B2(n_7),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_16),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_15),
.B(n_8),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_15),
.C(n_8),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.C(n_9),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_11),
.B1(n_10),
.B2(n_19),
.Y(n_29)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_16),
.B1(n_11),
.B2(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_29),
.B(n_30),
.C(n_2),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_5),
.A3(n_16),
.B1(n_12),
.B2(n_3),
.C1(n_0),
.C2(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_5),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_16),
.Y(n_39)
);


endmodule