module fake_jpeg_21321_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_31),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_13),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_15),
.B1(n_20),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_48),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_15),
.B1(n_20),
.B2(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_33),
.B1(n_36),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_49),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_36),
.B1(n_32),
.B2(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_60),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_28),
.B1(n_30),
.B2(n_26),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_26),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_24),
.B1(n_21),
.B2(n_14),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_21),
.B(n_24),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_63),
.B1(n_57),
.B2(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_49),
.B1(n_61),
.B2(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_62),
.C(n_63),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_72),
.C(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_92),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NOR4xp25_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_77),
.C(n_79),
.D(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_38),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_100),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_85),
.C(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_68),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_88),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_97),
.B(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_83),
.B1(n_80),
.B2(n_85),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_38),
.C(n_39),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_69),
.B1(n_12),
.B2(n_5),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_100),
.B1(n_95),
.B2(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_69),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_118),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_12),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_30),
.C(n_28),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_105),
.B(n_106),
.C(n_110),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_2),
.B(n_7),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_116),
.B1(n_39),
.B2(n_9),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_7),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_119),
.C(n_121),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B1(n_123),
.B2(n_9),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_2),
.B(n_7),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_130),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_28),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_129),
.B(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_132),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_28),
.Y(n_135)
);


endmodule