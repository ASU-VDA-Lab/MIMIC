module fake_jpeg_2363_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

INVx11_ASAP7_75t_SL g9 ( 
.A(n_4),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_5),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_15),
.B1(n_19),
.B2(n_16),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_19),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_20),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_23),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_19),
.B1(n_18),
.B2(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_19),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_23),
.C(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_12),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_31),
.C(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_30),
.B1(n_15),
.B2(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_38),
.B1(n_15),
.B2(n_2),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_38),
.C(n_39),
.Y(n_48)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_41),
.CI(n_43),
.CON(n_47),
.SN(n_47)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_48),
.B2(n_47),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_44),
.B(n_15),
.Y(n_50)
);

OAI31xp33_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_47),
.A3(n_48),
.B(n_6),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_7),
.C1(n_20),
.C2(n_17),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_3),
.Y(n_54)
);


endmodule