module fake_netlist_5_858_n_2086 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_2086);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2086;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_2001;
wire n_1494;
wire n_625;
wire n_1462;
wire n_854;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1243;
wire n_1016;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_1070;
wire n_777;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_464;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1538;
wire n_1162;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_1537;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_1989;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_512;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_1343;
wire n_1631;
wire n_1203;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_1937;
wire n_585;
wire n_1739;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_203),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_126),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_116),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_235),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_248),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_111),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_298),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

BUFx10_ASAP7_75t_L g405 ( 
.A(n_83),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_363),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_254),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_269),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_62),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_302),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_336),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_241),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_172),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_95),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_160),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_244),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_314),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_64),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_29),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_6),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_178),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_247),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_274),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_204),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_211),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_393),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_372),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_323),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_263),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_164),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_56),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_65),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_251),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_205),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_187),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_57),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_40),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_309),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_146),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_150),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_106),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_168),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_54),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_267),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_69),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_98),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_394),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_210),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_276),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_288),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_321),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_386),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_357),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_149),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_189),
.Y(n_461)
);

BUFx8_ASAP7_75t_SL g462 ( 
.A(n_43),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_137),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_342),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_318),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_378),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_125),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_358),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_306),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_325),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_31),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_310),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_91),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_14),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_39),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_215),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_220),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_207),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_34),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_285),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_315),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_395),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_190),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_332),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_30),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_43),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_152),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_166),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_209),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_49),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_221),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_287),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_183),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_346),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_50),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_67),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_359),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_322),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_252),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_112),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_200),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_326),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_292),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_256),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_345),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_148),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_223),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_195),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_319),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_29),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_79),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_333),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_17),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_15),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_381),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_3),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_119),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_268),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_127),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_213),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_206),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_331),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_36),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_356),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_7),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_158),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_197),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_253),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_352),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_388),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_182),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_330),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_142),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_245),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_387),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_141),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_85),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_81),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_301),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_360),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_120),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_143),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_316),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_351),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_277),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_129),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_123),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_340),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_305),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_59),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_163),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_341),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_238),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_36),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_246),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_344),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_218),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_58),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_364),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_37),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_133),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_374),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_40),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_117),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_202),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_173),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_355),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_156),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_233),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_121),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_328),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_165),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_384),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_3),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_61),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_232),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_97),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_1),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_258),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_70),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_28),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_377),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_100),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_339),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_317),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_21),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_243),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_266),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_131),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_82),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_334),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_313),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_144),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_8),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_212),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_389),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_124),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_47),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_10),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_371),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_385),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_396),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_280),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_350),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_383),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_201),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_132),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_278),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_257),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_327),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_118),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_373),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_264),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_18),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_349),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_90),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_300),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_31),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_8),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_49),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_369),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_41),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_180),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_74),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_225),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_236),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_32),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_9),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_271),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_4),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_228),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_175),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_161),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_299),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_297),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_139),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_234),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_311),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_335),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_19),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_101),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_329),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_159),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_21),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_250),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_96),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_136),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_11),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_6),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_366),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_35),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_38),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_240),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_5),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_255),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_50),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_237),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_354),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_260),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_63),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_368),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_105),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_337),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_68),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_9),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_99),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_296),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_135),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_103),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_320),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_227),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_138),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_275),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_379),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_42),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_194),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_42),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_343),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_7),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_87),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_22),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_279),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_370),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_361),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_108),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_226),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_231),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_171),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_188),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_308),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_46),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_11),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_273),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_282),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_128),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_80),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_47),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_107),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_35),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_113),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_283),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_94),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_185),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_353),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_153),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_174),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_193),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_365),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_324),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_147),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_392),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_230),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_92),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_41),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_169),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_362),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_45),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_347),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_491),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_398),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_645),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_462),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_405),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_645),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_645),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_397),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_645),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_692),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_645),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_400),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_491),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_491),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_645),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_491),
.Y(n_735)
);

CKINVDCx16_ASAP7_75t_R g736 ( 
.A(n_475),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_698),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_401),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_698),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_698),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_698),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_524),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_555),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_402),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_561),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_403),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_406),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_564),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_587),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_422),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_407),
.Y(n_751)
);

INVxp33_ASAP7_75t_SL g752 ( 
.A(n_423),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_620),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_621),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_629),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_452),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_641),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_693),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_700),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_455),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_408),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_628),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_461),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_399),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_409),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_666),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_404),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_411),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_413),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_415),
.Y(n_771)
);

INVxp33_ASAP7_75t_SL g772 ( 
.A(n_442),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_420),
.Y(n_773)
);

INVxp33_ASAP7_75t_SL g774 ( 
.A(n_471),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_579),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_425),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_490),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_492),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_432),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_427),
.Y(n_780)
);

INVxp67_ASAP7_75t_SL g781 ( 
.A(n_505),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_539),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_410),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_436),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_541),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_676),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_433),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_439),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_458),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_441),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_663),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_507),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_412),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_516),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_414),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_416),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_444),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_556),
.Y(n_798)
);

INVxp33_ASAP7_75t_SL g799 ( 
.A(n_476),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_676),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_446),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_454),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_417),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_456),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_537),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_576),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_418),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_405),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_428),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_469),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_463),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_585),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_473),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_419),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_474),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_479),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_484),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_480),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_488),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_591),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_421),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_608),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_500),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_510),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_637),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_486),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_518),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_428),
.Y(n_828)
);

INVxp33_ASAP7_75t_SL g829 ( 
.A(n_496),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_511),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_424),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_527),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_530),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_536),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_640),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_459),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_428),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_538),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_514),
.Y(n_839)
);

INVxp33_ASAP7_75t_L g840 ( 
.A(n_547),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_426),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_553),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_554),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_559),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_467),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_642),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_648),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_566),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_571),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_515),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_706),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_580),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_501),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_583),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_517),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_590),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_592),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_526),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_428),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_594),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_598),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_602),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_603),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_694),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_605),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_685),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_703),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_606),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_611),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_448),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_625),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_630),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_575),
.B(n_0),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_582),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_429),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_635),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_696),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_448),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_487),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_448),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_636),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_643),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_430),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_647),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_659),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_448),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_549),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_664),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_667),
.Y(n_889)
);

CKINVDCx16_ASAP7_75t_R g890 ( 
.A(n_459),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_671),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_673),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_683),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_691),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_595),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_701),
.Y(n_896)
);

INVxp33_ASAP7_75t_SL g897 ( 
.A(n_599),
.Y(n_897)
);

CKINVDCx14_ASAP7_75t_R g898 ( 
.A(n_481),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_431),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_468),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_434),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_708),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_713),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_435),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_600),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_437),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_714),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_468),
.Y(n_908)
);

CKINVDCx16_ASAP7_75t_R g909 ( 
.A(n_481),
.Y(n_909)
);

BUFx2_ASAP7_75t_SL g910 ( 
.A(n_568),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_615),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_438),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_717),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_443),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_440),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_445),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_498),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_519),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_447),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_449),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_523),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_619),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_568),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_468),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_525),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_658),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_468),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_503),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_450),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_503),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_503),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_451),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_453),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_503),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_631),
.Y(n_935)
);

INVxp33_ASAP7_75t_SL g936 ( 
.A(n_649),
.Y(n_936)
);

INVxp33_ASAP7_75t_SL g937 ( 
.A(n_650),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_567),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_652),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_567),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_567),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_567),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_457),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_464),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_618),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_618),
.Y(n_946)
);

INVxp33_ASAP7_75t_L g947 ( 
.A(n_618),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_618),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_653),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_465),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_596),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_699),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_466),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_655),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_470),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_657),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_472),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_678),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_680),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_682),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_718),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_460),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_482),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_662),
.Y(n_964)
);

INVx4_ASAP7_75t_R g965 ( 
.A(n_502),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_477),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_478),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_687),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_699),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_702),
.Y(n_970)
);

INVxp33_ASAP7_75t_L g971 ( 
.A(n_623),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_702),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_483),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_597),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_485),
.Y(n_975)
);

CKINVDCx16_ASAP7_75t_R g976 ( 
.A(n_508),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_489),
.Y(n_977)
);

CKINVDCx16_ASAP7_75t_R g978 ( 
.A(n_493),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_494),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_495),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_638),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_497),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_499),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_504),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_506),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_509),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_512),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_513),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_727),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_979),
.B(n_520),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_723),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_731),
.B(n_521),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_735),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_845),
.B(n_522),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_737),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_739),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_870),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_870),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_738),
.B(n_528),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_794),
.A2(n_531),
.B1(n_532),
.B2(n_529),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_740),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_741),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_870),
.Y(n_1003)
);

BUFx8_ASAP7_75t_L g1004 ( 
.A(n_786),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_878),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_780),
.Y(n_1006)
);

OA21x2_ASAP7_75t_L g1007 ( 
.A1(n_722),
.A2(n_534),
.B(n_533),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_880),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_720),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_784),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_886),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_900),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_744),
.B(n_535),
.Y(n_1013)
);

BUFx8_ASAP7_75t_L g1014 ( 
.A(n_969),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_811),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_720),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_924),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_949),
.B(n_540),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_753),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_732),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_732),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_746),
.B(n_542),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_910),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_733),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_729),
.A2(n_544),
.B1(n_545),
.B2(n_543),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_734),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_927),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_747),
.B(n_546),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_928),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_763),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_733),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_767),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_976),
.A2(n_550),
.B1(n_551),
.B2(n_548),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_930),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_749),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_853),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_724),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_L g1038 ( 
.A(n_791),
.B(n_552),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_800),
.A2(n_558),
.B1(n_560),
.B2(n_557),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_864),
.B(n_562),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_826),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_752),
.B(n_563),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_931),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_751),
.B(n_565),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_934),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_877),
.B(n_569),
.Y(n_1046)
);

INVx6_ASAP7_75t_L g1047 ( 
.A(n_808),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_762),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_938),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_836),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_766),
.B(n_570),
.Y(n_1051)
);

AND2x6_ASAP7_75t_L g1052 ( 
.A(n_725),
.B(n_52),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_800),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_940),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_742),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_941),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_942),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_946),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_948),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_858),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_743),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_726),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_745),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_809),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_SL g1065 ( 
.A(n_840),
.B(n_952),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_809),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_748),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_750),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_783),
.B(n_572),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_954),
.B(n_956),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_728),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_828),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_730),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_818),
.B(n_573),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_792),
.A2(n_577),
.B1(n_578),
.B2(n_574),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_772),
.B(n_581),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_754),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_755),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_757),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_828),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_758),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_759),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_874),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_760),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_793),
.B(n_584),
.Y(n_1085)
);

CKINVDCx14_ASAP7_75t_R g1086 ( 
.A(n_898),
.Y(n_1086)
);

OA21x2_ASAP7_75t_L g1087 ( 
.A1(n_837),
.A2(n_588),
.B(n_586),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_795),
.B(n_719),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_837),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_789),
.A2(n_593),
.B1(n_601),
.B2(n_589),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_774),
.B(n_604),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_796),
.B(n_607),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_915),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_765),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_859),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_818),
.B(n_609),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_958),
.B(n_610),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_768),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_859),
.A2(n_613),
.B(n_612),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_736),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_908),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_908),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_769),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_945),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_917),
.Y(n_1105)
);

INVx5_ASAP7_75t_L g1106 ( 
.A(n_890),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_918),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_945),
.A2(n_616),
.B(n_614),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_770),
.Y(n_1109)
);

AND2x2_ASAP7_75t_SL g1110 ( 
.A(n_909),
.B(n_0),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_921),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_895),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_771),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_773),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_863),
.A2(n_622),
.B1(n_624),
.B2(n_617),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_925),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_926),
.Y(n_1117)
);

AND2x2_ASAP7_75t_SL g1118 ( 
.A(n_923),
.B(n_1),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_776),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_779),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_803),
.B(n_626),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_807),
.B(n_716),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_978),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_959),
.B(n_627),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_830),
.B(n_632),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_960),
.B(n_633),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_799),
.B(n_634),
.Y(n_1127)
);

XOR2xp5_ASAP7_75t_L g1128 ( 
.A(n_971),
.B(n_2),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_787),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_866),
.Y(n_1130)
);

OAI22x1_ASAP7_75t_SL g1131 ( 
.A1(n_879),
.A2(n_712),
.B1(n_711),
.B2(n_710),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_961),
.B(n_639),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_788),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_867),
.A2(n_709),
.B1(n_707),
.B2(n_705),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_939),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_829),
.B(n_644),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_830),
.B(n_646),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_790),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_797),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_839),
.B(n_651),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_SL g1141 ( 
.A1(n_721),
.A2(n_704),
.B1(n_697),
.B2(n_695),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_814),
.B(n_690),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_801),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_973),
.B(n_654),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_805),
.A2(n_674),
.B1(n_688),
.B2(n_686),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_975),
.B(n_656),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_781),
.A2(n_672),
.B1(n_684),
.B2(n_681),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_802),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_L g1149 ( 
.A(n_980),
.B(n_660),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_821),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_883),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_831),
.B(n_689),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_804),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_906),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_810),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_813),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_897),
.B(n_935),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_982),
.B(n_661),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_841),
.B(n_679),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_983),
.B(n_665),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_815),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_816),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_817),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_819),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_823),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_839),
.B(n_850),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_824),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_875),
.B(n_677),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_970),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_850),
.B(n_668),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1100),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1062),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1071),
.Y(n_1173)
);

OAI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1033),
.A2(n_781),
.B1(n_951),
.B2(n_887),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1073),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1026),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1012),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1074),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1064),
.B(n_981),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1123),
.B(n_899),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1012),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1030),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1026),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_L g1184 ( 
.A(n_1166),
.B(n_905),
.C(n_855),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1072),
.B(n_936),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1123),
.B(n_990),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1053),
.B(n_855),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1030),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1007),
.A2(n_832),
.B(n_827),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1032),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1043),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1032),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1053),
.B(n_905),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1080),
.B(n_937),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1003),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_L g1196 ( 
.A(n_1052),
.B(n_984),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1049),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1089),
.B(n_901),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1047),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1037),
.B(n_911),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1049),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_922),
.C(n_911),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1054),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1054),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1056),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1056),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_997),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_992),
.B(n_904),
.Y(n_1208)
);

INVxp67_ASAP7_75t_R g1209 ( 
.A(n_1131),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1043),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_997),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1005),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1008),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1045),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1011),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_998),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1064),
.B(n_1066),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1045),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1066),
.B(n_988),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1057),
.Y(n_1220)
);

INVxp33_ASAP7_75t_L g1221 ( 
.A(n_1035),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_989),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1017),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1006),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_999),
.B(n_916),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1096),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_998),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1057),
.Y(n_1228)
);

AND3x2_ASAP7_75t_L g1229 ( 
.A(n_1023),
.B(n_775),
.C(n_951),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1027),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_1110),
.B(n_972),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1029),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1050),
.B(n_922),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1009),
.B(n_985),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1106),
.B(n_912),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1095),
.B(n_986),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1034),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1059),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1052),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_993),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1125),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1129),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1135),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_995),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_996),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1123),
.B(n_919),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1001),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1058),
.Y(n_1248)
);

AND2x6_ASAP7_75t_L g1249 ( 
.A(n_1149),
.B(n_987),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1095),
.B(n_920),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_1042),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1038),
.B(n_974),
.C(n_932),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1148),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1010),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_SL g1255 ( 
.A(n_1118),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1058),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_L g1257 ( 
.A(n_1052),
.B(n_929),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1106),
.B(n_933),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1002),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1013),
.B(n_944),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1120),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1019),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_994),
.B(n_950),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1019),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1153),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1155),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1165),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1047),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1101),
.B(n_957),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1101),
.B(n_967),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1015),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1102),
.B(n_977),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1167),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1141),
.A2(n_943),
.B1(n_953),
.B2(n_914),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1048),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1102),
.B(n_833),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1007),
.A2(n_1104),
.B(n_1009),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1104),
.B(n_775),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1036),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1137),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_SL g1281 ( 
.A(n_1151),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1093),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1105),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1120),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1161),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1107),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1161),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1116),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1077),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1098),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1163),
.Y(n_1291)
);

INVx8_ASAP7_75t_L g1292 ( 
.A(n_991),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1079),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1040),
.B(n_834),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1022),
.A2(n_842),
.B(n_838),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1081),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1163),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1113),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1082),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1098),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1103),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1143),
.Y(n_1302)
);

BUFx16f_ASAP7_75t_R g1303 ( 
.A(n_1014),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1130),
.B(n_1154),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1103),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1046),
.B(n_843),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1109),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1111),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1109),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_1041),
.B(n_963),
.C(n_962),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1106),
.B(n_1147),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1111),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1114),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1000),
.B(n_1025),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_L g1315 ( 
.A(n_1140),
.B(n_1170),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1114),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1150),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1119),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1119),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1138),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1117),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1138),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1018),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1097),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1070),
.B(n_964),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1156),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1222),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1268),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1187),
.B(n_1086),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1261),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1193),
.B(n_1083),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1261),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1284),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1284),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1285),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1285),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1212),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1287),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1287),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1291),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1268),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_R g1342 ( 
.A(n_1171),
.B(n_1130),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1275),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1200),
.B(n_1112),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1317),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1274),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1233),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1213),
.Y(n_1348)
);

XOR2x2_ASAP7_75t_L g1349 ( 
.A(n_1231),
.B(n_1128),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1215),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1291),
.Y(n_1351)
);

XOR2xp5_ASAP7_75t_L g1352 ( 
.A(n_1243),
.B(n_756),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1297),
.Y(n_1353)
);

NOR2xp67_ASAP7_75t_L g1354 ( 
.A(n_1184),
.B(n_1076),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1178),
.B(n_1028),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1223),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1297),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1265),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1308),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1304),
.Y(n_1360)
);

XNOR2xp5_ASAP7_75t_L g1361 ( 
.A(n_1304),
.B(n_761),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1266),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1250),
.B(n_955),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1269),
.B(n_966),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1270),
.B(n_1044),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1308),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1312),
.Y(n_1367)
);

BUFx8_ASAP7_75t_L g1368 ( 
.A(n_1281),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1312),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1321),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1273),
.Y(n_1371)
);

XOR2xp5_ASAP7_75t_L g1372 ( 
.A(n_1221),
.B(n_764),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_SL g1373 ( 
.A(n_1235),
.B(n_777),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1185),
.B(n_1060),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1321),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1191),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1278),
.B(n_1272),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1211),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1191),
.Y(n_1379)
);

INVxp33_ASAP7_75t_L g1380 ( 
.A(n_1202),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1262),
.B(n_1016),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1210),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1198),
.B(n_1051),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1210),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1194),
.B(n_1157),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1226),
.B(n_1069),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1208),
.B(n_1225),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1292),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1214),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1214),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1218),
.Y(n_1391)
);

XOR2xp5_ASAP7_75t_L g1392 ( 
.A(n_1252),
.B(n_778),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1218),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1260),
.B(n_1091),
.Y(n_1394)
);

XOR2xp5_ASAP7_75t_L g1395 ( 
.A(n_1314),
.B(n_782),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1220),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1292),
.Y(n_1397)
);

INVxp33_ASAP7_75t_L g1398 ( 
.A(n_1325),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1281),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1220),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_SL g1401 ( 
.A(n_1251),
.B(n_785),
.Y(n_1401)
);

BUFx5_ASAP7_75t_L g1402 ( 
.A(n_1172),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1228),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1251),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1241),
.B(n_1085),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1294),
.B(n_1127),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1228),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_SL g1408 ( 
.A(n_1255),
.B(n_798),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1248),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1248),
.Y(n_1410)
);

CKINVDCx16_ASAP7_75t_R g1411 ( 
.A(n_1255),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1256),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_SL g1413 ( 
.A(n_1199),
.B(n_806),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1256),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1298),
.Y(n_1415)
);

XNOR2xp5_ASAP7_75t_L g1416 ( 
.A(n_1311),
.B(n_812),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1298),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1302),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1302),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1229),
.Y(n_1420)
);

NAND2xp33_ASAP7_75t_SL g1421 ( 
.A(n_1323),
.B(n_1039),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1289),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1293),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1296),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1280),
.B(n_1088),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1299),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1282),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1306),
.B(n_1136),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1180),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1283),
.Y(n_1430)
);

BUFx5_ASAP7_75t_L g1431 ( 
.A(n_1172),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1286),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1288),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1224),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1263),
.B(n_1124),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1254),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1173),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1264),
.B(n_1020),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1246),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1271),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1279),
.Y(n_1441)
);

XOR2x2_ASAP7_75t_L g1442 ( 
.A(n_1258),
.B(n_1128),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1316),
.B(n_1021),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1217),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1316),
.B(n_1126),
.Y(n_1445)
);

XOR2xp5_ASAP7_75t_L g1446 ( 
.A(n_1186),
.B(n_820),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1230),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1234),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1232),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1237),
.Y(n_1450)
);

INVxp33_ASAP7_75t_L g1451 ( 
.A(n_1325),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1238),
.Y(n_1452)
);

NOR2x2_ASAP7_75t_L g1453 ( 
.A(n_1349),
.B(n_1437),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1381),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1374),
.B(n_1324),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1330),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1347),
.B(n_1182),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1332),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1387),
.A2(n_1236),
.B1(n_1219),
.B2(n_1179),
.C(n_1315),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1383),
.A2(n_1295),
.B1(n_1249),
.B2(n_1099),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1365),
.A2(n_1394),
.B1(n_1444),
.B2(n_1385),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1328),
.B(n_1188),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1381),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1333),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1395),
.A2(n_1174),
.B1(n_1075),
.B2(n_1065),
.C(n_849),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1406),
.B(n_1239),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1438),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1428),
.B(n_822),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1405),
.B(n_1249),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1425),
.B(n_1249),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1331),
.B(n_1115),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1377),
.B(n_1249),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1334),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1363),
.B(n_825),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_SL g1475 ( 
.A(n_1327),
.B(n_835),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1335),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1364),
.A2(n_847),
.B1(n_851),
.B2(n_846),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1354),
.B(n_1239),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1415),
.A2(n_1099),
.B1(n_1108),
.B2(n_1087),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1438),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1336),
.B(n_1092),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1341),
.B(n_1190),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1338),
.B(n_1121),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1339),
.B(n_1122),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1340),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1417),
.A2(n_1257),
.B(n_1196),
.C(n_1090),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1351),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1337),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1344),
.B(n_1239),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1378),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_1404),
.B(n_1310),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1353),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1378),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1357),
.B(n_1142),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1359),
.B(n_1152),
.Y(n_1495)
);

AO22x1_ASAP7_75t_L g1496 ( 
.A1(n_1380),
.A2(n_1004),
.B1(n_1169),
.B2(n_1132),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1448),
.B(n_1159),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1378),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1366),
.B(n_1168),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1367),
.B(n_1276),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1348),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1355),
.B(n_1134),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1421),
.A2(n_892),
.B1(n_844),
.B2(n_848),
.C(n_852),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_SL g1504 ( 
.A1(n_1418),
.A2(n_1419),
.B(n_1370),
.C(n_1375),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1435),
.B(n_1144),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1386),
.B(n_1145),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1350),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1445),
.B(n_1192),
.Y(n_1508)
);

AND2x6_ASAP7_75t_SL g1509 ( 
.A(n_1329),
.B(n_1303),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1343),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1398),
.B(n_1146),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1369),
.B(n_1173),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1373),
.B(n_1402),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1451),
.B(n_1158),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1376),
.B(n_1175),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1356),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1379),
.A2(n_1160),
.B1(n_1108),
.B2(n_1087),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1382),
.A2(n_1175),
.B(n_1176),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1402),
.B(n_1290),
.Y(n_1519)
);

AND2x6_ASAP7_75t_SL g1520 ( 
.A(n_1372),
.B(n_1209),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1384),
.B(n_1024),
.Y(n_1521)
);

OR2x6_ASAP7_75t_SL g1522 ( 
.A(n_1399),
.B(n_965),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1402),
.B(n_1290),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1389),
.B(n_1031),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1390),
.B(n_1277),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1391),
.A2(n_1189),
.B(n_1240),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1393),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1396),
.A2(n_1244),
.B1(n_1247),
.B2(n_1245),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1400),
.A2(n_1259),
.B1(n_1253),
.B2(n_1242),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1403),
.A2(n_1195),
.B1(n_1253),
.B2(n_1242),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1407),
.A2(n_1267),
.B1(n_1183),
.B2(n_1300),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1409),
.B(n_1183),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1358),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1420),
.B(n_1301),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1402),
.B(n_1267),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1345),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1410),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1431),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1342),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1412),
.A2(n_1318),
.B1(n_1305),
.B2(n_1309),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1461),
.B(n_1414),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1455),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1500),
.B(n_1431),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1496),
.B(n_1443),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1508),
.B(n_1434),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1431),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1456),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1534),
.B(n_1436),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1481),
.B(n_1431),
.Y(n_1549)
);

BUFx4f_ASAP7_75t_L g1550 ( 
.A(n_1493),
.Y(n_1550)
);

AND2x6_ASAP7_75t_L g1551 ( 
.A(n_1537),
.B(n_1440),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1453),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1508),
.B(n_1441),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1537),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1527),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1510),
.B(n_1388),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_SL g1557 ( 
.A(n_1468),
.B(n_1411),
.C(n_1416),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1483),
.B(n_1422),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1471),
.A2(n_1401),
.B1(n_1408),
.B2(n_1413),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1484),
.B(n_1423),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1493),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1539),
.Y(n_1562)
);

AND2x6_ASAP7_75t_L g1563 ( 
.A(n_1537),
.B(n_1458),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1536),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1462),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1464),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1474),
.A2(n_1346),
.B1(n_1439),
.B2(n_1429),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1493),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1469),
.B(n_1470),
.Y(n_1569)
);

AND2x2_ASAP7_75t_SL g1570 ( 
.A(n_1475),
.B(n_1442),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1454),
.B(n_1463),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1467),
.B(n_1480),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1457),
.B(n_1452),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1462),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1473),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1502),
.B(n_1361),
.C(n_670),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1476),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1477),
.B(n_1352),
.Y(n_1578)
);

AND3x1_ASAP7_75t_L g1579 ( 
.A(n_1465),
.B(n_1313),
.C(n_1307),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1538),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1534),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1472),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1485),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1494),
.B(n_1392),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1487),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1492),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1512),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1495),
.B(n_1426),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1499),
.B(n_1450),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1490),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1515),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_SL g1592 ( 
.A(n_1505),
.B(n_1397),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1511),
.B(n_1446),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1457),
.B(n_1427),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1549),
.A2(n_1538),
.B(n_1513),
.Y(n_1595)
);

AO31x2_ASAP7_75t_L g1596 ( 
.A1(n_1546),
.A2(n_1486),
.A3(n_1525),
.B(n_1518),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1587),
.B(n_1521),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1543),
.A2(n_1459),
.B(n_1460),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1569),
.A2(n_1526),
.B(n_1504),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1541),
.A2(n_1478),
.B(n_1535),
.Y(n_1600)
);

BUFx12f_ASAP7_75t_L g1601 ( 
.A(n_1564),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1550),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1580),
.A2(n_1466),
.B(n_1479),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1591),
.B(n_1506),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1558),
.B(n_1524),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1580),
.A2(n_1523),
.B(n_1519),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1547),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1554),
.A2(n_1532),
.B(n_1517),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1554),
.A2(n_1579),
.B(n_1528),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1542),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1560),
.A2(n_1529),
.B(n_1489),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1555),
.A2(n_1501),
.B(n_1488),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1514),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1588),
.A2(n_1540),
.B(n_1432),
.Y(n_1616)
);

BUFx8_ASAP7_75t_SL g1617 ( 
.A(n_1552),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1585),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1589),
.A2(n_1516),
.B(n_1507),
.Y(n_1619)
);

AO31x2_ASAP7_75t_L g1620 ( 
.A1(n_1575),
.A2(n_1433),
.A3(n_1447),
.B(n_1430),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

AO32x1_ASAP7_75t_L g1622 ( 
.A1(n_1583),
.A2(n_1449),
.A3(n_968),
.B1(n_857),
.B2(n_860),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1571),
.B(n_1498),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1556),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1572),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1573),
.Y(n_1627)
);

NAND2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1590),
.B(n_1181),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1593),
.B(n_1491),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1531),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1562),
.Y(n_1631)
);

AND3x4_ASAP7_75t_L g1632 ( 
.A(n_1557),
.B(n_1520),
.C(n_1522),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1576),
.A2(n_1371),
.B(n_1424),
.C(n_1362),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1601),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1598),
.A2(n_1559),
.B(n_1592),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1631),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1607),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1608),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1595),
.A2(n_1605),
.B(n_1604),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1597),
.A2(n_1614),
.B(n_1633),
.C(n_1578),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1597),
.B(n_1567),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1612),
.A2(n_1570),
.B(n_1545),
.C(n_1553),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1615),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1618),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1625),
.B(n_1594),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1599),
.A2(n_1544),
.B(n_1582),
.Y(n_1646)
);

AO22x2_ASAP7_75t_L g1647 ( 
.A1(n_1632),
.A2(n_1553),
.B1(n_1545),
.B2(n_1565),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1621),
.Y(n_1648)
);

AOI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1603),
.A2(n_1177),
.B(n_1544),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1600),
.A2(n_1530),
.B(n_1320),
.Y(n_1650)
);

AO31x2_ASAP7_75t_L g1651 ( 
.A1(n_1619),
.A2(n_856),
.A3(n_861),
.B(n_854),
.Y(n_1651)
);

BUFx12f_ASAP7_75t_L g1652 ( 
.A(n_1602),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1611),
.A2(n_1503),
.B1(n_889),
.B2(n_891),
.C(n_862),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1602),
.B(n_1590),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1629),
.B(n_1581),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1622),
.A2(n_868),
.A3(n_869),
.B(n_865),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1612),
.A2(n_1322),
.B(n_1319),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1616),
.A2(n_1563),
.B(n_1548),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1609),
.A2(n_1326),
.B(n_1201),
.Y(n_1659)
);

BUFx12f_ASAP7_75t_L g1660 ( 
.A(n_1624),
.Y(n_1660)
);

NAND3x1_ASAP7_75t_L g1661 ( 
.A(n_1626),
.B(n_1368),
.C(n_1117),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1620),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1627),
.B(n_1574),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1620),
.Y(n_1664)
);

AO31x2_ASAP7_75t_L g1665 ( 
.A1(n_1622),
.A2(n_872),
.A3(n_876),
.B(n_871),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1616),
.A2(n_882),
.B(n_881),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1628),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1631),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1606),
.A2(n_1203),
.B(n_1197),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1630),
.A2(n_1360),
.B1(n_1548),
.B2(n_1551),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1610),
.A2(n_1204),
.B(n_1181),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1613),
.A2(n_1551),
.B(n_1563),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1617),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1623),
.A2(n_1551),
.B1(n_1563),
.B2(n_1368),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1622),
.A2(n_1563),
.B(n_1551),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1637),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1638),
.Y(n_1677)
);

OAI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1641),
.A2(n_1623),
.B1(n_873),
.B2(n_1590),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1668),
.B(n_1620),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1635),
.A2(n_885),
.B(n_884),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1636),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1652),
.Y(n_1682)
);

CKINVDCx6p67_ASAP7_75t_R g1683 ( 
.A(n_1673),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1662),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1643),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1647),
.A2(n_1646),
.B1(n_1658),
.B2(n_1655),
.Y(n_1686)
);

CKINVDCx11_ASAP7_75t_R g1687 ( 
.A(n_1660),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1644),
.Y(n_1688)
);

BUFx8_ASAP7_75t_L g1689 ( 
.A(n_1634),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1645),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1647),
.A2(n_1205),
.B1(n_1206),
.B2(n_1078),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1663),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1648),
.B(n_1561),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1670),
.A2(n_1568),
.B1(n_947),
.B2(n_1482),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1674),
.A2(n_1482),
.B1(n_669),
.B2(n_675),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1639),
.A2(n_1205),
.B1(n_1206),
.B2(n_1084),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1654),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1664),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1653),
.A2(n_1666),
.B1(n_1657),
.B2(n_1650),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1649),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1651),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1651),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1667),
.A2(n_1063),
.B1(n_1078),
.B2(n_1084),
.Y(n_1703)
);

CKINVDCx11_ASAP7_75t_R g1704 ( 
.A(n_1654),
.Y(n_1704)
);

INVx6_ASAP7_75t_L g1705 ( 
.A(n_1667),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1661),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1642),
.A2(n_888),
.B1(n_893),
.B2(n_894),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1672),
.A2(n_1061),
.B1(n_1063),
.B2(n_1162),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1675),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1640),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1669),
.A2(n_1061),
.B1(n_1164),
.B2(n_1156),
.Y(n_1711)
);

CKINVDCx6p67_ASAP7_75t_R g1712 ( 
.A(n_1656),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1656),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1659),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1665),
.B(n_1227),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1671),
.Y(n_1717)
);

CKINVDCx16_ASAP7_75t_R g1718 ( 
.A(n_1690),
.Y(n_1718)
);

OAI21xp33_ASAP7_75t_SL g1719 ( 
.A1(n_1691),
.A2(n_902),
.B(n_896),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1681),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1676),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1692),
.Y(n_1722)
);

BUFx12f_ASAP7_75t_L g1723 ( 
.A(n_1687),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1677),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1704),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1684),
.Y(n_1726)
);

OR2x6_ASAP7_75t_L g1727 ( 
.A(n_1701),
.B(n_1596),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1679),
.B(n_1596),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1698),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1710),
.A2(n_907),
.B(n_903),
.Y(n_1730)
);

AO21x2_ASAP7_75t_L g1731 ( 
.A1(n_1702),
.A2(n_913),
.B(n_1596),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1686),
.B(n_2),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1688),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1685),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1707),
.A2(n_1164),
.B1(n_1162),
.B2(n_1055),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1713),
.Y(n_1737)
);

BUFx12f_ASAP7_75t_L g1738 ( 
.A(n_1689),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1714),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1693),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1717),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1716),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1680),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1712),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1709),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1715),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1706),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1680),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1699),
.B(n_4),
.Y(n_1750)
);

INVx5_ASAP7_75t_SL g1751 ( 
.A(n_1683),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1707),
.B(n_5),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1697),
.B(n_10),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1705),
.B(n_1708),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1689),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1705),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1682),
.Y(n_1757)
);

INVxp33_ASAP7_75t_L g1758 ( 
.A(n_1694),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1682),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1682),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1694),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1695),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1678),
.B(n_1067),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1696),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1711),
.Y(n_1765)
);

AO21x2_ASAP7_75t_L g1766 ( 
.A1(n_1703),
.A2(n_1509),
.B(n_12),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1710),
.A2(n_1176),
.B(n_1133),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1676),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1721),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1739),
.A2(n_12),
.B(n_13),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1094),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1735),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1735),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1746),
.B(n_13),
.Y(n_1774)
);

AO21x2_ASAP7_75t_L g1775 ( 
.A1(n_1744),
.A2(n_14),
.B(n_15),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1724),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1768),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1729),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1739),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1749),
.B(n_16),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1720),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1733),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1742),
.B(n_16),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1761),
.B(n_17),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1749),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1761),
.B(n_18),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1745),
.B(n_19),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1734),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1725),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1747),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1742),
.B(n_1139),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1741),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1757),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1725),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1725),
.Y(n_1798)
);

OA21x2_ASAP7_75t_L g1799 ( 
.A1(n_1743),
.A2(n_20),
.B(n_22),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1747),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1727),
.B(n_20),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1740),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1727),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1743),
.B(n_23),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1727),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1747),
.Y(n_1806)
);

OAI21xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1750),
.A2(n_23),
.B(n_24),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1748),
.Y(n_1808)
);

OAI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1748),
.A2(n_1216),
.B(n_1207),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1776),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1777),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1788),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1782),
.B(n_1758),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1778),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1792),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1805),
.B(n_1757),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1782),
.B(n_1718),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1788),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1779),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1788),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1805),
.B(n_1760),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1807),
.A2(n_1732),
.B(n_1750),
.C(n_1762),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1803),
.B(n_1760),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1799),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1787),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1798),
.B(n_1802),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1793),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1772),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1780),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1725),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1784),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1780),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1795),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1793),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1797),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1836),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1814),
.B(n_1816),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1826),
.B(n_1771),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1837),
.B(n_1801),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1810),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1829),
.B(n_1793),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1838),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1820),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1811),
.B(n_1783),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1832),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1818),
.B(n_1800),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1812),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1815),
.Y(n_1853)
);

NAND2x1_ASAP7_75t_L g1854 ( 
.A(n_1819),
.B(n_1770),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1820),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1821),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1838),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1828),
.B(n_1800),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1817),
.B(n_1806),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1817),
.B(n_1806),
.Y(n_1861)
);

BUFx2_ASAP7_75t_SL g1862 ( 
.A(n_1833),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1834),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1806),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1841),
.B(n_1826),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1862),
.B(n_1817),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1842),
.B(n_1823),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1844),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1852),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1853),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1857),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1823),
.Y(n_1872)
);

CKINVDCx16_ASAP7_75t_R g1873 ( 
.A(n_1847),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1858),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1863),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1839),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1849),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1850),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1847),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1850),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1842),
.B(n_1823),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1848),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1851),
.B(n_1825),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1848),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1840),
.B(n_1856),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1860),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1864),
.B(n_1801),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1856),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1854),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1843),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1861),
.B(n_1846),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1846),
.B(n_1855),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1843),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1859),
.B(n_1827),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1855),
.B(n_1825),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1845),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1873),
.B(n_1864),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1878),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1878),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1879),
.B(n_1723),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1885),
.B(n_1804),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1868),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1867),
.B(n_1845),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1881),
.B(n_1825),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1869),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1877),
.B(n_1832),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1879),
.B(n_1723),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1872),
.B(n_1755),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1874),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1887),
.B(n_1781),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1870),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1872),
.B(n_1755),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1887),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1871),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1875),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1865),
.B(n_1824),
.Y(n_1916)
);

NAND2xp33_ASAP7_75t_SL g1917 ( 
.A(n_1897),
.B(n_1866),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1900),
.B(n_1880),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1909),
.B(n_1887),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1908),
.B(n_1866),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1912),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1900),
.B(n_1775),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1907),
.B(n_1775),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1907),
.B(n_1738),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1913),
.B(n_1876),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1898),
.B(n_1890),
.Y(n_1926)
);

OAI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1916),
.A2(n_1758),
.B1(n_1886),
.B2(n_1896),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1899),
.B(n_1893),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1910),
.B(n_1891),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1910),
.B(n_1891),
.Y(n_1930)
);

NOR4xp25_ASAP7_75t_SL g1931 ( 
.A(n_1902),
.B(n_1889),
.C(n_1882),
.D(n_1835),
.Y(n_1931)
);

INVxp67_ASAP7_75t_SL g1932 ( 
.A(n_1918),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1920),
.B(n_1903),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1922),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1924),
.B(n_1738),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1929),
.B(n_1901),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1921),
.B(n_1905),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1926),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1917),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1919),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1939),
.B(n_1930),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1937),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1936),
.Y(n_1943)
);

AOI21xp33_ASAP7_75t_L g1944 ( 
.A1(n_1932),
.A2(n_1927),
.B(n_1923),
.Y(n_1944)
);

NAND4xp25_ASAP7_75t_L g1945 ( 
.A(n_1940),
.B(n_1928),
.C(n_1925),
.D(n_1914),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1933),
.B(n_1911),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1938),
.B(n_1915),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1941),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1943),
.A2(n_1934),
.B1(n_1931),
.B2(n_1935),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1946),
.B(n_1935),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1947),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1944),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1952),
.A2(n_1945),
.B1(n_1942),
.B2(n_1906),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1948),
.B(n_1950),
.Y(n_1954)
);

AOI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1949),
.A2(n_1774),
.B(n_1790),
.C(n_1753),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1954),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1955),
.Y(n_1957)
);

NOR3xp33_ASAP7_75t_L g1958 ( 
.A(n_1956),
.B(n_1951),
.C(n_1953),
.Y(n_1958)
);

NAND4xp25_ASAP7_75t_L g1959 ( 
.A(n_1957),
.B(n_1730),
.C(n_1767),
.D(n_1786),
.Y(n_1959)
);

NAND2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1956),
.B(n_1759),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1958),
.A2(n_1906),
.B(n_1789),
.C(n_1763),
.Y(n_1961)
);

NAND4xp25_ASAP7_75t_L g1962 ( 
.A(n_1959),
.B(n_1759),
.C(n_1722),
.D(n_1752),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1960),
.B(n_1766),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1961),
.B(n_1751),
.Y(n_1964)
);

NOR4xp25_ASAP7_75t_L g1965 ( 
.A(n_1962),
.B(n_1888),
.C(n_1884),
.D(n_1794),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1965),
.B(n_1884),
.Y(n_1966)
);

XNOR2x1_ASAP7_75t_L g1967 ( 
.A(n_1964),
.B(n_24),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1963),
.B(n_1904),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_R g1969 ( 
.A(n_1963),
.B(n_25),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1968),
.B(n_1888),
.Y(n_1970)
);

AND4x1_ASAP7_75t_L g1971 ( 
.A(n_1967),
.B(n_1751),
.C(n_1752),
.D(n_27),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1966),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1969),
.B(n_1892),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1973),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1971),
.B(n_1766),
.Y(n_1975)
);

NOR4xp75_ASAP7_75t_L g1976 ( 
.A(n_1970),
.B(n_1759),
.C(n_26),
.D(n_27),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1973),
.A2(n_1799),
.B1(n_1751),
.B2(n_1781),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1973),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1973),
.Y(n_1979)
);

BUFx8_ASAP7_75t_L g1980 ( 
.A(n_1972),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1973),
.A2(n_1892),
.B1(n_1781),
.B2(n_1799),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1975),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1976),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1978),
.A2(n_1895),
.B1(n_1756),
.B2(n_1785),
.Y(n_1984)
);

AO22x2_ASAP7_75t_L g1985 ( 
.A1(n_1979),
.A2(n_1756),
.B1(n_1894),
.B2(n_1883),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1980),
.Y(n_1986)
);

INVx3_ASAP7_75t_L g1987 ( 
.A(n_1977),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1981),
.A2(n_1719),
.B1(n_1770),
.B2(n_1831),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1974),
.A2(n_1736),
.B1(n_1813),
.B2(n_1770),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1974),
.A2(n_1736),
.B1(n_1813),
.B2(n_1819),
.Y(n_1990)
);

OAI22x1_ASAP7_75t_L g1991 ( 
.A1(n_1974),
.A2(n_1822),
.B1(n_1754),
.B2(n_32),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1974),
.A2(n_1822),
.B1(n_1211),
.B2(n_1791),
.Y(n_1992)
);

AO22x1_ASAP7_75t_L g1993 ( 
.A1(n_1980),
.A2(n_25),
.B1(n_30),
.B2(n_33),
.Y(n_1993)
);

OAI22x1_ASAP7_75t_L g1994 ( 
.A1(n_1974),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_1994)
);

OAI22x1_ASAP7_75t_L g1995 ( 
.A1(n_1974),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1974),
.A2(n_1207),
.B1(n_1216),
.B2(n_1211),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1974),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1975),
.Y(n_1998)
);

AO22x2_ASAP7_75t_L g1999 ( 
.A1(n_1974),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1974),
.A2(n_1830),
.B1(n_1765),
.B2(n_1808),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1975),
.Y(n_2001)
);

AOI22x1_ASAP7_75t_L g2002 ( 
.A1(n_1974),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_2002)
);

AO22x2_ASAP7_75t_L g2003 ( 
.A1(n_1974),
.A2(n_48),
.B1(n_51),
.B2(n_1830),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_2003),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1991),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1993),
.B(n_55),
.Y(n_2006)
);

AND3x2_ASAP7_75t_L g2007 ( 
.A(n_1986),
.B(n_60),
.C(n_66),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1983),
.A2(n_1765),
.B1(n_1764),
.B2(n_73),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1997),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1999),
.Y(n_2010)
);

NAND3x1_ASAP7_75t_L g2011 ( 
.A(n_1982),
.B(n_71),
.C(n_72),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1987),
.B(n_75),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1994),
.B(n_76),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_SL g2014 ( 
.A1(n_1995),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1998),
.A2(n_1773),
.B1(n_88),
.B2(n_89),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1984),
.A2(n_86),
.B1(n_93),
.B2(n_102),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_2002),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2001),
.B(n_104),
.Y(n_2018)
);

OA21x2_ASAP7_75t_L g2019 ( 
.A1(n_1996),
.A2(n_1809),
.B(n_110),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1985),
.A2(n_1731),
.B1(n_114),
.B2(n_115),
.Y(n_2020)
);

AO21x2_ASAP7_75t_L g2021 ( 
.A1(n_1990),
.A2(n_2000),
.B(n_1988),
.Y(n_2021)
);

INVx3_ASAP7_75t_SL g2022 ( 
.A(n_1992),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_SL g2023 ( 
.A1(n_1989),
.A2(n_109),
.B1(n_122),
.B2(n_130),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_SL g2024 ( 
.A1(n_1983),
.A2(n_134),
.B1(n_140),
.B2(n_145),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1986),
.B(n_151),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1986),
.Y(n_2026)
);

OA22x2_ASAP7_75t_L g2027 ( 
.A1(n_1991),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1993),
.B(n_162),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1986),
.Y(n_2029)
);

NAND2x1p5_ASAP7_75t_L g2030 ( 
.A(n_1986),
.B(n_167),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2026),
.Y(n_2031)
);

NAND4xp25_ASAP7_75t_L g2032 ( 
.A(n_2029),
.B(n_170),
.C(n_176),
.D(n_177),
.Y(n_2032)
);

AOI221x1_ASAP7_75t_L g2033 ( 
.A1(n_2010),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.C(n_186),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_2027),
.A2(n_191),
.B(n_192),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_2011),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2005),
.A2(n_196),
.B(n_198),
.Y(n_2036)
);

AO21x2_ASAP7_75t_L g2037 ( 
.A1(n_2018),
.A2(n_199),
.B(n_208),
.Y(n_2037)
);

INVx3_ASAP7_75t_L g2038 ( 
.A(n_2009),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2006),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2028),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_2012),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_SL g2042 ( 
.A1(n_2004),
.A2(n_2017),
.B1(n_2013),
.B2(n_2030),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_2009),
.A2(n_1731),
.B1(n_222),
.B2(n_224),
.Y(n_2043)
);

OAI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_2020),
.A2(n_219),
.B(n_229),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2007),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2025),
.Y(n_2046)
);

OAI32xp33_ASAP7_75t_L g2047 ( 
.A1(n_2016),
.A2(n_239),
.A3(n_242),
.B1(n_249),
.B2(n_259),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2014),
.A2(n_261),
.B1(n_262),
.B2(n_265),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_2035),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2037),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_2034),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_2038),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2031),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_2045),
.A2(n_2008),
.B1(n_2023),
.B2(n_2015),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_2048),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_2046),
.Y(n_2056)
);

BUFx6f_ASAP7_75t_L g2057 ( 
.A(n_2039),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2042),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_2040),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2044),
.Y(n_2060)
);

CKINVDCx20_ASAP7_75t_R g2061 ( 
.A(n_2036),
.Y(n_2061)
);

BUFx2_ASAP7_75t_L g2062 ( 
.A(n_2032),
.Y(n_2062)
);

NAND2xp33_ASAP7_75t_R g2063 ( 
.A(n_2033),
.B(n_2019),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2041),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2049),
.B(n_2021),
.Y(n_2065)
);

OR2x6_ASAP7_75t_L g2066 ( 
.A(n_2050),
.B(n_2024),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2058),
.B(n_2022),
.Y(n_2067)
);

AOI21xp33_ASAP7_75t_SL g2068 ( 
.A1(n_2053),
.A2(n_2047),
.B(n_2043),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2056),
.B(n_270),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_2052),
.B(n_272),
.Y(n_2070)
);

XNOR2xp5_ASAP7_75t_L g2071 ( 
.A(n_2059),
.B(n_390),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2051),
.A2(n_281),
.B(n_284),
.Y(n_2072)
);

NAND2x1p5_ASAP7_75t_L g2073 ( 
.A(n_2057),
.B(n_286),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2063),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2055),
.B(n_289),
.Y(n_2075)
);

AO22x2_ASAP7_75t_L g2076 ( 
.A1(n_2065),
.A2(n_2064),
.B1(n_2060),
.B2(n_2061),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2074),
.A2(n_2054),
.B1(n_2057),
.B2(n_2062),
.Y(n_2077)
);

OAI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2069),
.A2(n_290),
.B1(n_291),
.B2(n_293),
.Y(n_2078)
);

OAI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2067),
.A2(n_294),
.B1(n_295),
.B2(n_303),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_2075),
.A2(n_304),
.B1(n_307),
.B2(n_312),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2076),
.B(n_2068),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2077),
.Y(n_2082)
);

OAI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2079),
.A2(n_2066),
.B(n_2072),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2081),
.A2(n_2066),
.B(n_2073),
.Y(n_2084)
);

OAI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_2084),
.A2(n_2082),
.B1(n_2083),
.B2(n_2070),
.Y(n_2085)
);

AOI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2085),
.A2(n_2078),
.B(n_2071),
.C(n_2080),
.Y(n_2086)
);


endmodule