module fake_jpeg_3304_n_687 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_687);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_687;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_352;
wire n_150;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_70),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_63),
.Y(n_193)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_8),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_65),
.B(n_36),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_66),
.Y(n_170)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_33),
.B(n_8),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_14),
.Y(n_155)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_75),
.Y(n_198)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_79),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_90),
.Y(n_148)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_8),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_94),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_100),
.Y(n_230)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_103),
.Y(n_211)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_9),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_115),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_114),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_9),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

BUFx4f_ASAP7_75t_SL g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_58),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_28),
.B(n_9),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_13),
.Y(n_167)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_34),
.Y(n_130)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_34),
.Y(n_131)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_63),
.B(n_31),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_140),
.B(n_146),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_46),
.B1(n_41),
.B2(n_52),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_142),
.A2(n_165),
.B1(n_214),
.B2(n_58),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_81),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_155),
.B(n_168),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_51),
.B1(n_55),
.B2(n_31),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_156),
.A2(n_166),
.B1(n_172),
.B2(n_185),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_80),
.A2(n_41),
.B1(n_46),
.B2(n_52),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_159),
.A2(n_229),
.B1(n_54),
.B2(n_1),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_86),
.A2(n_46),
.B1(n_52),
.B2(n_41),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_103),
.A2(n_51),
.B1(n_55),
.B2(n_31),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_167),
.B(n_195),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_44),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_105),
.A2(n_48),
.B1(n_55),
.B2(n_28),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_48),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_174),
.B(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_26),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_184),
.B(n_222),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_72),
.A2(n_48),
.B1(n_52),
.B2(n_46),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_77),
.B(n_53),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_94),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_192),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_87),
.B(n_44),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_201),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_78),
.B(n_27),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_84),
.B(n_41),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_98),
.B(n_53),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_223),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_111),
.A2(n_37),
.B1(n_44),
.B2(n_36),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_125),
.B(n_37),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_121),
.B(n_35),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_127),
.B(n_53),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_232),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_95),
.A2(n_36),
.B1(n_37),
.B2(n_27),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_131),
.B(n_45),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_100),
.B(n_45),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_58),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_234),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_235),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_237),
.Y(n_336)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_240),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_241),
.A2(n_244),
.B1(n_276),
.B2(n_283),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_165),
.A2(n_126),
.B1(n_122),
.B2(n_117),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_242),
.A2(n_264),
.B1(n_273),
.B2(n_278),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_147),
.A2(n_125),
.B(n_45),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_243),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_195),
.A2(n_116),
.B1(n_113),
.B2(n_110),
.Y(n_244)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_250),
.Y(n_350)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_253),
.Y(n_358)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_151),
.Y(n_256)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_156),
.A2(n_106),
.B1(n_27),
.B2(n_35),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_SL g341 ( 
.A1(n_258),
.A2(n_263),
.B(n_268),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_151),
.A2(n_35),
.B1(n_120),
.B2(n_38),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_209),
.B1(n_134),
.B2(n_133),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g382 ( 
.A(n_266),
.B(n_312),
.C(n_315),
.Y(n_382)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_151),
.A2(n_38),
.B1(n_22),
.B2(n_30),
.Y(n_268)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_269),
.Y(n_368)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_270),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_149),
.B(n_22),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_291),
.Y(n_325)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_154),
.Y(n_272)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_272),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_184),
.A2(n_38),
.B1(n_22),
.B2(n_30),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_148),
.B(n_9),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_275),
.B(n_309),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

INVx4_ASAP7_75t_SL g354 ( 
.A(n_277),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_182),
.A2(n_54),
.B1(n_7),
.B2(n_10),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_160),
.Y(n_280)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_162),
.A2(n_54),
.B1(n_7),
.B2(n_13),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_161),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_199),
.A2(n_54),
.B1(n_7),
.B2(n_13),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_287),
.A2(n_294),
.B1(n_305),
.B2(n_183),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_185),
.A2(n_54),
.B1(n_6),
.B2(n_15),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_288),
.A2(n_313),
.B1(n_316),
.B2(n_318),
.Y(n_366)
);

BUFx16f_ASAP7_75t_L g289 ( 
.A(n_171),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_289),
.Y(n_360)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_190),
.Y(n_290)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_145),
.B(n_6),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_292),
.B(n_298),
.Y(n_365)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_136),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_299),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_170),
.A2(n_54),
.B1(n_19),
.B2(n_18),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_139),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_300),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_135),
.A2(n_19),
.B(n_17),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_138),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_143),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_303),
.Y(n_355)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_210),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_306),
.Y(n_337)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_180),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_304),
.B(n_307),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_152),
.A2(n_17),
.B1(n_15),
.B2(n_2),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_138),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_157),
.Y(n_309)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_139),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_216),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_157),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_166),
.A2(n_17),
.B1(n_15),
.B2(n_2),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_203),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_172),
.B1(n_231),
.B2(n_221),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_225),
.B(n_0),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_164),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_181),
.B(n_0),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_164),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_319),
.B(n_321),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_169),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_320),
.B(n_250),
.Y(n_383)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_175),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_323),
.A2(n_327),
.B1(n_339),
.B2(n_342),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_241),
.A2(n_257),
.B1(n_242),
.B2(n_251),
.Y(n_327)
);

AND2x4_ASAP7_75t_SL g329 ( 
.A(n_255),
.B(n_183),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_329),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_338),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_248),
.A2(n_224),
.B1(n_175),
.B2(n_173),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_248),
.A2(n_243),
.B1(n_260),
.B2(n_296),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_340),
.A2(n_348),
.B1(n_370),
.B2(n_278),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_257),
.A2(n_224),
.B1(n_173),
.B2(n_176),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_254),
.A2(n_230),
.B1(n_217),
.B2(n_211),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_252),
.B(n_169),
.C(n_204),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_359),
.C(n_235),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_252),
.A2(n_158),
.B(n_178),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_352),
.A2(n_268),
.B(n_263),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_239),
.A2(n_204),
.B1(n_231),
.B2(n_221),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_353),
.A2(n_373),
.B1(n_375),
.B2(n_380),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_245),
.B(n_230),
.C(n_178),
.Y(n_359)
);

AOI32xp33_ASAP7_75t_L g361 ( 
.A1(n_297),
.A2(n_178),
.A3(n_205),
.B1(n_219),
.B2(n_150),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_256),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_290),
.A2(n_137),
.B1(n_202),
.B2(n_194),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_258),
.A2(n_202),
.B1(n_194),
.B2(n_177),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_273),
.A2(n_137),
.B1(n_150),
.B2(n_219),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_244),
.B(n_177),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_379),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_285),
.B(n_0),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_314),
.A2(n_205),
.B1(n_1),
.B2(n_2),
.Y(n_380)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_387),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_390),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_238),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_391),
.B(n_408),
.C(n_422),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_383),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_392),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_334),
.Y(n_435)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_384),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_395),
.B(n_397),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_330),
.B(n_265),
.Y(n_397)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_305),
.B(n_294),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_407),
.B(n_424),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_401),
.B(n_415),
.Y(n_459)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_330),
.B(n_306),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_404),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_351),
.B(n_259),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_300),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_418),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_349),
.A2(n_287),
.B(n_284),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_279),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_412),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_327),
.A2(n_262),
.B1(n_246),
.B2(n_319),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_413),
.A2(n_414),
.B1(n_416),
.B2(n_419),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_333),
.A2(n_377),
.B1(n_378),
.B2(n_366),
.Y(n_414)
);

INVx3_ASAP7_75t_SL g415 ( 
.A(n_354),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_333),
.A2(n_323),
.B1(n_328),
.B2(n_341),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_352),
.A2(n_318),
.B(n_316),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_417),
.A2(n_350),
.B(n_343),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_337),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_366),
.A2(n_269),
.B1(n_247),
.B2(n_307),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_420),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_359),
.B(n_310),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_421),
.B(n_427),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_270),
.C(n_267),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_373),
.A2(n_274),
.B1(n_277),
.B2(n_261),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_423),
.A2(n_426),
.B1(n_434),
.B2(n_336),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_365),
.A2(n_289),
.B(n_298),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_325),
.B(n_311),
.C(n_289),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_350),
.C(n_372),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_353),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_337),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_354),
.A2(n_295),
.B1(n_304),
.B2(n_286),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_428),
.A2(n_432),
.B1(n_332),
.B2(n_367),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_337),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_429),
.Y(n_457)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

AO22x1_ASAP7_75t_L g431 ( 
.A1(n_364),
.A2(n_249),
.B1(n_1),
.B2(n_3),
.Y(n_431)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_431),
.A2(n_369),
.B1(n_332),
.B2(n_356),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_368),
.A2(n_5),
.B1(n_0),
.B2(n_4),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_433),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_364),
.A2(n_4),
.B1(n_322),
.B2(n_324),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_435),
.B(n_437),
.C(n_463),
.Y(n_495)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_334),
.C(n_346),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_436),
.B(n_408),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_358),
.Y(n_437)
);

AO22x1_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_322),
.B1(n_334),
.B2(n_324),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_439),
.B(n_431),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_442),
.A2(n_431),
.B(n_415),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_407),
.A2(n_326),
.B(n_360),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_443),
.A2(n_428),
.B(n_402),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_362),
.B1(n_346),
.B2(n_374),
.Y(n_444)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_444),
.A2(n_464),
.B1(n_477),
.B2(n_415),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_416),
.A2(n_362),
.B1(n_347),
.B2(n_343),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_447),
.B1(n_461),
.B2(n_472),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_389),
.A2(n_347),
.B1(n_343),
.B2(n_374),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_452),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_389),
.A2(n_356),
.B1(n_326),
.B2(n_357),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_401),
.A2(n_369),
.B1(n_331),
.B2(n_372),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_403),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_465),
.B(n_385),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_434),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_466),
.B(n_427),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_336),
.C(n_367),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_474),
.C(n_417),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_469),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_398),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_391),
.B(n_345),
.C(n_4),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_419),
.A2(n_4),
.B1(n_345),
.B2(n_392),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_476),
.Y(n_478)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_462),
.A2(n_413),
.B1(n_398),
.B2(n_426),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_479),
.A2(n_481),
.B1(n_487),
.B2(n_499),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_422),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_480),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_482),
.B(n_454),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_501),
.Y(n_518)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_455),
.Y(n_484)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_484),
.Y(n_527)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_485),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_476),
.A2(n_388),
.B1(n_385),
.B2(n_396),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_386),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_435),
.C(n_454),
.Y(n_526)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_489),
.Y(n_533)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_458),
.Y(n_490)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_491),
.A2(n_492),
.B1(n_493),
.B2(n_498),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_451),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_440),
.A2(n_394),
.B1(n_396),
.B2(n_400),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_424),
.Y(n_496)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_496),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_500),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_441),
.A2(n_423),
.B1(n_405),
.B2(n_397),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_441),
.A2(n_418),
.B1(n_429),
.B2(n_390),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_450),
.B(n_425),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_475),
.B(n_395),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_437),
.B(n_387),
.Y(n_503)
);

INVxp33_ASAP7_75t_SL g555 ( 
.A(n_503),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_457),
.B(n_412),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_508),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_505),
.A2(n_509),
.B(n_496),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_451),
.B(n_399),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_506),
.B(n_449),
.Y(n_550)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_507),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_457),
.B(n_420),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_448),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_511),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_448),
.B(n_430),
.Y(n_511)
);

AO22x1_ASAP7_75t_SL g512 ( 
.A1(n_461),
.A2(n_459),
.B1(n_445),
.B2(n_446),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_512),
.B(n_513),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_453),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_515),
.A2(n_452),
.B1(n_473),
.B2(n_470),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_446),
.B(n_409),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_516),
.Y(n_553)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_517),
.B(n_471),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_526),
.B(n_537),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_481),
.A2(n_460),
.B1(n_459),
.B2(n_447),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_529),
.A2(n_534),
.B1(n_539),
.B2(n_540),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_481),
.A2(n_460),
.B1(n_459),
.B2(n_468),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_493),
.A2(n_468),
.B1(n_466),
.B2(n_439),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_536),
.A2(n_502),
.B1(n_514),
.B2(n_510),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_488),
.B(n_467),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_497),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_478),
.A2(n_439),
.B1(n_469),
.B2(n_463),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_504),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_541),
.B(n_545),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_495),
.B(n_474),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_544),
.C(n_549),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_495),
.B(n_443),
.C(n_442),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_508),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_501),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_546),
.B(n_548),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_511),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_482),
.B(n_473),
.C(n_449),
.Y(n_549)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_550),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_514),
.A2(n_479),
.B1(n_513),
.B2(n_491),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_551),
.A2(n_496),
.B1(n_486),
.B2(n_509),
.Y(n_559)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_554),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_556),
.A2(n_569),
.B1(n_571),
.B2(n_575),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_522),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_558),
.B(n_567),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_559),
.A2(n_576),
.B1(n_552),
.B2(n_529),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_525),
.B(n_500),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_562),
.B(n_555),
.Y(n_594)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_522),
.Y(n_564)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_564),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_537),
.Y(n_591)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_533),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_523),
.A2(n_499),
.B1(n_486),
.B2(n_489),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_533),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_570),
.B(n_577),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_536),
.A2(n_486),
.B1(n_487),
.B2(n_498),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_521),
.B(n_485),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_572),
.B(n_530),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_526),
.B(n_512),
.C(n_505),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_573),
.B(n_578),
.C(n_542),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_520),
.A2(n_512),
.B1(n_516),
.B2(n_484),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_551),
.A2(n_512),
.B1(n_507),
.B2(n_494),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_530),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_543),
.B(n_490),
.C(n_449),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_534),
.Y(n_597)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_519),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_583),
.Y(n_593)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_518),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_452),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_584),
.B(n_549),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_528),
.A2(n_517),
.B1(n_438),
.B2(n_471),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_585),
.A2(n_539),
.B1(n_540),
.B2(n_528),
.Y(n_587)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_519),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_586),
.B(n_527),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_587),
.A2(n_595),
.B1(n_603),
.B2(n_559),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_588),
.B(n_571),
.Y(n_630)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_591),
.B(n_598),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_600),
.Y(n_620)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_594),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_568),
.A2(n_547),
.B1(n_524),
.B2(n_552),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_597),
.A2(n_569),
.B(n_561),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_578),
.B(n_573),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_560),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_599),
.B(n_608),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_544),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_601),
.B(n_606),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_565),
.B(n_547),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_SL g622 ( 
.A(n_602),
.B(n_604),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_576),
.A2(n_524),
.B1(n_553),
.B2(n_527),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_SL g604 ( 
.A(n_574),
.B(n_563),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_579),
.A2(n_542),
.B(n_535),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_605),
.A2(n_579),
.B(n_581),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_531),
.C(n_535),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_531),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_610),
.B(n_561),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_586),
.B(n_438),
.C(n_456),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_611),
.B(n_471),
.Y(n_629)
);

AOI21x1_ASAP7_75t_SL g648 ( 
.A1(n_614),
.A2(n_632),
.B(n_628),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_607),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_615),
.B(n_617),
.Y(n_645)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_616),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_596),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_608),
.B(n_566),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_619),
.B(n_606),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_592),
.Y(n_641)
);

BUFx12f_ASAP7_75t_SL g623 ( 
.A(n_588),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_623),
.A2(n_593),
.B(n_604),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_612),
.A2(n_567),
.B1(n_570),
.B2(n_580),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_625),
.A2(n_432),
.B1(n_632),
.B2(n_616),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_609),
.B(n_582),
.Y(n_627)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_627),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_605),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_629),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_630),
.B(n_633),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_597),
.A2(n_556),
.B(n_575),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_626),
.B(n_557),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_634),
.B(n_649),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_630),
.B(n_598),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_635),
.B(n_637),
.Y(n_652)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_638),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_626),
.B(n_591),
.C(n_601),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_SL g656 ( 
.A(n_640),
.B(n_624),
.Y(n_656)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_641),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_627),
.B(n_610),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_642),
.B(n_651),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_618),
.A2(n_595),
.B(n_589),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_643),
.B(n_650),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_621),
.A2(n_603),
.B1(n_564),
.B2(n_585),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_644),
.A2(n_613),
.B1(n_622),
.B2(n_641),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_648),
.A2(n_614),
.B(n_620),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_631),
.B(n_611),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_623),
.A2(n_602),
.B(n_433),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_635),
.B(n_640),
.C(n_624),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_654),
.B(n_656),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_647),
.B(n_633),
.C(n_620),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_661),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_639),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_662),
.B(n_664),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_636),
.B(n_625),
.C(n_622),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_663),
.B(n_646),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_655),
.B(n_645),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_666),
.B(n_671),
.Y(n_676)
);

AOI21xp33_ASAP7_75t_L g678 ( 
.A1(n_667),
.A2(n_657),
.B(n_659),
.Y(n_678)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_654),
.B(n_662),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_669),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_639),
.Y(n_669)
);

OAI21x1_ASAP7_75t_SL g670 ( 
.A1(n_653),
.A2(n_648),
.B(n_641),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_670),
.A2(n_661),
.B(n_663),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_652),
.B(n_660),
.Y(n_671)
);

OAI211xp5_ASAP7_75t_L g679 ( 
.A1(n_675),
.A2(n_678),
.B(n_676),
.C(n_665),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_R g677 ( 
.A(n_672),
.B(n_652),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_677),
.A2(n_673),
.B(n_671),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_679),
.A2(n_680),
.B(n_673),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_674),
.B(n_669),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_681),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_683),
.B(n_660),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_682),
.C(n_644),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_685),
.A2(n_642),
.B(n_684),
.Y(n_686)
);

BUFx24_ASAP7_75t_SL g687 ( 
.A(n_686),
.Y(n_687)
);


endmodule