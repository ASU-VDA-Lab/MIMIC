module fake_jpeg_20362_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_27),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_73),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_57),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_63),
.B1(n_46),
.B2(n_54),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_80),
.B1(n_60),
.B2(n_65),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_55),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_66),
.B(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_61),
.B1(n_65),
.B2(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_57),
.B1(n_60),
.B2(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_52),
.B1(n_59),
.B2(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_91),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_49),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_58),
.B(n_1),
.C(n_2),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_50),
.C(n_29),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_0),
.C(n_1),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_108),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_20),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_15),
.B(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_116),
.B1(n_103),
.B2(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_14),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_23),
.Y(n_119)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_121),
.C(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_114),
.C(n_33),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_123),
.C(n_114),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_30),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_120),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_34),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_35),
.B(n_38),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_42),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_107),
.Y(n_133)
);


endmodule