module real_jpeg_49_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_2),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_102),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_2),
.A2(n_39),
.B1(n_45),
.B2(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_34),
.B(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_98),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_51),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_3),
.A2(n_26),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_39),
.C(n_88),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_3),
.B(n_42),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_92),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_39),
.B1(n_45),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_4),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_6),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_6),
.A2(n_44),
.B1(n_52),
.B2(n_53),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_8),
.A2(n_39),
.B1(n_45),
.B2(n_59),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_63),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_9),
.A2(n_39),
.B1(n_45),
.B2(n_63),
.Y(n_157)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_12),
.A2(n_39),
.B1(n_45),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_13),
.A2(n_32),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_13),
.A2(n_39),
.B1(n_45),
.B2(n_70),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_15),
.A2(n_39),
.B1(n_45),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_16),
.A2(n_32),
.B1(n_35),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_73),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_16),
.A2(n_39),
.B1(n_45),
.B2(n_73),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_109),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_109),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_74),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_49),
.C(n_64),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_24),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_25),
.B(n_37),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.A3(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_26),
.A2(n_53),
.A3(n_55),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_27),
.B(n_153),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_38),
.A2(n_42),
.B1(n_78),
.B2(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_38),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_38),
.A2(n_42),
.B1(n_157),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_38),
.A2(n_42),
.B1(n_153),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_38),
.A2(n_42),
.B1(n_196),
.B2(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_45),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_39),
.B(n_194),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_41),
.A2(n_47),
.B1(n_79),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_41),
.A2(n_108),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_41),
.A2(n_108),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_64),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_49)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_50),
.A2(n_58),
.B1(n_60),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_50),
.A2(n_60),
.B1(n_119),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_50),
.A2(n_60),
.B1(n_133),
.B2(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_62),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AO22x2_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_53),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_52),
.B(n_56),
.Y(n_154)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_53),
.B(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_72),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_94),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_93),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_90),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_92),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_92),
.B1(n_116),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_86),
.A2(n_92),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_86),
.A2(n_92),
.B1(n_166),
.B2(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_90),
.A2(n_106),
.B1(n_149),
.B2(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_107),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_120),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_141),
.B(n_216),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_139),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_126),
.B(n_139),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_131),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_131),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_161),
.B(n_215),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_159),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_159),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_150),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_150),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_210),
.B(n_214),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_179),
.B(n_209),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_171),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_168),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_174),
.C(n_177),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_190),
.B(n_208),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_202),
.B(n_207),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B(n_201),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_206),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_213),
.Y(n_214)
);


endmodule