module fake_jpeg_27526_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_18),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_31),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_57),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_17),
.B(n_29),
.C(n_27),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_42),
.C(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_20),
.B1(n_30),
.B2(n_16),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_39),
.B1(n_38),
.B2(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_70),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_36),
.C(n_42),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_30),
.B1(n_16),
.B2(n_23),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_34),
.B1(n_41),
.B2(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_30),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_56),
.B1(n_54),
.B2(n_44),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_22),
.B1(n_33),
.B2(n_19),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_100)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_51),
.B(n_53),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_108),
.B(n_75),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_98),
.B1(n_104),
.B2(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_32),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_54),
.B1(n_34),
.B2(n_41),
.Y(n_104)
);

OAI22x1_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_36),
.B1(n_42),
.B2(n_40),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_111),
.B1(n_114),
.B2(n_72),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_21),
.B(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_24),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_54),
.B1(n_56),
.B2(n_52),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_68),
.C(n_85),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_56),
.B1(n_50),
.B2(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_56),
.B1(n_21),
.B2(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_75),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_127),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_58),
.C(n_77),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_69),
.B(n_87),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_135),
.B(n_144),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_133),
.B(n_95),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_65),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_24),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_125),
.A2(n_109),
.B1(n_80),
.B2(n_78),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_62),
.B1(n_90),
.B2(n_67),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_132),
.B1(n_143),
.B2(n_93),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_64),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_86),
.B1(n_74),
.B2(n_71),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_108),
.B(n_110),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_100),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_93),
.B1(n_103),
.B2(n_92),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_102),
.B(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_92),
.B(n_28),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_89),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_147),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_28),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_77),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_138),
.B(n_123),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_152),
.B(n_164),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_106),
.B(n_109),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_157),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_28),
.B1(n_9),
.B2(n_10),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_31),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_171),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_178),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_66),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_95),
.B(n_1),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_172),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_174),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_32),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_153),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_128),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_144),
.B1(n_147),
.B2(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_119),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_182),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_125),
.B1(n_126),
.B2(n_135),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_126),
.B1(n_143),
.B2(n_121),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_190),
.B1(n_194),
.B2(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_193),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_174),
.B1(n_161),
.B2(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

XOR2x1_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_120),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_5),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_141),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_140),
.B1(n_77),
.B2(n_32),
.Y(n_201)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_155),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_32),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_0),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_149),
.B(n_28),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_169),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_172),
.B1(n_149),
.B2(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_5),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_161),
.B1(n_158),
.B2(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_213),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_227),
.B1(n_228),
.B2(n_209),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_163),
.B(n_156),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_221),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_159),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_175),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_154),
.B1(n_163),
.B2(n_171),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_235),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_236),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_188),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_5),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_224),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_192),
.C(n_200),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_245),
.C(n_247),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_187),
.C(n_203),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_220),
.C(n_227),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_215),
.B1(n_232),
.B2(n_201),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_189),
.C(n_196),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_257),
.C(n_199),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_232),
.B1(n_228),
.B2(n_193),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_256),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_189),
.C(n_207),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_237),
.B(n_207),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_273),
.B(n_10),
.Y(n_285)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_265),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_254),
.B(n_257),
.C(n_216),
.D(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_238),
.B(n_237),
.CI(n_235),
.CON(n_267),
.SN(n_267)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_274),
.Y(n_275)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_199),
.C(n_208),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_271),
.C(n_249),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_201),
.C(n_7),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_7),
.B(n_11),
.Y(n_273)
);

OAI322xp33_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_241),
.A3(n_244),
.B1(n_249),
.B2(n_240),
.C1(n_243),
.C2(n_245),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_259),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_282),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_268),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_261),
.B1(n_258),
.B2(n_271),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_287),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_4),
.B(n_2),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_11),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_259),
.C(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_3),
.C(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_264),
.B1(n_270),
.B2(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_300),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_267),
.B1(n_15),
.B2(n_4),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_299),
.B1(n_285),
.B2(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_15),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_306),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_275),
.B1(n_288),
.B2(n_2),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_307),
.C(n_304),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_295),
.B(n_299),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_305),
.B(n_294),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_311),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_291),
.B(n_3),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_310),
.B(n_315),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_314),
.B1(n_308),
.B2(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_301),
.C(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_309),
.Y(n_323)
);


endmodule