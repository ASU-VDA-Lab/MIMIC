module real_aes_7848_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g432 ( .A(n_0), .Y(n_432) );
INVx1_ASAP7_75t_L g471 ( .A(n_1), .Y(n_471) );
INVx1_ASAP7_75t_L g181 ( .A(n_2), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_3), .A2(n_35), .B1(n_137), .B2(n_487), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g161 ( .A1(n_4), .A2(n_118), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_5), .B(n_111), .Y(n_462) );
AND2x6_ASAP7_75t_L g123 ( .A(n_6), .B(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_7), .A2(n_220), .B(n_221), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_8), .B(n_36), .Y(n_433) );
INVx1_ASAP7_75t_L g168 ( .A(n_9), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_10), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g116 ( .A(n_11), .Y(n_116) );
INVx1_ASAP7_75t_L g466 ( .A(n_12), .Y(n_466) );
INVx1_ASAP7_75t_L g226 ( .A(n_13), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_14), .B(n_149), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_15), .B(n_112), .Y(n_443) );
AO32x2_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_111), .A3(n_146), .B1(n_449), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_17), .B(n_137), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_18), .B(n_132), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_19), .B(n_112), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_20), .A2(n_49), .B1(n_137), .B2(n_487), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_21), .B(n_118), .Y(n_192) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_22), .A2(n_73), .B1(n_137), .B2(n_149), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_23), .B(n_137), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_24), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_25), .A2(n_224), .B(n_225), .C(n_227), .Y(n_223) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_26), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_27), .B(n_170), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_28), .B(n_166), .Y(n_183) );
INVx1_ASAP7_75t_L g155 ( .A(n_29), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_30), .B(n_170), .Y(n_510) );
INVx2_ASAP7_75t_L g121 ( .A(n_31), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_32), .B(n_137), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_33), .B(n_170), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_34), .A2(n_123), .B(n_127), .C(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g153 ( .A(n_37), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_38), .B(n_166), .Y(n_236) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_39), .A2(n_42), .B1(n_101), .B2(n_713), .C1(n_718), .C2(n_719), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g718 ( .A(n_39), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_40), .B(n_137), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_41), .A2(n_84), .B1(n_199), .B2(n_487), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_43), .B(n_137), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_44), .B(n_137), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_45), .Y(n_738) );
CKINVDCx16_ASAP7_75t_R g156 ( .A(n_46), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_47), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_48), .B(n_118), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_50), .A2(n_59), .B1(n_137), .B2(n_149), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_51), .A2(n_127), .B1(n_149), .B2(n_151), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_52), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_53), .B(n_137), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_54), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_55), .B(n_137), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_56), .A2(n_136), .B(n_165), .C(n_167), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_57), .Y(n_240) );
INVx1_ASAP7_75t_L g163 ( .A(n_58), .Y(n_163) );
INVx1_ASAP7_75t_L g124 ( .A(n_60), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_61), .B(n_137), .Y(n_472) );
INVx1_ASAP7_75t_L g115 ( .A(n_62), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_63), .Y(n_726) );
AO32x2_ASAP7_75t_L g490 ( .A1(n_64), .A2(n_111), .A3(n_206), .B1(n_449), .B2(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g529 ( .A(n_65), .Y(n_529) );
INVx1_ASAP7_75t_L g505 ( .A(n_66), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_SL g131 ( .A1(n_67), .A2(n_132), .B(n_133), .C(n_136), .Y(n_131) );
INVxp67_ASAP7_75t_L g134 ( .A(n_68), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_69), .B(n_149), .Y(n_506) );
INVx1_ASAP7_75t_L g725 ( .A(n_70), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_71), .Y(n_159) );
INVx1_ASAP7_75t_L g233 ( .A(n_72), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_74), .A2(n_123), .B(n_127), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_75), .B(n_487), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_76), .A2(n_99), .B1(n_721), .B2(n_730), .C1(n_741), .C2(n_747), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_76), .A2(n_102), .B1(n_103), .B2(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_76), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_77), .B(n_149), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_78), .B(n_182), .Y(n_195) );
INVx2_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_80), .B(n_132), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_81), .B(n_149), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_82), .A2(n_123), .B(n_127), .C(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g430 ( .A(n_83), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g435 ( .A(n_83), .Y(n_435) );
OR2x2_ASAP7_75t_L g729 ( .A(n_83), .B(n_720), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_85), .A2(n_97), .B1(n_149), .B2(n_150), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_86), .B(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_87), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_88), .A2(n_123), .B(n_127), .C(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_89), .Y(n_216) );
INVx1_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g222 ( .A(n_91), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_92), .B(n_182), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_93), .B(n_149), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_94), .B(n_111), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_95), .A2(n_118), .B(n_125), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_96), .B(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22x1_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_428), .B1(n_434), .B2(n_436), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_103), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_713) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_365), .Y(n_103) );
NOR4xp25_ASAP7_75t_L g104 ( .A(n_105), .B(n_295), .C(n_326), .D(n_345), .Y(n_104) );
NAND4xp25_ASAP7_75t_L g105 ( .A(n_106), .B(n_253), .C(n_268), .D(n_286), .Y(n_105) );
AOI222xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_188), .B1(n_229), .B2(n_241), .C1(n_246), .C2(n_248), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_171), .Y(n_107) );
INVx1_ASAP7_75t_L g309 ( .A(n_108), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_142), .Y(n_108) );
AND2x2_ASAP7_75t_L g172 ( .A(n_109), .B(n_160), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_109), .B(n_175), .Y(n_338) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g245 ( .A(n_110), .B(n_144), .Y(n_245) );
AND2x2_ASAP7_75t_L g254 ( .A(n_110), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g280 ( .A(n_110), .Y(n_280) );
AND2x2_ASAP7_75t_L g301 ( .A(n_110), .B(n_144), .Y(n_301) );
BUFx2_ASAP7_75t_L g324 ( .A(n_110), .Y(n_324) );
AND2x2_ASAP7_75t_L g348 ( .A(n_110), .B(n_145), .Y(n_348) );
AND2x2_ASAP7_75t_L g412 ( .A(n_110), .B(n_160), .Y(n_412) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_117), .B(n_139), .Y(n_110) );
INVx4_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_111), .A2(n_454), .B(n_462), .Y(n_453) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g146 ( .A(n_112), .Y(n_146) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_113), .B(n_114), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
BUFx2_ASAP7_75t_L g220 ( .A(n_118), .Y(n_220) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
NAND2x1p5_ASAP7_75t_L g157 ( .A(n_119), .B(n_123), .Y(n_157) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g461 ( .A(n_120), .Y(n_461) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g128 ( .A(n_121), .Y(n_128) );
INVx1_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
INVx1_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
INVx1_ASAP7_75t_L g132 ( .A(n_122), .Y(n_132) );
INVx3_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx4_ASAP7_75t_SL g138 ( .A(n_123), .Y(n_138) );
BUFx3_ASAP7_75t_L g449 ( .A(n_123), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_123), .A2(n_455), .B(n_458), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_123), .A2(n_465), .B(n_469), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_123), .A2(n_480), .B(n_484), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_123), .A2(n_504), .B(n_507), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_130), .B(n_131), .C(n_138), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_126), .A2(n_138), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_126), .A2(n_138), .B(n_222), .C(n_223), .Y(n_221) );
INVx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_128), .Y(n_137) );
BUFx3_ASAP7_75t_L g199 ( .A(n_128), .Y(n_199) );
INVx1_ASAP7_75t_L g487 ( .A(n_128), .Y(n_487) );
INVx1_ASAP7_75t_L g483 ( .A(n_132), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_135), .B(n_168), .Y(n_167) );
INVx5_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_135), .A2(n_166), .B1(n_492), .B2(n_493), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_SL g504 ( .A1(n_136), .A2(n_182), .B(n_505), .C(n_506), .Y(n_504) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g147 ( .A1(n_138), .A2(n_148), .B1(n_156), .B2(n_157), .Y(n_147) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_140), .A2(n_161), .B(n_169), .Y(n_160) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_SL g201 ( .A(n_141), .B(n_202), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_141), .B(n_445), .C(n_449), .Y(n_444) );
AO21x1_ASAP7_75t_L g537 ( .A1(n_141), .A2(n_445), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g313 ( .A(n_142), .B(n_244), .Y(n_313) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_143), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_160), .Y(n_143) );
OR2x2_ASAP7_75t_L g273 ( .A(n_144), .B(n_176), .Y(n_273) );
AND2x2_ASAP7_75t_L g285 ( .A(n_144), .B(n_244), .Y(n_285) );
BUFx2_ASAP7_75t_L g417 ( .A(n_144), .Y(n_417) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g174 ( .A(n_145), .B(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g267 ( .A(n_145), .B(n_176), .Y(n_267) );
AND2x2_ASAP7_75t_L g320 ( .A(n_145), .B(n_160), .Y(n_320) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_145), .Y(n_356) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_158), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_146), .B(n_159), .Y(n_158) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_146), .A2(n_177), .B(n_185), .Y(n_176) );
INVx2_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
INVx2_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_151) );
INVx2_ASAP7_75t_L g154 ( .A(n_152), .Y(n_154) );
INVx4_ASAP7_75t_L g224 ( .A(n_152), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_157), .A2(n_178), .B(n_179), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_233), .B(n_234), .Y(n_232) );
AND2x2_ASAP7_75t_L g243 ( .A(n_160), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_SL g255 ( .A(n_160), .Y(n_255) );
INVx2_ASAP7_75t_L g266 ( .A(n_160), .Y(n_266) );
BUFx2_ASAP7_75t_L g290 ( .A(n_160), .Y(n_290) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_160), .B(n_348), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_165), .A2(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_L g528 ( .A1(n_165), .A2(n_470), .B(n_529), .C(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_166), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_166), .A2(n_447), .B1(n_497), .B2(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
INVx2_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_170), .A2(n_219), .B(n_228), .Y(n_218) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_170), .A2(n_479), .B(n_488), .Y(n_478) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_170), .A2(n_503), .B(n_510), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
AOI332xp33_ASAP7_75t_L g268 ( .A1(n_172), .A2(n_269), .A3(n_273), .B1(n_274), .B2(n_278), .B3(n_281), .C1(n_282), .C2(n_284), .Y(n_268) );
NAND2x1_ASAP7_75t_L g353 ( .A(n_172), .B(n_244), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_172), .B(n_258), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_SL g286 ( .A1(n_173), .A2(n_287), .B(n_290), .C(n_291), .Y(n_286) );
AND2x2_ASAP7_75t_L g425 ( .A(n_173), .B(n_266), .Y(n_425) );
INVx3_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
OR2x2_ASAP7_75t_L g322 ( .A(n_174), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g327 ( .A(n_174), .B(n_324), .Y(n_327) );
INVx1_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
AND2x2_ASAP7_75t_L g361 ( .A(n_175), .B(n_320), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_175), .B(n_301), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_175), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_175), .B(n_279), .Y(n_387) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g244 ( .A(n_176), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .C(n_184), .Y(n_180) );
INVx2_ASAP7_75t_L g447 ( .A(n_182), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_182), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_182), .A2(n_526), .B(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_184), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_187), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_187), .B(n_240), .Y(n_239) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_188), .A2(n_347), .A3(n_354), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_203), .Y(n_188) );
AND2x2_ASAP7_75t_L g229 ( .A(n_189), .B(n_230), .Y(n_229) );
NAND2x1_ASAP7_75t_SL g249 ( .A(n_189), .B(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_189), .Y(n_336) );
AND2x2_ASAP7_75t_L g341 ( .A(n_189), .B(n_252), .Y(n_341) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_190), .A2(n_254), .B(n_256), .C(n_259), .Y(n_253) );
OR2x2_ASAP7_75t_L g270 ( .A(n_190), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g283 ( .A(n_190), .Y(n_283) );
AND2x2_ASAP7_75t_L g289 ( .A(n_190), .B(n_231), .Y(n_289) );
INVx2_ASAP7_75t_L g307 ( .A(n_190), .Y(n_307) );
AND2x2_ASAP7_75t_L g318 ( .A(n_190), .B(n_272), .Y(n_318) );
AND2x2_ASAP7_75t_L g350 ( .A(n_190), .B(n_308), .Y(n_350) );
AND2x2_ASAP7_75t_L g354 ( .A(n_190), .B(n_277), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_190), .B(n_203), .Y(n_359) );
AND2x2_ASAP7_75t_L g393 ( .A(n_190), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_190), .B(n_296), .Y(n_427) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
AOI21xp5_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_193), .B(n_200), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
INVx1_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_200), .A2(n_464), .B(n_473), .Y(n_463) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_200), .A2(n_524), .B(n_531), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_203), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g335 ( .A(n_203), .Y(n_335) );
AND2x2_ASAP7_75t_L g397 ( .A(n_203), .B(n_318), .Y(n_397) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_217), .Y(n_203) );
OR2x2_ASAP7_75t_L g251 ( .A(n_204), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g261 ( .A(n_204), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_204), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g369 ( .A(n_204), .Y(n_369) );
AND2x2_ASAP7_75t_L g386 ( .A(n_204), .B(n_231), .Y(n_386) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g277 ( .A(n_205), .B(n_217), .Y(n_277) );
AND2x2_ASAP7_75t_L g306 ( .A(n_205), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g317 ( .A(n_205), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_205), .B(n_272), .Y(n_408) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_215), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_214), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g230 ( .A(n_218), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
AND2x2_ASAP7_75t_L g308 ( .A(n_218), .B(n_272), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_224), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g468 ( .A(n_224), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_224), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g410 ( .A(n_229), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_230), .Y(n_414) );
INVx2_ASAP7_75t_L g272 ( .A(n_231), .Y(n_272) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_238), .B(n_239), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_245), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_243), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_243), .B(n_348), .Y(n_406) );
OR2x2_ASAP7_75t_L g247 ( .A(n_244), .B(n_245), .Y(n_247) );
INVx1_ASAP7_75t_SL g299 ( .A(n_244), .Y(n_299) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_250), .A2(n_303), .B1(n_305), .B2(n_309), .C(n_310), .Y(n_302) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g330 ( .A(n_251), .B(n_294), .Y(n_330) );
INVx2_ASAP7_75t_L g262 ( .A(n_252), .Y(n_262) );
INVx1_ASAP7_75t_L g288 ( .A(n_252), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_252), .B(n_272), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_252), .B(n_275), .Y(n_382) );
INVx1_ASAP7_75t_L g390 ( .A(n_252), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_254), .B(n_258), .Y(n_304) );
AND2x4_ASAP7_75t_L g279 ( .A(n_255), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g392 ( .A(n_258), .B(n_348), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_261), .B(n_293), .Y(n_292) );
INVxp67_ASAP7_75t_L g400 ( .A(n_262), .Y(n_400) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g300 ( .A(n_266), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g372 ( .A(n_266), .B(n_348), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_266), .B(n_285), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g332 ( .A1(n_267), .A2(n_301), .A3(n_308), .B1(n_333), .B2(n_336), .C1(n_337), .C2(n_339), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_267), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g398 ( .A(n_270), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g344 ( .A(n_271), .Y(n_344) );
INVx2_ASAP7_75t_L g275 ( .A(n_272), .Y(n_275) );
INVx1_ASAP7_75t_L g334 ( .A(n_272), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g281 ( .A(n_273), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g370 ( .A(n_275), .B(n_283), .Y(n_370) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g282 ( .A(n_277), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g325 ( .A(n_277), .B(n_318), .Y(n_325) );
AND2x2_ASAP7_75t_L g329 ( .A(n_277), .B(n_289), .Y(n_329) );
OAI21xp33_ASAP7_75t_SL g339 ( .A1(n_278), .A2(n_340), .B(n_342), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_278), .A2(n_410), .B1(n_411), .B2(n_413), .Y(n_409) );
INVx3_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g284 ( .A(n_279), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_279), .B(n_299), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_281), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g421 ( .A(n_288), .Y(n_421) );
INVx4_ASAP7_75t_L g294 ( .A(n_289), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_289), .B(n_316), .Y(n_364) );
INVx1_ASAP7_75t_SL g376 ( .A(n_290), .Y(n_376) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g389 ( .A(n_294), .B(n_390), .Y(n_389) );
OAI211xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_297), .B(n_302), .C(n_319), .Y(n_295) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_297), .A2(n_335), .B1(n_414), .B2(n_416), .C(n_418), .Y(n_415) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_299), .B(n_412), .Y(n_411) );
OAI31xp33_ASAP7_75t_L g391 ( .A1(n_300), .A2(n_377), .A3(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g331 ( .A(n_301), .Y(n_331) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g381 ( .A(n_306), .Y(n_381) );
AND2x2_ASAP7_75t_L g394 ( .A(n_308), .B(n_317), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_314), .Y(n_310) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_318), .B(n_421), .Y(n_420) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B(n_325), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_328), .B1(n_330), .B2(n_331), .C(n_332), .Y(n_326) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_327), .A2(n_396), .B(n_398), .C(n_401), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_330), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g357 ( .A(n_338), .Y(n_357) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g343 ( .A(n_341), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g385 ( .A(n_341), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI211xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B(n_351), .C(n_360), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_349), .A2(n_359), .B1(n_423), .B2(n_424), .C(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B1(n_355), .B2(n_358), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_SL g423 ( .A(n_362), .Y(n_423) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_395), .C(n_415), .D(n_422), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B(n_373), .C(n_391), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B(n_379), .C(n_383), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g402 ( .A(n_380), .Y(n_402) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
OR2x2_ASAP7_75t_L g413 ( .A(n_381), .B(n_414), .Y(n_413) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_412), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g714 ( .A(n_429), .Y(n_714) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g434 ( .A(n_431), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g720 ( .A(n_431), .Y(n_720) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g716 ( .A(n_434), .Y(n_716) );
NOR2x2_ASAP7_75t_L g719 ( .A(n_435), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g717 ( .A(n_436), .Y(n_717) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_438), .B(n_647), .Y(n_437) );
NOR5xp2_ASAP7_75t_L g438 ( .A(n_439), .B(n_560), .C(n_606), .D(n_619), .E(n_631), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_474), .B(n_514), .C(n_541), .Y(n_439) );
INVx1_ASAP7_75t_SL g642 ( .A(n_440), .Y(n_642) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_450), .Y(n_440) );
AND2x2_ASAP7_75t_L g566 ( .A(n_441), .B(n_451), .Y(n_566) );
AND2x2_ASAP7_75t_L g594 ( .A(n_441), .B(n_540), .Y(n_594) );
AND2x2_ASAP7_75t_L g602 ( .A(n_441), .B(n_545), .Y(n_602) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g532 ( .A(n_442), .B(n_452), .Y(n_532) );
INVx2_ASAP7_75t_L g544 ( .A(n_442), .Y(n_544) );
AND2x2_ASAP7_75t_L g669 ( .A(n_442), .B(n_611), .Y(n_669) );
OR2x2_ASAP7_75t_L g671 ( .A(n_442), .B(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g538 ( .A(n_443), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_447), .A2(n_459), .B(n_460), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_447), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_449), .A2(n_525), .B(n_528), .Y(n_524) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g582 ( .A(n_451), .B(n_554), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_451), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g696 ( .A(n_451), .B(n_536), .Y(n_696) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .Y(n_451) );
AND2x2_ASAP7_75t_L g539 ( .A(n_452), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g586 ( .A(n_452), .Y(n_586) );
AND2x2_ASAP7_75t_L g611 ( .A(n_452), .B(n_523), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_452), .B(n_644), .Y(n_681) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g545 ( .A(n_453), .B(n_523), .Y(n_545) );
AND2x2_ASAP7_75t_L g559 ( .A(n_453), .B(n_522), .Y(n_559) );
AND2x2_ASAP7_75t_L g576 ( .A(n_453), .B(n_463), .Y(n_576) );
AND2x2_ASAP7_75t_L g633 ( .A(n_453), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_453), .B(n_540), .Y(n_646) );
AND2x2_ASAP7_75t_L g698 ( .A(n_453), .B(n_623), .Y(n_698) );
INVx2_ASAP7_75t_L g470 ( .A(n_461), .Y(n_470) );
AND2x2_ASAP7_75t_L g521 ( .A(n_463), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g540 ( .A(n_463), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_463), .B(n_523), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_499), .B(n_511), .Y(n_474) );
INVx1_ASAP7_75t_SL g630 ( .A(n_475), .Y(n_630) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_489), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_477), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g513 ( .A(n_478), .Y(n_513) );
INVx1_ASAP7_75t_L g550 ( .A(n_478), .Y(n_550) );
AND2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_494), .Y(n_571) );
AND2x2_ASAP7_75t_L g605 ( .A(n_478), .B(n_495), .Y(n_605) );
OR2x2_ASAP7_75t_L g624 ( .A(n_478), .B(n_501), .Y(n_624) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_478), .Y(n_638) );
AND2x2_ASAP7_75t_L g651 ( .A(n_478), .B(n_652), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_483), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_489), .A2(n_573), .B1(n_574), .B2(n_583), .Y(n_572) );
AND2x2_ASAP7_75t_L g656 ( .A(n_489), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
INVx1_ASAP7_75t_L g517 ( .A(n_490), .Y(n_517) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
INVx1_ASAP7_75t_L g565 ( .A(n_490), .Y(n_565) );
AND2x2_ASAP7_75t_L g580 ( .A(n_490), .B(n_495), .Y(n_580) );
OR2x2_ASAP7_75t_L g534 ( .A(n_494), .B(n_519), .Y(n_534) );
AND2x2_ASAP7_75t_L g564 ( .A(n_494), .B(n_565), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g652 ( .A(n_494), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g512 ( .A(n_495), .B(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g621 ( .A(n_495), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_499), .B(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g599 ( .A(n_500), .B(n_565), .Y(n_599) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g511 ( .A(n_501), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g570 ( .A(n_501), .Y(n_570) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g519 ( .A(n_502), .Y(n_519) );
OR2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_502), .Y(n_604) );
AOI32xp33_ASAP7_75t_L g641 ( .A1(n_511), .A2(n_571), .A3(n_642), .B1(n_643), .B2(n_645), .Y(n_641) );
AND2x2_ASAP7_75t_L g567 ( .A(n_512), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_512), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_512), .B(n_599), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_512), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_520), .B1(n_533), .B2(n_535), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
AND2x2_ASAP7_75t_L g620 ( .A(n_516), .B(n_621), .Y(n_620) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_517), .B(n_519), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_518), .A2(n_542), .B1(n_546), .B2(n_556), .Y(n_541) );
AND2x2_ASAP7_75t_L g563 ( .A(n_518), .B(n_564), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_518), .A2(n_532), .B(n_580), .C(n_615), .Y(n_614) );
OAI332xp33_ASAP7_75t_L g619 ( .A1(n_518), .A2(n_620), .A3(n_622), .B1(n_624), .B2(n_625), .B3(n_627), .C1(n_628), .C2(n_630), .Y(n_619) );
INVx2_ASAP7_75t_L g660 ( .A(n_518), .Y(n_660) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_519), .Y(n_578) );
INVx1_ASAP7_75t_L g653 ( .A(n_519), .Y(n_653) );
AND2x2_ASAP7_75t_L g707 ( .A(n_519), .B(n_571), .Y(n_707) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
AND2x2_ASAP7_75t_L g587 ( .A(n_522), .B(n_537), .Y(n_587) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g536 ( .A(n_523), .B(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g635 ( .A(n_523), .B(n_537), .Y(n_635) );
INVx1_ASAP7_75t_L g644 ( .A(n_523), .Y(n_644) );
INVx1_ASAP7_75t_L g618 ( .A(n_532), .Y(n_618) );
INVxp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g702 ( .A(n_534), .B(n_554), .Y(n_702) );
INVx1_ASAP7_75t_SL g613 ( .A(n_535), .Y(n_613) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
AND2x2_ASAP7_75t_L g640 ( .A(n_536), .B(n_598), .Y(n_640) );
INVx1_ASAP7_75t_L g659 ( .A(n_536), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_536), .B(n_626), .Y(n_661) );
INVx1_ASAP7_75t_L g558 ( .A(n_537), .Y(n_558) );
AND2x2_ASAP7_75t_L g562 ( .A(n_539), .B(n_543), .Y(n_562) );
AND2x2_ASAP7_75t_L g629 ( .A(n_539), .B(n_587), .Y(n_629) );
INVx2_ASAP7_75t_L g672 ( .A(n_539), .Y(n_672) );
INVx2_ASAP7_75t_L g555 ( .A(n_540), .Y(n_555) );
AND2x2_ASAP7_75t_L g557 ( .A(n_540), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_544), .B(n_617), .Y(n_623) );
OR2x2_ASAP7_75t_L g687 ( .A(n_544), .B(n_646), .Y(n_687) );
INVx1_ASAP7_75t_L g711 ( .A(n_544), .Y(n_711) );
INVx1_ASAP7_75t_L g667 ( .A(n_545), .Y(n_667) );
AND2x2_ASAP7_75t_L g712 ( .A(n_545), .B(n_555), .Y(n_712) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_549), .A2(n_575), .B1(n_577), .B2(n_581), .Y(n_574) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI322xp33_ASAP7_75t_SL g658 ( .A1(n_552), .A2(n_659), .A3(n_660), .B1(n_661), .B2(n_662), .C1(n_665), .C2(n_667), .Y(n_658) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g655 ( .A(n_553), .B(n_571), .Y(n_655) );
OR2x2_ASAP7_75t_L g689 ( .A(n_553), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g692 ( .A(n_553), .B(n_624), .Y(n_692) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g637 ( .A(n_554), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g693 ( .A(n_554), .B(n_624), .Y(n_693) );
INVx3_ASAP7_75t_L g626 ( .A(n_555), .Y(n_626) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g682 ( .A(n_557), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g561 ( .A1(n_559), .A2(n_562), .B1(n_563), .B2(n_566), .C1(n_567), .C2(n_569), .Y(n_561) );
INVx1_ASAP7_75t_L g592 ( .A(n_559), .Y(n_592) );
NAND3xp33_ASAP7_75t_SL g560 ( .A(n_561), .B(n_572), .C(n_589), .Y(n_560) );
AND2x2_ASAP7_75t_L g677 ( .A(n_564), .B(n_578), .Y(n_677) );
BUFx2_ASAP7_75t_L g568 ( .A(n_565), .Y(n_568) );
INVx1_ASAP7_75t_L g609 ( .A(n_565), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_566), .A2(n_602), .B1(n_655), .B2(n_656), .C(n_658), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_568), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_571), .Y(n_595) );
AND2x2_ASAP7_75t_L g608 ( .A(n_571), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_576), .B(n_587), .Y(n_588) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_578), .A2(n_584), .B(n_588), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_578), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g675 ( .A(n_580), .B(n_657), .Y(n_675) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g598 ( .A(n_586), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_587), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g704 ( .A(n_587), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .B1(n_596), .B2(n_599), .C(n_600), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_591), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g700 ( .A(n_599), .B(n_605), .Y(n_700) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OAI31xp33_ASAP7_75t_SL g668 ( .A1(n_603), .A2(n_642), .A3(n_669), .B(n_670), .Y(n_668) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g657 ( .A(n_604), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_605), .B(n_609), .Y(n_708) );
OAI221xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_610), .B1(n_612), .B2(n_613), .C(n_614), .Y(n_606) );
INVx1_ASAP7_75t_L g612 ( .A(n_608), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_611), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g627 ( .A(n_620), .Y(n_627) );
INVx2_ASAP7_75t_L g663 ( .A(n_621), .Y(n_663) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g649 ( .A(n_626), .B(n_635), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_626), .A2(n_643), .B(n_700), .C(n_701), .Y(n_699) );
OAI221xp5_ASAP7_75t_SL g631 ( .A1(n_627), .A2(n_632), .B1(n_636), .B2(n_639), .C(n_641), .Y(n_631) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_630), .A2(n_695), .B(n_697), .C(n_699), .Y(n_694) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_633), .A2(n_684), .B1(n_686), .B2(n_688), .C(n_691), .Y(n_683) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_673), .C(n_694), .D(n_705), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_654), .C(n_668), .Y(n_648) );
INVx1_ASAP7_75t_SL g703 ( .A(n_655), .Y(n_703) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g666 ( .A(n_664), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_671), .A2(n_680), .B1(n_692), .B2(n_693), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_678), .C(n_683), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI31xp33_ASAP7_75t_L g705 ( .A1(n_676), .A2(n_706), .A3(n_708), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
NOR2xp33_ASAP7_75t_SL g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_SL g746 ( .A(n_724), .Y(n_746) );
INVx1_ASAP7_75t_L g745 ( .A(n_726), .Y(n_745) );
OA21x2_ASAP7_75t_L g748 ( .A1(n_726), .A2(n_746), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_729), .Y(n_736) );
INVx2_ASAP7_75t_L g740 ( .A(n_729), .Y(n_740) );
BUFx2_ASAP7_75t_L g749 ( .A(n_729), .Y(n_749) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B(n_737), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
CKINVDCx6p67_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
endmodule