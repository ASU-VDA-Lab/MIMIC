module fake_jpeg_27453_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_60),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_34),
.B1(n_16),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_40),
.B1(n_42),
.B2(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_16),
.B1(n_34),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_55),
.B1(n_40),
.B2(n_42),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_16),
.B1(n_34),
.B2(n_28),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_29),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_70),
.B1(n_85),
.B2(n_93),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_72),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_28),
.B1(n_21),
.B2(n_31),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_41),
.B(n_36),
.C(n_38),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_83),
.C(n_94),
.Y(n_108)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_21),
.B1(n_44),
.B2(n_27),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_77),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_36),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_42),
.B1(n_40),
.B2(n_44),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_92),
.B1(n_51),
.B2(n_60),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_27),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_40),
.B1(n_44),
.B2(n_35),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_26),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_74),
.B1(n_89),
.B2(n_91),
.Y(n_134)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_105),
.B1(n_100),
.B2(n_110),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_35),
.B1(n_63),
.B2(n_39),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_116),
.B1(n_83),
.B2(n_92),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_39),
.B1(n_26),
.B2(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_118),
.Y(n_138)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_77),
.B1(n_73),
.B2(n_84),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_123),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_29),
.C(n_24),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_71),
.C(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_124),
.A2(n_134),
.B1(n_66),
.B2(n_43),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_65),
.B(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_149),
.B(n_99),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_127),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_139),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_108),
.C(n_114),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_147),
.C(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_85),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_147),
.B1(n_138),
.B2(n_130),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_23),
.B(n_31),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_152),
.B(n_20),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_23),
.C(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_24),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_24),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_146),
.B(n_151),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_81),
.C(n_80),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_32),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_43),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_91),
.B(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_29),
.B(n_32),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_133),
.B(n_149),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_161),
.Y(n_196)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_159),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_165),
.C(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_107),
.C(n_105),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_107),
.B(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_171),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_78),
.B(n_1),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_152),
.B(n_129),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_173),
.B1(n_175),
.B2(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_184),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_117),
.B1(n_115),
.B2(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_144),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_74),
.B1(n_98),
.B2(n_112),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_180),
.B1(n_186),
.B2(n_188),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_18),
.B1(n_17),
.B2(n_33),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_78),
.C(n_37),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_37),
.C(n_20),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_182),
.C(n_0),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_37),
.C(n_20),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_125),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_32),
.B(n_1),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_139),
.A2(n_18),
.B1(n_17),
.B2(n_33),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_145),
.B(n_32),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_153),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_18),
.B1(n_17),
.B2(n_9),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_197),
.B(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_203),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_144),
.Y(n_197)
);

NAND2x1_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_141),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_169),
.B1(n_178),
.B2(n_171),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_207),
.B1(n_215),
.B2(n_188),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_141),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_184),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_144),
.B1(n_140),
.B2(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_168),
.B1(n_186),
.B2(n_157),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_140),
.B1(n_17),
.B2(n_9),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_162),
.B1(n_163),
.B2(n_174),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_172),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_176),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_160),
.C(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_232),
.C(n_236),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_158),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_180),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_233),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_243),
.B1(n_210),
.B2(n_206),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_166),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_182),
.C(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_14),
.C(n_12),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_12),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_241),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_240),
.B(n_215),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_0),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_196),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_234),
.B1(n_191),
.B2(n_207),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_200),
.B(n_189),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_196),
.C(n_199),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_194),
.C(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_259),
.C(n_221),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_194),
.C(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_189),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_192),
.B(n_190),
.C(n_198),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_281),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_232),
.C(n_220),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.C(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_225),
.C(n_224),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_231),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_248),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_273),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_205),
.Y(n_274)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_190),
.C(n_193),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_206),
.B(n_191),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_251),
.B(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_198),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_264),
.B(n_250),
.Y(n_290)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_233),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_245),
.C(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_244),
.C(n_257),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_269),
.C(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_3),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_253),
.C(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_3),
.C(n_4),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_253),
.B(n_2),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_295),
.B(n_0),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_278),
.B1(n_267),
.B2(n_277),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_281),
.C(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_3),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_294),
.C(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_284),
.B(n_283),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_308),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_4),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_314),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_286),
.B(n_285),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_316),
.B(n_317),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_293),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_297),
.C(n_300),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_293),
.C(n_296),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_304),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.C(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_5),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_5),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_323),
.B(n_321),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B1(n_326),
.B2(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_5),
.C(n_6),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_7),
.C(n_8),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_7),
.B(n_8),
.Y(n_331)
);


endmodule