module fake_jpeg_1841_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_50),
.B1(n_61),
.B2(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_74),
.B1(n_71),
.B2(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_81),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_50),
.B1(n_61),
.B2(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_54),
.B(n_46),
.C(n_47),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_51),
.B1(n_55),
.B2(n_49),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_70),
.B1(n_71),
.B2(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_51),
.B1(n_47),
.B2(n_48),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_70),
.B1(n_58),
.B2(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_96),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_71),
.A3(n_62),
.B1(n_59),
.B2(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_99),
.B1(n_76),
.B2(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_101),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_58),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_6),
.Y(n_101)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_75),
.CI(n_9),
.CON(n_107),
.SN(n_107)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_19),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_115),
.B1(n_117),
.B2(n_18),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_75),
.C(n_76),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_83),
.C(n_26),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_93),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_29),
.B1(n_44),
.B2(n_43),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_15),
.B(n_16),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_14),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_132),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_108),
.B(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_127),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_16),
.B(n_17),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_18),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_19),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_35),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_113),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_107),
.B(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_38),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_127),
.Y(n_151)
);

AND2x4_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_33),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_112),
.C(n_106),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_143),
.C(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_117),
.C(n_24),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_45),
.B1(n_25),
.B2(n_28),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_20),
.A3(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_153),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_20),
.B1(n_42),
.B2(n_41),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_121),
.B(n_128),
.C(n_139),
.D(n_138),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_161),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_140),
.C(n_151),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_166),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_143),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_167),
.Y(n_168)
);

AOI321xp33_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_154),
.A3(n_141),
.B1(n_147),
.B2(n_149),
.C(n_152),
.Y(n_167)
);

XOR2x2_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_163),
.B1(n_165),
.B2(n_158),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_172),
.B1(n_168),
.B2(n_169),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_172),
.C(n_153),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_156),
.C(n_130),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_139),
.B(n_123),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_125),
.B(n_132),
.Y(n_177)
);


endmodule