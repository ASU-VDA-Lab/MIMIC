module fake_ariane_2976_n_1803 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1803);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1803;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_82),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_91),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_50),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_38),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_55),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_3),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_58),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_42),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_35),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_77),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_83),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_26),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_72),
.B(n_60),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_107),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_79),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_36),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_13),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_88),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_41),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_92),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_23),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_93),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_56),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_13),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_41),
.Y(n_211)
);

BUFx8_ASAP7_75t_SL g212 ( 
.A(n_3),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_138),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_8),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_50),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_84),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_97),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_29),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_64),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_23),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_52),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g226 ( 
.A(n_26),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_76),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_6),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_49),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_143),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_158),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_135),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_129),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_46),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_75),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_90),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_112),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_140),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_113),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_80),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_28),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_2),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_142),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_111),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_46),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_68),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_85),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_130),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_37),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_43),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_127),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_94),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_1),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_43),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_16),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_105),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_117),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_42),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_15),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_134),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_108),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_44),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_36),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_53),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_24),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_8),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_57),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_58),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_128),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_98),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_17),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_121),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_10),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_144),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_100),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_40),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_150),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_27),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_48),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_47),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_157),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_106),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_74),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_31),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_69),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_30),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_22),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_95),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_116),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_14),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_34),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_37),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_147),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_12),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_24),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_7),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_25),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_176),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_212),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_233),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_232),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_194),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_239),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_249),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_176),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_312),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_176),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_167),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_165),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_205),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_176),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_176),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_240),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_240),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_207),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_216),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_240),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_240),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_226),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_240),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_217),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_209),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_218),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_204),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_208),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_204),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_235),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_166),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_235),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_223),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_261),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_225),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_236),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_261),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_282),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_268),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_288),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_161),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_245),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_211),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_215),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_265),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_265),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_169),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_192),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_300),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_177),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_180),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_198),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_317),
.B(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_335),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_318),
.B(n_193),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_326),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_319),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_319),
.B(n_320),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

AND3x2_ASAP7_75t_L g405 ( 
.A(n_325),
.B(n_227),
.C(n_186),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_342),
.A2(n_170),
.B1(n_161),
.B2(n_310),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_375),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_374),
.B(n_186),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_361),
.B(n_306),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_329),
.B(n_159),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_330),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_360),
.B(n_192),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_170),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_363),
.B(n_192),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_375),
.B(n_306),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_166),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_338),
.A2(n_172),
.B(n_168),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_377),
.B(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_339),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_173),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_322),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_340),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_334),
.A2(n_284),
.B1(n_175),
.B2(n_310),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_340),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_323),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_344),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_384),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_367),
.A2(n_190),
.B1(n_187),
.B2(n_309),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_345),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_345),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_379),
.B(n_183),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_380),
.B(n_191),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_365),
.B(n_287),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_347),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_348),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_348),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_350),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_350),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_404),
.Y(n_463)
);

INVxp33_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_413),
.B(n_343),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_413),
.B(n_351),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_404),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_383),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_414),
.B(n_356),
.Y(n_472)
);

CKINVDCx6p67_ASAP7_75t_R g473 ( 
.A(n_450),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_393),
.B(n_362),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_428),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_408),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_393),
.B(n_364),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_396),
.B(n_366),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_414),
.B(n_160),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

BUFx6f_ASAP7_75t_SL g490 ( 
.A(n_416),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_430),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_422),
.B(n_427),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_422),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_396),
.B(n_353),
.Y(n_495)
);

BUFx4f_ASAP7_75t_L g496 ( 
.A(n_437),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_427),
.B(n_389),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

INVx11_ASAP7_75t_L g499 ( 
.A(n_443),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_406),
.B(n_376),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_392),
.B(n_355),
.C(n_354),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_380),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_406),
.B(n_381),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_394),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_418),
.B(n_160),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_418),
.B(n_162),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_457),
.B(n_441),
.Y(n_514)
);

CKINVDCx6p67_ASAP7_75t_R g515 ( 
.A(n_450),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_445),
.A2(n_224),
.B1(n_270),
.B2(n_256),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_426),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g518 ( 
.A(n_398),
.B(n_399),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_457),
.B(n_162),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_457),
.B(n_381),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_394),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_397),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_397),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_409),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_400),
.B(n_163),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_409),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_411),
.B(n_382),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

AND3x2_ASAP7_75t_L g534 ( 
.A(n_416),
.B(n_263),
.C(n_230),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_445),
.B(n_163),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_420),
.B(n_382),
.Y(n_537)
);

AND3x2_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_292),
.C(n_201),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_412),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_421),
.A2(n_386),
.B(n_385),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_447),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_416),
.A2(n_295),
.B1(n_187),
.B2(n_185),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_L g550 ( 
.A(n_424),
.B(n_164),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_416),
.B(n_164),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_425),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_425),
.B(n_412),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_412),
.B(n_171),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_412),
.B(n_171),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_447),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_461),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_412),
.B(n_435),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_423),
.B(n_391),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_405),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_417),
.B(n_355),
.C(n_354),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_417),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_431),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_431),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_442),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_436),
.B(n_385),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_403),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_407),
.B(n_389),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_407),
.A2(n_295),
.B1(n_185),
.B2(n_182),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_435),
.B(n_178),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

INVxp33_ASAP7_75t_SL g585 ( 
.A(n_448),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_395),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_433),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_436),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_433),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_434),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_434),
.Y(n_591)
);

INVxp33_ASAP7_75t_SL g592 ( 
.A(n_423),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_437),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_451),
.A2(n_327),
.B1(n_369),
.B2(n_372),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_434),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_444),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_451),
.B(n_390),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_444),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_447),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_395),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_439),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_436),
.B(n_386),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_455),
.B(n_182),
.C(n_175),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_447),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_439),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_447),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_436),
.B(n_387),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_447),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_453),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_453),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_435),
.B(n_178),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_436),
.A2(n_315),
.B1(n_302),
.B2(n_388),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_453),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_523),
.B(n_571),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_540),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_485),
.B(n_435),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_494),
.B(n_435),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_518),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_571),
.B(n_405),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_471),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_495),
.B(n_455),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_523),
.B(n_179),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_467),
.A2(n_437),
.B1(n_387),
.B2(n_388),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_540),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_501),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_493),
.A2(n_237),
.B1(n_280),
.B2(n_296),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_523),
.B(n_179),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_493),
.A2(n_237),
.B1(n_280),
.B2(n_296),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_523),
.B(n_184),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_501),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_494),
.B(n_497),
.Y(n_632)
);

NAND2x1p5_ASAP7_75t_L g633 ( 
.A(n_588),
.B(n_541),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_510),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_467),
.B(n_184),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_514),
.B(n_456),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_510),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_521),
.B(n_456),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_468),
.B(n_463),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_601),
.B(n_605),
.Y(n_640)
);

BUFx8_ASAP7_75t_L g641 ( 
.A(n_586),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_601),
.B(n_196),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_605),
.B(n_243),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_481),
.B(n_378),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_540),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_588),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_468),
.B(n_188),
.Y(n_647)
);

A2O1A1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_465),
.A2(n_242),
.B(n_246),
.C(n_197),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_463),
.B(n_188),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_471),
.B(n_500),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_475),
.B(n_189),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_482),
.B(n_189),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_497),
.B(n_390),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_588),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_585),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_478),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_469),
.B(n_260),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_229),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_490),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_507),
.B(n_304),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_463),
.B(n_304),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_557),
.B(n_560),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_536),
.B(n_241),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_506),
.B(n_311),
.Y(n_665)
);

O2A1O1Ixp5_ASAP7_75t_L g666 ( 
.A1(n_554),
.A2(n_214),
.B(n_271),
.C(n_258),
.Y(n_666)
);

NOR3xp33_ASAP7_75t_L g667 ( 
.A(n_581),
.B(n_279),
.C(n_190),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_541),
.B(n_311),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_490),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_669)
);

NAND2x1p5_ASAP7_75t_L g670 ( 
.A(n_564),
.B(n_437),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_466),
.B(n_206),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_527),
.A2(n_391),
.B(n_371),
.C(n_370),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_551),
.B(n_486),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_483),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_510),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_516),
.A2(n_285),
.B1(n_279),
.B2(n_284),
.C(n_290),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_499),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_586),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_567),
.B(n_285),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_580),
.A2(n_287),
.B1(n_174),
.B2(n_276),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_478),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_492),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_578),
.B(n_247),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_466),
.B(n_248),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_602),
.B(n_251),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_568),
.B(n_357),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_567),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_607),
.B(n_255),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_580),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_479),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_472),
.B(n_568),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_580),
.B(n_321),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_479),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_491),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_466),
.B(n_252),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_490),
.A2(n_281),
.B1(n_283),
.B2(n_254),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_511),
.B(n_259),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_470),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_513),
.B(n_262),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_583),
.B(n_264),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_531),
.B(n_269),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_537),
.B(n_273),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_603),
.B(n_309),
.C(n_291),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_470),
.B(n_274),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_522),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_522),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_470),
.A2(n_297),
.B(n_303),
.C(n_305),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_522),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_474),
.B(n_275),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_611),
.B(n_277),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_491),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_524),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_552),
.A2(n_402),
.B(n_415),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_524),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_474),
.B(n_476),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_499),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_524),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_474),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_526),
.A2(n_368),
.B(n_359),
.C(n_371),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_526),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_476),
.B(n_290),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_526),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_476),
.B(n_291),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_530),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_473),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_480),
.B(n_484),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_490),
.B(n_294),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_480),
.B(n_294),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_530),
.A2(n_402),
.B(n_415),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_528),
.A2(n_293),
.B1(n_199),
.B2(n_213),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_480),
.B(n_299),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_530),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_550),
.A2(n_195),
.B1(n_219),
.B2(n_220),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_533),
.A2(n_402),
.B(n_415),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_484),
.B(n_487),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_498),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_484),
.B(n_299),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_473),
.B(n_301),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_487),
.B(n_301),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_515),
.B(n_287),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_487),
.B(n_307),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_488),
.B(n_307),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_580),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_488),
.B(n_308),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_534),
.B(n_357),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_488),
.B(n_308),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_489),
.B(n_174),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_489),
.B(n_222),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_515),
.B(n_359),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_489),
.B(n_558),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_533),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_533),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_498),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_549),
.B(n_370),
.C(n_368),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_503),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_561),
.A2(n_462),
.B(n_453),
.C(n_266),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_503),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_547),
.B(n_228),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_508),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_547),
.B(n_231),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_580),
.A2(n_272),
.B1(n_234),
.B2(n_238),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_504),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_504),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_508),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_505),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_547),
.B(n_244),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_572),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_561),
.B(n_174),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_538),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_572),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_558),
.B(n_453),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_572),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_563),
.B(n_276),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_558),
.B(n_565),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_565),
.B(n_253),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_563),
.B(n_276),
.Y(n_777)
);

AO21x2_ASAP7_75t_L g778 ( 
.A1(n_505),
.A2(n_462),
.B(n_453),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_565),
.B(n_257),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_509),
.B(n_267),
.Y(n_780)
);

INVx8_ASAP7_75t_L g781 ( 
.A(n_597),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_509),
.B(n_453),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_597),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_597),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_597),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_SL g786 ( 
.A(n_612),
.B(n_462),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_768),
.Y(n_787)
);

BUFx8_ASAP7_75t_L g788 ( 
.A(n_717),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_645),
.B(n_569),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_645),
.B(n_569),
.Y(n_790)
);

AO22x1_ASAP7_75t_L g791 ( 
.A1(n_658),
.A2(n_592),
.B1(n_464),
.B2(n_594),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_621),
.B(n_597),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_649),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_657),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_658),
.B(n_512),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_768),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_771),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_660),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_675),
.Y(n_799)
);

INVxp33_ASAP7_75t_L g800 ( 
.A(n_644),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_SL g801 ( 
.A(n_678),
.B(n_512),
.C(n_559),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_656),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_682),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_660),
.B(n_566),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_651),
.A2(n_556),
.B1(n_544),
.B2(n_548),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_688),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_771),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_660),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_640),
.A2(n_496),
.B(n_517),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_SL g810 ( 
.A(n_630),
.B(n_553),
.C(n_520),
.Y(n_810)
);

INVx5_ASAP7_75t_L g811 ( 
.A(n_646),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_638),
.B(n_520),
.Y(n_812)
);

BUFx12f_ASAP7_75t_L g813 ( 
.A(n_641),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_656),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_646),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_691),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_694),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_646),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_632),
.B(n_525),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_620),
.B(n_278),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_646),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_632),
.B(n_278),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_636),
.B(n_525),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_616),
.B(n_529),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_641),
.Y(n_825)
);

NOR2x1_ASAP7_75t_L g826 ( 
.A(n_618),
.B(n_570),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_652),
.B(n_529),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_695),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_712),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_726),
.B(n_496),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_750),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_737),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_642),
.B(n_532),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_785),
.A2(n_496),
.B1(n_566),
.B2(n_593),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_639),
.A2(n_496),
.B(n_566),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_643),
.B(n_532),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_645),
.B(n_543),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_674),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_687),
.B(n_535),
.Y(n_839)
);

NAND2x1_ASAP7_75t_L g840 ( 
.A(n_615),
.B(n_543),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_726),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_655),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_687),
.B(n_535),
.Y(n_843)
);

NAND2x2_ASAP7_75t_L g844 ( 
.A(n_680),
.B(n_278),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_654),
.B(n_544),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_664),
.B(n_556),
.C(n_559),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_754),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_681),
.A2(n_593),
.B1(n_566),
.B2(n_545),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_654),
.B(n_545),
.Y(n_849)
);

OAI221xp5_ASAP7_75t_L g850 ( 
.A1(n_681),
.A2(n_555),
.B1(n_548),
.B2(n_553),
.C(n_570),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_617),
.B(n_555),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_683),
.B(n_502),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_679),
.B(n_575),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_781),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_664),
.A2(n_593),
.B1(n_610),
.B2(n_606),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_617),
.B(n_575),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_690),
.B(n_577),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_615),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_781),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_653),
.B(n_619),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_773),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_647),
.B(n_577),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_739),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_781),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_744),
.B(n_508),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_661),
.B(n_582),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_783),
.A2(n_593),
.B1(n_606),
.B2(n_610),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_756),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_655),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_667),
.B(n_502),
.C(n_542),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_645),
.B(n_543),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_623),
.A2(n_584),
.B1(n_582),
.B2(n_596),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_773),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_665),
.B(n_584),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_760),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_746),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_R g877 ( 
.A(n_741),
.B(n_542),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_702),
.B(n_596),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_698),
.B(n_613),
.C(n_609),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_623),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_699),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_626),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_758),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_625),
.A2(n_539),
.B1(n_517),
.B2(n_508),
.Y(n_884)
);

BUFx4f_ASAP7_75t_L g885 ( 
.A(n_633),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_703),
.B(n_596),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_748),
.B(n_598),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_645),
.B(n_543),
.Y(n_888)
);

AND2x6_ASAP7_75t_L g889 ( 
.A(n_625),
.B(n_599),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_746),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_763),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_693),
.B(n_598),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_633),
.Y(n_893)
);

NOR2x1p5_ASAP7_75t_L g894 ( 
.A(n_668),
.B(n_546),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_645),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_699),
.Y(n_896)
);

NOR2x2_ASAP7_75t_L g897 ( 
.A(n_677),
.B(n_599),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_765),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_748),
.B(n_598),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_769),
.B(n_517),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_765),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_764),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_SL g903 ( 
.A1(n_784),
.A2(n_209),
.B1(n_250),
.B2(n_608),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_626),
.A2(n_573),
.B1(n_574),
.B2(n_576),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_769),
.B(n_774),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_765),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_614),
.B(n_546),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_719),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_774),
.B(n_517),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_762),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_777),
.B(n_539),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_760),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_728),
.Y(n_913)
);

AND2x6_ASAP7_75t_L g914 ( 
.A(n_766),
.B(n_599),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_716),
.A2(n_539),
.B(n_562),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_663),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_770),
.B(n_604),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_639),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_SL g919 ( 
.A(n_698),
.B(n_613),
.C(n_609),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_777),
.B(n_539),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_692),
.B(n_673),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_631),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_728),
.B(n_604),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_634),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_673),
.B(n_604),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_719),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_765),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_635),
.B(n_573),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_622),
.A2(n_546),
.B1(n_562),
.B2(n_608),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_635),
.B(n_573),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_637),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_732),
.B(n_574),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_637),
.A2(n_574),
.B1(n_576),
.B2(n_587),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_670),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_676),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_676),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_732),
.B(n_576),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_706),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_706),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_755),
.B(n_546),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_663),
.B(n_587),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_722),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_707),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_SL g944 ( 
.A(n_622),
.B(n_0),
.C(n_1),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_628),
.A2(n_562),
.B1(n_609),
.B2(n_608),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_707),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_709),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_709),
.A2(n_595),
.B1(n_591),
.B2(n_590),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_614),
.A2(n_613),
.B(n_562),
.C(n_591),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_684),
.B(n_587),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_713),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_713),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_724),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_727),
.A2(n_579),
.B(n_591),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_715),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_715),
.A2(n_595),
.B1(n_590),
.B2(n_589),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_670),
.B(n_589),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_729),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_SL g959 ( 
.A(n_628),
.B(n_4),
.C(n_5),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_718),
.Y(n_960)
);

BUFx4f_ASAP7_75t_L g961 ( 
.A(n_718),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_721),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_738),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_686),
.B(n_589),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_627),
.B(n_590),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_689),
.B(n_595),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_721),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_700),
.B(n_579),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_700),
.B(n_579),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_736),
.A2(n_579),
.B(n_419),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_659),
.A2(n_711),
.B1(n_701),
.B2(n_731),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_723),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_723),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_725),
.A2(n_462),
.B1(n_209),
.B2(n_250),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_740),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_725),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_812),
.A2(n_751),
.B(n_775),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_792),
.B(n_659),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_823),
.A2(n_751),
.B(n_782),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_793),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_905),
.A2(n_648),
.B(n_711),
.C(n_701),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_808),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_808),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_808),
.Y(n_984)
);

INVx8_ASAP7_75t_L g985 ( 
.A(n_813),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_916),
.B(n_629),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_795),
.A2(n_780),
.B(n_704),
.C(n_666),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_806),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_916),
.B(n_669),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_795),
.A2(n_752),
.B(n_753),
.C(n_733),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_860),
.B(n_733),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_971),
.A2(n_753),
.B1(n_752),
.B2(n_743),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_860),
.B(n_697),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_L g994 ( 
.A(n_791),
.B(n_685),
.C(n_747),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_794),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_913),
.B(n_734),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_895),
.A2(n_650),
.B(n_662),
.Y(n_997)
);

AOI221xp5_ASAP7_75t_L g998 ( 
.A1(n_800),
.A2(n_910),
.B1(n_806),
.B2(n_822),
.C(n_848),
.Y(n_998)
);

OAI22x1_ASAP7_75t_L g999 ( 
.A1(n_863),
.A2(n_921),
.B1(n_831),
.B2(n_892),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_819),
.B(n_742),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_805),
.A2(n_745),
.B1(n_705),
.B2(n_710),
.Y(n_1001)
);

AOI33xp33_ASAP7_75t_L g1002 ( 
.A1(n_803),
.A2(n_672),
.A3(n_720),
.B1(n_624),
.B2(n_12),
.B3(n_14),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_838),
.B(n_624),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_819),
.B(n_759),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_824),
.A2(n_650),
.B1(n_662),
.B2(n_761),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_845),
.B(n_767),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_814),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_895),
.A2(n_772),
.B(n_714),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_814),
.Y(n_1009)
);

AOI33xp33_ASAP7_75t_L g1010 ( 
.A1(n_816),
.A2(n_7),
.A3(n_9),
.B1(n_10),
.B2(n_15),
.B3(n_17),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_849),
.B(n_671),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_838),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_854),
.B(n_671),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_802),
.B(n_885),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_851),
.A2(n_696),
.B1(n_779),
.B2(n_776),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_825),
.B(n_696),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_799),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_788),
.B(n_786),
.Y(n_1018)
);

OR2x6_ASAP7_75t_SL g1019 ( 
.A(n_853),
.B(n_749),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_788),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_808),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_827),
.B(n_778),
.Y(n_1022)
);

OAI22x1_ASAP7_75t_L g1023 ( 
.A1(n_921),
.A2(n_772),
.B1(n_708),
.B2(n_778),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_885),
.B(n_757),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_827),
.A2(n_735),
.B(n_730),
.C(n_462),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_820),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_800),
.A2(n_462),
.B1(n_250),
.B2(n_209),
.C(n_579),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_809),
.A2(n_579),
.B(n_419),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_846),
.A2(n_462),
.B(n_209),
.C(n_250),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_958),
.B(n_438),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_815),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_841),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_817),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_842),
.B(n_250),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_975),
.B(n_18),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_876),
.B(n_19),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_900),
.A2(n_429),
.B(n_419),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_975),
.B(n_20),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_833),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_890),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_815),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_836),
.B(n_25),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_942),
.A2(n_27),
.B(n_31),
.C(n_32),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_909),
.A2(n_920),
.B(n_911),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_830),
.B(n_438),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_839),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_953),
.A2(n_33),
.B(n_38),
.C(n_39),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_866),
.A2(n_429),
.B(n_419),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_963),
.B(n_40),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_815),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_SL g1051 ( 
.A1(n_848),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_830),
.B(n_438),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_862),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_826),
.Y(n_1054)
);

BUFx4f_ASAP7_75t_L g1055 ( 
.A(n_917),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_801),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_SL g1057 ( 
.A1(n_907),
.A2(n_438),
.B(n_286),
.C(n_419),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_811),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_843),
.B(n_54),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_SL g1060 ( 
.A(n_944),
.B(n_55),
.C(n_56),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_798),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_887),
.A2(n_429),
.B(n_419),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_874),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_880),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_798),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_878),
.A2(n_429),
.B(n_419),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_858),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_886),
.A2(n_915),
.B(n_968),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_857),
.B(n_61),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_944),
.B(n_429),
.C(n_403),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_869),
.B(n_62),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_858),
.A2(n_438),
.B1(n_429),
.B2(n_403),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_959),
.A2(n_286),
.B(n_438),
.C(n_403),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_859),
.B(n_429),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_959),
.A2(n_286),
.B(n_438),
.C(n_403),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_810),
.A2(n_403),
.B(n_286),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_815),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_852),
.B(n_864),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_828),
.B(n_438),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_811),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_829),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_832),
.B(n_286),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_869),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_969),
.A2(n_403),
.B(n_70),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_877),
.B(n_286),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_850),
.A2(n_286),
.B(n_71),
.C(n_81),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_811),
.B(n_65),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_810),
.A2(n_286),
.B(n_96),
.C(n_99),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_847),
.B(n_86),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_868),
.B(n_102),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_877),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_883),
.A2(n_109),
.B1(n_118),
.B2(n_123),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_804),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_891),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_865),
.A2(n_131),
.B1(n_139),
.B2(n_145),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_902),
.A2(n_146),
.B(n_148),
.C(n_152),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_865),
.A2(n_154),
.B(n_156),
.C(n_855),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_842),
.B(n_811),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_801),
.A2(n_965),
.B(n_918),
.C(n_941),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_925),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_835),
.A2(n_949),
.B(n_954),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_972),
.B(n_893),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_917),
.B(n_893),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_917),
.B(n_804),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_949),
.A2(n_970),
.B(n_789),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_922),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_925),
.B(n_923),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_925),
.B(n_923),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_899),
.A2(n_937),
.B(n_932),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_950),
.A2(n_964),
.B(n_966),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_856),
.B(n_881),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_879),
.A2(n_870),
.B(n_940),
.C(n_961),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_961),
.B(n_875),
.Y(n_1114)
);

AO32x1_ASAP7_75t_L g1115 ( 
.A1(n_924),
.A2(n_943),
.A3(n_955),
.B1(n_973),
.B2(n_935),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_SL g1116 ( 
.A1(n_912),
.A2(n_927),
.B(n_870),
.C(n_929),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_818),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_818),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_939),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_818),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_896),
.B(n_908),
.Y(n_1121)
);

OAI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_940),
.A2(n_867),
.B(n_928),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_926),
.B(n_976),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_SL g1124 ( 
.A(n_903),
.B(n_821),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_907),
.B(n_930),
.C(n_945),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_978),
.B(n_946),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_980),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_1022),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1044),
.A2(n_837),
.B(n_888),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_981),
.A2(n_923),
.B(n_967),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_989),
.B(n_962),
.Y(n_1131)
);

O2A1O1Ixp5_ASAP7_75t_SL g1132 ( 
.A1(n_1085),
.A2(n_789),
.B(n_790),
.C(n_934),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_986),
.B(n_934),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1068),
.A2(n_947),
.A3(n_960),
.B(n_882),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_993),
.B(n_821),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1110),
.A2(n_888),
.B(n_871),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1086),
.A2(n_894),
.B(n_919),
.C(n_834),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1009),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1111),
.A2(n_837),
.B(n_871),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1035),
.A2(n_1038),
.B(n_987),
.C(n_994),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_1097),
.A2(n_790),
.B(n_840),
.C(n_912),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1099),
.A2(n_884),
.B(n_834),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_1062),
.A2(n_951),
.B(n_947),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_995),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1008),
.A2(n_957),
.B(n_906),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_985),
.B(n_804),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_1105),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1033),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_988),
.A2(n_875),
.B1(n_872),
.B2(n_906),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1102),
.A2(n_951),
.B(n_960),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1012),
.B(n_1003),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1012),
.B(n_952),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1101),
.B(n_976),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_985),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1104),
.B(n_818),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_985),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1103),
.B(n_952),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1081),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1125),
.A2(n_872),
.B(n_914),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1094),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1125),
.A2(n_914),
.B(n_889),
.Y(n_1161)
);

NAND2xp33_ASAP7_75t_R g1162 ( 
.A(n_1018),
.B(n_957),
.Y(n_1162)
);

BUFx8_ASAP7_75t_L g1163 ( 
.A(n_1020),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1106),
.A2(n_787),
.B(n_796),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1004),
.B(n_875),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1042),
.A2(n_897),
.B(n_927),
.C(n_936),
.Y(n_1166)
);

NAND3x1_ASAP7_75t_L g1167 ( 
.A(n_1010),
.B(n_998),
.C(n_1049),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1000),
.B(n_938),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1083),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1026),
.B(n_1040),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_991),
.B(n_931),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_996),
.B(n_787),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1006),
.B(n_796),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_1105),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1046),
.A2(n_957),
.B(n_807),
.C(n_861),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1058),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1005),
.A2(n_914),
.B(n_889),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1066),
.A2(n_797),
.B(n_873),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1005),
.A2(n_914),
.B(n_889),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_1091),
.B(n_906),
.Y(n_1180)
);

INVx3_ASAP7_75t_SL g1181 ( 
.A(n_1056),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1037),
.A2(n_797),
.B(n_873),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1107),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1055),
.B(n_875),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1028),
.A2(n_1048),
.B(n_1084),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1057),
.A2(n_904),
.B(n_956),
.Y(n_1186)
);

NOR4xp25_ASAP7_75t_L g1187 ( 
.A(n_1060),
.B(n_844),
.C(n_974),
.D(n_933),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1015),
.A2(n_901),
.A3(n_974),
.B(n_904),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_977),
.A2(n_898),
.B(n_901),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_979),
.A2(n_933),
.B(n_948),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1036),
.B(n_948),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1119),
.Y(n_1192)
);

AO21x2_ASAP7_75t_L g1193 ( 
.A1(n_1113),
.A2(n_889),
.B(n_956),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1001),
.A2(n_898),
.B(n_844),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_992),
.A2(n_898),
.B(n_1034),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1001),
.A2(n_898),
.B(n_992),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1082),
.A2(n_1024),
.B(n_1090),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1032),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1023),
.A2(n_1108),
.B(n_1109),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1069),
.B(n_1019),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1064),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1046),
.A2(n_1067),
.B(n_1047),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1051),
.A2(n_1059),
.B1(n_1011),
.B2(n_1071),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1007),
.B(n_999),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1070),
.A2(n_1122),
.B1(n_1065),
.B2(n_1061),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1054),
.B(n_1112),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_982),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1002),
.A2(n_997),
.B(n_1088),
.C(n_1063),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1089),
.A2(n_1072),
.B(n_1117),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_990),
.A2(n_1029),
.A3(n_1025),
.B(n_1115),
.Y(n_1210)
);

O2A1O1Ixp5_ASAP7_75t_L g1211 ( 
.A1(n_1116),
.A2(n_1092),
.B(n_1070),
.C(n_1117),
.Y(n_1211)
);

AOI31xp67_ASAP7_75t_L g1212 ( 
.A1(n_1095),
.A2(n_1079),
.A3(n_1045),
.B(n_1052),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1078),
.B(n_1013),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1096),
.A2(n_1092),
.B(n_1114),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1073),
.A2(n_1075),
.B(n_1027),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1031),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1124),
.A2(n_1115),
.B(n_1074),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1121),
.Y(n_1218)
);

AOI31xp67_ASAP7_75t_L g1219 ( 
.A1(n_1115),
.A2(n_1098),
.A3(n_1030),
.B(n_1013),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1124),
.A2(n_1074),
.B(n_1076),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1123),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1100),
.B(n_1014),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1016),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1016),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1058),
.A2(n_1080),
.A3(n_1053),
.B(n_1039),
.Y(n_1225)
);

AOI221x1_ASAP7_75t_L g1226 ( 
.A1(n_1031),
.A2(n_1118),
.B1(n_1077),
.B2(n_1050),
.C(n_1061),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1016),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1065),
.A2(n_1043),
.B(n_1093),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1080),
.B(n_1041),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1120),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1031),
.A2(n_1050),
.B(n_1077),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1087),
.A2(n_982),
.B1(n_983),
.B2(n_984),
.Y(n_1232)
);

AOI221x1_ASAP7_75t_L g1233 ( 
.A1(n_1050),
.A2(n_1077),
.B1(n_1118),
.B2(n_984),
.C(n_1021),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1074),
.A2(n_1118),
.B(n_983),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1021),
.B(n_978),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1009),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_978),
.B(n_651),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_978),
.A2(n_795),
.B(n_905),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_L g1239 ( 
.A1(n_1097),
.A2(n_1068),
.B(n_1088),
.C(n_1015),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1012),
.B(n_688),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1037),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1012),
.B(n_688),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_978),
.B(n_795),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_L g1244 ( 
.A(n_1056),
.B(n_678),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_985),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_985),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_978),
.B(n_651),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1102),
.A2(n_1068),
.B(n_1106),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1037),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_978),
.A2(n_795),
.B(n_905),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1044),
.A2(n_895),
.B(n_1068),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_978),
.A2(n_971),
.B(n_981),
.C(n_795),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_SL g1253 ( 
.A(n_981),
.B(n_971),
.C(n_905),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1044),
.A2(n_895),
.B(n_1068),
.Y(n_1254)
);

BUFx4_ASAP7_75t_SL g1255 ( 
.A(n_1020),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1037),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1009),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_978),
.A2(n_795),
.B(n_905),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_978),
.B(n_651),
.Y(n_1259)
);

NAND3x1_ASAP7_75t_L g1260 ( 
.A(n_989),
.B(n_971),
.C(n_658),
.Y(n_1260)
);

CKINVDCx6p67_ASAP7_75t_R g1261 ( 
.A(n_985),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_985),
.B(n_660),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1102),
.A2(n_1068),
.B(n_1106),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1068),
.A2(n_1110),
.A3(n_1022),
.B(n_1015),
.Y(n_1264)
);

NOR3xp33_ASAP7_75t_L g1265 ( 
.A(n_981),
.B(n_905),
.C(n_795),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_985),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1017),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1068),
.A2(n_1110),
.A3(n_1022),
.B(n_1015),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1217),
.A2(n_1143),
.B(n_1196),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1251),
.A2(n_1254),
.B(n_1249),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1147),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1254),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1203),
.A2(n_1243),
.B1(n_1258),
.B2(n_1250),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1252),
.A2(n_1140),
.B(n_1238),
.C(n_1253),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1260),
.A2(n_1167),
.B1(n_1259),
.B2(n_1247),
.Y(n_1276)
);

INVx3_ASAP7_75t_SL g1277 ( 
.A(n_1261),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1265),
.A2(n_1202),
.B(n_1175),
.C(n_1253),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1127),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1134),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1138),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1251),
.A2(n_1185),
.B(n_1145),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1145),
.A2(n_1139),
.B(n_1136),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1239),
.A2(n_1265),
.B(n_1179),
.Y(n_1285)
);

OAI22x1_ASAP7_75t_L g1286 ( 
.A1(n_1200),
.A2(n_1133),
.B1(n_1223),
.B2(n_1224),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1134),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1163),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1237),
.B(n_1131),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1133),
.B(n_1235),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1144),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1175),
.A2(n_1208),
.B(n_1239),
.C(n_1177),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1151),
.B(n_1206),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1178),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1139),
.A2(n_1136),
.B(n_1129),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1129),
.A2(n_1182),
.B(n_1209),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1148),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1163),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1217),
.A2(n_1150),
.B(n_1164),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1197),
.A2(n_1189),
.B(n_1190),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1147),
.B(n_1174),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1206),
.B(n_1126),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1135),
.A2(n_1169),
.B1(n_1142),
.B2(n_1267),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1255),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1166),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1211),
.A2(n_1130),
.B(n_1195),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1255),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1178),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1137),
.A2(n_1132),
.B(n_1205),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1236),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1198),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1194),
.B(n_1187),
.C(n_1152),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1159),
.A2(n_1220),
.B(n_1214),
.C(n_1161),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1169),
.B(n_1257),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1128),
.A2(n_1189),
.B(n_1220),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1141),
.A2(n_1152),
.B(n_1228),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1248),
.A2(n_1263),
.B(n_1141),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1158),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1181),
.B(n_1191),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1181),
.A2(n_1245),
.B(n_1146),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1160),
.B(n_1183),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1248),
.A2(n_1263),
.B(n_1186),
.Y(n_1322)
);

AO21x2_ASAP7_75t_L g1323 ( 
.A1(n_1143),
.A2(n_1128),
.B(n_1199),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1165),
.B(n_1204),
.C(n_1227),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1234),
.A2(n_1231),
.B(n_1226),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1171),
.A2(n_1233),
.B(n_1149),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1147),
.B(n_1174),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1172),
.A2(n_1173),
.B(n_1192),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1212),
.A2(n_1244),
.B(n_1157),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1146),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1201),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1246),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1176),
.A2(n_1229),
.B(n_1232),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1222),
.Y(n_1334)
);

AOI221xp5_ASAP7_75t_L g1335 ( 
.A1(n_1213),
.A2(n_1170),
.B1(n_1218),
.B2(n_1153),
.C(n_1168),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1232),
.A2(n_1147),
.B(n_1174),
.C(n_1221),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1174),
.B(n_1155),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_L g1338 ( 
.A(n_1180),
.B(n_1216),
.Y(n_1338)
);

OAI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1180),
.A2(n_1266),
.B(n_1230),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1216),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1193),
.A2(n_1184),
.B(n_1264),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1219),
.A2(n_1210),
.A3(n_1268),
.B(n_1264),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1264),
.A2(n_1268),
.B(n_1210),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1146),
.A2(n_1154),
.B1(n_1156),
.B2(n_1262),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1216),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1262),
.A2(n_1210),
.B(n_1225),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1216),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1264),
.A2(n_1268),
.B(n_1210),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1193),
.A2(n_1188),
.B(n_1225),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1188),
.A2(n_1225),
.B(n_1162),
.Y(n_1350)
);

INVx4_ASAP7_75t_SL g1351 ( 
.A(n_1262),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1154),
.A2(n_1156),
.B1(n_1225),
.B2(n_1162),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1188),
.B(n_1207),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1188),
.A2(n_1252),
.B(n_1253),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1251),
.A2(n_1254),
.B(n_1249),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1260),
.A2(n_1252),
.B(n_1250),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1203),
.A2(n_978),
.B1(n_1243),
.B2(n_1238),
.Y(n_1357)
);

AOI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1217),
.A2(n_1062),
.B(n_1220),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1252),
.A2(n_1253),
.B(n_1250),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1127),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1260),
.A2(n_1238),
.B1(n_1258),
.B2(n_1250),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1252),
.A2(n_978),
.B(n_981),
.C(n_971),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1251),
.A2(n_1254),
.B(n_1249),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1146),
.Y(n_1368)
);

NAND2x1p5_ASAP7_75t_L g1369 ( 
.A(n_1147),
.B(n_1174),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1127),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1261),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1127),
.Y(n_1372)
);

BUFx8_ASAP7_75t_L g1373 ( 
.A(n_1138),
.Y(n_1373)
);

AO21x1_ASAP7_75t_L g1374 ( 
.A1(n_1265),
.A2(n_1203),
.B(n_981),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1203),
.A2(n_978),
.B1(n_1243),
.B2(n_1238),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1203),
.A2(n_971),
.B1(n_792),
.B2(n_993),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1147),
.B(n_1174),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1127),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1217),
.A2(n_1062),
.B(n_1220),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1134),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1175),
.B(n_1146),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_SL g1385 ( 
.A1(n_1252),
.A2(n_1140),
.B(n_1250),
.C(n_1238),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1261),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1260),
.A2(n_1238),
.B1(n_1258),
.B2(n_1250),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1388)
);

AOI21xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1181),
.A2(n_585),
.B(n_678),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1252),
.A2(n_1253),
.B(n_1250),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1252),
.A2(n_1140),
.B(n_1243),
.C(n_1238),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1243),
.B(n_1133),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1249),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1203),
.A2(n_592),
.B1(n_323),
.B2(n_327),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1302),
.B(n_1290),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1283),
.A2(n_1284),
.B(n_1343),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1397),
.B(n_1293),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1388),
.B(n_1314),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1280),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1365),
.A2(n_1376),
.B(n_1385),
.C(n_1362),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1284),
.A2(n_1348),
.B(n_1343),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1399),
.A2(n_1375),
.B1(n_1357),
.B2(n_1365),
.C(n_1276),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1397),
.B(n_1289),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1291),
.B(n_1297),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1274),
.B(n_1360),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1282),
.B(n_1310),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1385),
.A2(n_1393),
.B(n_1275),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1274),
.B(n_1387),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1356),
.A2(n_1396),
.B(n_1279),
.C(n_1305),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1334),
.B(n_1321),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1279),
.A2(n_1292),
.B(n_1336),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1292),
.A2(n_1336),
.B(n_1383),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1303),
.B(n_1318),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1342),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1383),
.A2(n_1301),
.B(n_1327),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1354),
.A2(n_1285),
.B(n_1357),
.C(n_1375),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1373),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1361),
.B(n_1370),
.Y(n_1423)
);

CKINVDCx16_ASAP7_75t_R g1424 ( 
.A(n_1288),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1288),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1342),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1335),
.B(n_1372),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_1374),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1331),
.B(n_1324),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1313),
.A2(n_1309),
.B(n_1329),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1340),
.B(n_1345),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1347),
.B(n_1286),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1373),
.B(n_1339),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1348),
.A2(n_1295),
.B(n_1273),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1337),
.B(n_1332),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1353),
.B(n_1350),
.Y(n_1436)
);

OA22x2_ASAP7_75t_L g1437 ( 
.A1(n_1352),
.A2(n_1316),
.B1(n_1330),
.B2(n_1368),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1389),
.A2(n_1312),
.B(n_1320),
.C(n_1313),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_SL g1439 ( 
.A1(n_1371),
.A2(n_1386),
.B(n_1277),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1373),
.B(n_1328),
.Y(n_1440)
);

AOI21x1_ASAP7_75t_SL g1441 ( 
.A1(n_1371),
.A2(n_1386),
.B(n_1277),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1322),
.A2(n_1317),
.B(n_1296),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1307),
.A2(n_1344),
.B1(n_1304),
.B2(n_1298),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1342),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1298),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1346),
.B(n_1333),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1341),
.B(n_1338),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1304),
.A2(n_1311),
.B1(n_1306),
.B2(n_1369),
.Y(n_1448)
);

O2A1O1Ixp5_ASAP7_75t_L g1449 ( 
.A1(n_1358),
.A2(n_1379),
.B(n_1308),
.C(n_1294),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1301),
.A2(n_1327),
.B(n_1377),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1311),
.A2(n_1306),
.B1(n_1377),
.B2(n_1327),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1306),
.A2(n_1271),
.B1(n_1315),
.B2(n_1270),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1269),
.A2(n_1308),
.B(n_1294),
.C(n_1278),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1349),
.A2(n_1326),
.B(n_1271),
.C(n_1300),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1325),
.B(n_1323),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1270),
.A2(n_1367),
.B1(n_1355),
.B2(n_1299),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1300),
.B(n_1317),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1281),
.A2(n_1287),
.B(n_1382),
.C(n_1296),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1382),
.A2(n_1355),
.B(n_1367),
.C(n_1299),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1359),
.A2(n_1363),
.B(n_1364),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1363),
.A2(n_1364),
.B1(n_1366),
.B2(n_1380),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1366),
.B(n_1380),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1381),
.A2(n_1384),
.B1(n_1390),
.B2(n_1391),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1392),
.B(n_1398),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1392),
.A2(n_1394),
.B1(n_1395),
.B2(n_1398),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1394),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1395),
.B(n_1351),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1365),
.A2(n_1252),
.B(n_1140),
.C(n_1243),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1357),
.A2(n_1375),
.B1(n_1260),
.B2(n_1274),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1365),
.A2(n_1252),
.B(n_1250),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1283),
.A2(n_1284),
.B(n_1343),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1283),
.A2(n_1284),
.B(n_1343),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1365),
.A2(n_1252),
.B(n_1250),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1319),
.B(n_1272),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1288),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1290),
.B(n_1293),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1365),
.A2(n_1252),
.B(n_1250),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1319),
.B(n_1272),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1302),
.B(n_1290),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1280),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1365),
.A2(n_1252),
.B(n_1175),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1302),
.B(n_1290),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1290),
.B(n_1293),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1404),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1414),
.B(n_1410),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1449),
.A2(n_1430),
.B(n_1460),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1456),
.A2(n_1459),
.B(n_1452),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1419),
.B(n_1426),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1420),
.B(n_1417),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1420),
.B(n_1417),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1467),
.Y(n_1491)
);

AOI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1461),
.A2(n_1463),
.B(n_1465),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1428),
.B(n_1418),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1409),
.B(n_1421),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1480),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1409),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1423),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1444),
.B(n_1406),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1406),
.B(n_1457),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1455),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1429),
.Y(n_1501)
);

AND3x2_ASAP7_75t_L g1502 ( 
.A(n_1416),
.B(n_1481),
.C(n_1450),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1447),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1466),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1431),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1440),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1435),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1432),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1475),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1458),
.A2(n_1421),
.B(n_1454),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1436),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1446),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1446),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1414),
.A2(n_1412),
.B(n_1470),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1462),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1415),
.B(n_1413),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1403),
.B(n_1483),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1464),
.B(n_1434),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1458),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1434),
.B(n_1401),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1401),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1427),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1437),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1442),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1454),
.A2(n_1453),
.B(n_1416),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1476),
.B(n_1402),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1503),
.B(n_1408),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1499),
.B(n_1434),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1524),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1499),
.B(n_1401),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1524),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1503),
.B(n_1400),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1524),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1524),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1484),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1493),
.B(n_1500),
.Y(n_1539)
);

AOI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1485),
.A2(n_1407),
.B1(n_1469),
.B2(n_1405),
.C(n_1477),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1500),
.B(n_1478),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1485),
.B(n_1482),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1524),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1516),
.B(n_1474),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1516),
.B(n_1411),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1490),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1507),
.Y(n_1548)
);

OAI211xp5_ASAP7_75t_L g1549 ( 
.A1(n_1514),
.A2(n_1468),
.B(n_1473),
.C(n_1481),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1507),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1518),
.B(n_1472),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1498),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1494),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1494),
.B(n_1479),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1520),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1542),
.B(n_1526),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1539),
.B(n_1516),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_L g1558 ( 
.A1(n_1540),
.A2(n_1514),
.B1(n_1522),
.B2(n_1506),
.C(n_1523),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1547),
.B(n_1489),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1549),
.A2(n_1438),
.B(n_1522),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1527),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1533),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1547),
.B(n_1491),
.Y(n_1564)
);

AOI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1540),
.A2(n_1506),
.B1(n_1510),
.B2(n_1501),
.C(n_1508),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1542),
.B(n_1526),
.Y(n_1566)
);

AOI221x1_ASAP7_75t_L g1567 ( 
.A1(n_1527),
.A2(n_1523),
.B1(n_1443),
.B2(n_1448),
.C(n_1501),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1539),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_L g1569 ( 
.A(n_1549),
.B(n_1513),
.C(n_1512),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1553),
.A2(n_1510),
.B1(n_1508),
.B2(n_1498),
.C(n_1519),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_R g1571 ( 
.A(n_1532),
.B(n_1509),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1534),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1553),
.A2(n_1510),
.B1(n_1525),
.B2(n_1437),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1554),
.A2(n_1510),
.B1(n_1525),
.B2(n_1511),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1554),
.B(n_1486),
.C(n_1498),
.Y(n_1576)
);

AOI33xp33_ASAP7_75t_L g1577 ( 
.A1(n_1528),
.A2(n_1496),
.A3(n_1518),
.B1(n_1505),
.B2(n_1495),
.B3(n_1488),
.Y(n_1577)
);

OAI211xp5_ASAP7_75t_L g1578 ( 
.A1(n_1555),
.A2(n_1521),
.B(n_1492),
.C(n_1515),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1532),
.B(n_1526),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1539),
.B(n_1517),
.Y(n_1580)
);

AOI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1555),
.A2(n_1510),
.B1(n_1519),
.B2(n_1525),
.C(n_1497),
.Y(n_1581)
);

OAI211xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1529),
.A2(n_1543),
.B(n_1531),
.C(n_1535),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1529),
.A2(n_1521),
.B(n_1487),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1548),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1537),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1517),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1545),
.B(n_1517),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1547),
.A2(n_1502),
.B1(n_1525),
.B2(n_1490),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1537),
.Y(n_1591)
);

OAI211xp5_ASAP7_75t_L g1592 ( 
.A1(n_1536),
.A2(n_1528),
.B(n_1530),
.C(n_1538),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1496),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1583),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1583),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1560),
.B(n_1486),
.C(n_1521),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1571),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1577),
.B(n_1548),
.Y(n_1598)
);

AOI21xp33_ASAP7_75t_L g1599 ( 
.A1(n_1558),
.A2(n_1525),
.B(n_1486),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1567),
.A2(n_1489),
.B(n_1490),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1562),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1583),
.Y(n_1602)
);

INVx8_ASAP7_75t_L g1603 ( 
.A(n_1559),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1562),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1583),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1584),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1586),
.B(n_1528),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1586),
.B(n_1530),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1563),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1585),
.B(n_1530),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1563),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1559),
.B(n_1489),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1572),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1585),
.B(n_1538),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1573),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1587),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1591),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1591),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1568),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1589),
.Y(n_1624)
);

INVx3_ASAP7_75t_SL g1625 ( 
.A(n_1557),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1578),
.A2(n_1567),
.B(n_1576),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1561),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1606),
.B(n_1556),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1626),
.B(n_1566),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1625),
.B(n_1588),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1626),
.A2(n_1565),
.B1(n_1570),
.B2(n_1574),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1623),
.B(n_1580),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1604),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1424),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1604),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1610),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1625),
.B(n_1589),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1545),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.B(n_1592),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1599),
.B(n_1579),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1610),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1611),
.B(n_1593),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1612),
.Y(n_1648)
);

OAI21xp33_ASAP7_75t_L g1649 ( 
.A1(n_1596),
.A2(n_1576),
.B(n_1575),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1593),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1612),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1538),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1614),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1598),
.B(n_1541),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1594),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1597),
.B(n_1425),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1614),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1607),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1617),
.B(n_1544),
.Y(n_1659)
);

OAI211xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1596),
.A2(n_1475),
.B(n_1422),
.C(n_1546),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1615),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1615),
.Y(n_1662)
);

NAND4xp25_ASAP7_75t_L g1663 ( 
.A(n_1599),
.B(n_1569),
.C(n_1544),
.D(n_1551),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1616),
.B(n_1541),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1617),
.B(n_1544),
.Y(n_1665)
);

AOI321xp33_ASAP7_75t_L g1666 ( 
.A1(n_1594),
.A2(n_1590),
.A3(n_1551),
.B1(n_1451),
.B2(n_1513),
.C(n_1512),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1600),
.B(n_1425),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1616),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1618),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1653),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1630),
.B(n_1608),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1649),
.C(n_1663),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1669),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1617),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1658),
.A2(n_1600),
.B1(n_1603),
.B2(n_1613),
.Y(n_1675)
);

AOI21xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1638),
.A2(n_1628),
.B(n_1654),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1631),
.B(n_1608),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1629),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1647),
.B(n_1608),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1669),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1639),
.B(n_1609),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1639),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1656),
.B(n_1621),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1635),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1656),
.B(n_1445),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1635),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1627),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1621),
.Y(n_1689)
);

OAI21xp33_ASAP7_75t_SL g1690 ( 
.A1(n_1644),
.A2(n_1609),
.B(n_1621),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1650),
.B(n_1618),
.Y(n_1691)
);

NAND2x1p5_ASAP7_75t_L g1692 ( 
.A(n_1667),
.B(n_1550),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1640),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1645),
.B(n_1619),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1640),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1632),
.B(n_1619),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1445),
.Y(n_1697)
);

OAI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1666),
.A2(n_1582),
.B(n_1590),
.C(n_1536),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1654),
.B(n_1564),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1641),
.Y(n_1700)
);

NOR2xp67_ASAP7_75t_SL g1701 ( 
.A(n_1642),
.B(n_1439),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1632),
.B(n_1620),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1636),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1641),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1634),
.B(n_1620),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1688),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_R g1707 ( 
.A(n_1676),
.B(n_1644),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1684),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1674),
.B(n_1652),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1674),
.B(n_1652),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1688),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1673),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1680),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1692),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1672),
.B(n_1646),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1694),
.B(n_1646),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1659),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1703),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1686),
.Y(n_1720)
);

AO21x1_ASAP7_75t_L g1721 ( 
.A1(n_1671),
.A2(n_1627),
.B(n_1655),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1703),
.Y(n_1722)
);

NOR2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1670),
.B(n_1634),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1683),
.A2(n_1655),
.B(n_1648),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1682),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1687),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1677),
.B(n_1659),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1681),
.B(n_1665),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1681),
.B(n_1665),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1693),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1725),
.B(n_1678),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1721),
.A2(n_1690),
.B1(n_1698),
.B2(n_1602),
.C(n_1605),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1713),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1707),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1713),
.Y(n_1735)
);

OAI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1715),
.A2(n_1683),
.B(n_1682),
.C(n_1697),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1715),
.B(n_1700),
.C(n_1695),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1715),
.A2(n_1701),
.B(n_1675),
.C(n_1602),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1740)
);

AOI21xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1707),
.A2(n_1699),
.B(n_1692),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1708),
.Y(n_1742)
);

OAI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1724),
.A2(n_1699),
.B(n_1689),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1724),
.A2(n_1696),
.B1(n_1702),
.B2(n_1705),
.C(n_1595),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1720),
.A2(n_1699),
.B1(n_1679),
.B2(n_1685),
.Y(n_1745)
);

AOI21xp33_ASAP7_75t_L g1746 ( 
.A1(n_1721),
.A2(n_1704),
.B(n_1702),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1708),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1721),
.A2(n_1595),
.B1(n_1602),
.B2(n_1605),
.C(n_1696),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1719),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1723),
.A2(n_1595),
.B1(n_1605),
.B2(n_1701),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1739),
.Y(n_1751)
);

OAI31xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1736),
.A2(n_1720),
.A3(n_1716),
.B(n_1728),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1733),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1734),
.B(n_1722),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1740),
.B(n_1723),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1731),
.B(n_1716),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1737),
.B(n_1719),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1716),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1749),
.B(n_1735),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1741),
.B(n_1714),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1750),
.B(n_1714),
.Y(n_1761)
);

AO22x1_ASAP7_75t_L g1762 ( 
.A1(n_1757),
.A2(n_1743),
.B1(n_1722),
.B2(n_1714),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1744),
.B(n_1746),
.C(n_1738),
.Y(n_1763)
);

NOR4xp25_ASAP7_75t_L g1764 ( 
.A(n_1759),
.B(n_1712),
.C(n_1742),
.D(n_1747),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1751),
.B(n_1718),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1752),
.A2(n_1750),
.B(n_1732),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1760),
.A2(n_1748),
.B1(n_1714),
.B2(n_1745),
.C(n_1717),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1755),
.A2(n_1711),
.B1(n_1706),
.B2(n_1714),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1754),
.A2(n_1712),
.B(n_1722),
.Y(n_1769)
);

NAND3xp33_ASAP7_75t_L g1770 ( 
.A(n_1756),
.B(n_1722),
.C(n_1711),
.Y(n_1770)
);

OAI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1766),
.A2(n_1706),
.B1(n_1711),
.B2(n_1717),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1763),
.A2(n_1758),
.B(n_1722),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1767),
.A2(n_1758),
.B1(n_1706),
.B2(n_1711),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1764),
.A2(n_1753),
.B(n_1730),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1762),
.A2(n_1770),
.B(n_1765),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1773),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1774),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1771),
.A2(n_1769),
.B(n_1768),
.Y(n_1778)
);

NAND2x1_ASAP7_75t_L g1779 ( 
.A(n_1772),
.B(n_1726),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1775),
.A2(n_1730),
.B(n_1726),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1773),
.A2(n_1706),
.B1(n_1717),
.B2(n_1705),
.C(n_1727),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1781),
.B(n_1718),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1780),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1777),
.B(n_1718),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1778),
.B(n_1727),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1776),
.Y(n_1786)
);

CKINVDCx12_ASAP7_75t_R g1787 ( 
.A(n_1784),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1785),
.B(n_1727),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1783),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1788),
.Y(n_1790)
);

AOI322xp5_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1789),
.A3(n_1786),
.B1(n_1779),
.B2(n_1782),
.C1(n_1787),
.C2(n_1729),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1791),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1791),
.A2(n_1729),
.B(n_1728),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1793),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1792),
.A2(n_1729),
.B1(n_1728),
.B2(n_1710),
.Y(n_1795)
);

NAND5xp2_ASAP7_75t_L g1796 ( 
.A(n_1794),
.B(n_1441),
.C(n_1710),
.D(n_1709),
.E(n_1433),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1795),
.A2(n_1689),
.B1(n_1648),
.B2(n_1668),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1797),
.Y(n_1798)
);

OA21x2_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1796),
.B(n_1710),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1799),
.B(n_1709),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1800),
.A2(n_1709),
.B1(n_1668),
.B2(n_1661),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_1637),
.B1(n_1651),
.B2(n_1662),
.C(n_1657),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1664),
.B(n_1643),
.C(n_1622),
.Y(n_1803)
);


endmodule