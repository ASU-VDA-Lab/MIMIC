module fake_jpeg_26925_n_88 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_16),
.B1(n_6),
.B2(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22x1_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_20),
.B1(n_23),
.B2(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_63)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_51),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_8),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_55),
.B(n_56),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_25),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_46),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_26),
.B(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_76),
.B1(n_66),
.B2(n_69),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_26),
.B1(n_41),
.B2(n_29),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_61),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_71),
.C(n_65),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_78),
.B1(n_74),
.B2(n_63),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_82),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_64),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_60),
.B(n_50),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.C(n_83),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_69),
.B(n_39),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_28),
.B(n_42),
.Y(n_88)
);


endmodule