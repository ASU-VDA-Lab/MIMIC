module fake_jpeg_19565_n_148 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_32),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_80),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_76),
.Y(n_85)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_2),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_73),
.B(n_53),
.C(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_66),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_70),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_106),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_104),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_84),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_62),
.B1(n_54),
.B2(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_103),
.B1(n_65),
.B2(n_69),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_63),
.B1(n_49),
.B2(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_3),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_28),
.B1(n_34),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_52),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_65),
.B(n_71),
.C(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_113),
.Y(n_126)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_67),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_19),
.C(n_21),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_4),
.B1(n_6),
.B2(n_13),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_43),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_14),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_115),
.B1(n_117),
.B2(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_111),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_116),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_134),
.B1(n_137),
.B2(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_135),
.B1(n_126),
.B2(n_124),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_132),
.C(n_128),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_120),
.C(n_110),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_127),
.B(n_125),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_30),
.B(n_31),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_39),
.B(n_131),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_119),
.Y(n_148)
);


endmodule