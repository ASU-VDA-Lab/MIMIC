module fake_netlist_1_7693_n_952 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_952);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_952;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_948;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g113 ( .A(n_38), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_5), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_55), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_58), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_35), .Y(n_120) );
INVx2_ASAP7_75t_SL g121 ( .A(n_91), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_53), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_72), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_99), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_24), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_62), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_10), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_12), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_45), .Y(n_132) );
BUFx5_ASAP7_75t_L g133 ( .A(n_13), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
INVx2_ASAP7_75t_SL g136 ( .A(n_71), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_103), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_18), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_87), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_11), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_13), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_23), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_4), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_35), .Y(n_145) );
INVx1_ASAP7_75t_SL g146 ( .A(n_92), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_16), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_27), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_0), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_52), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_63), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_15), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_41), .Y(n_155) );
INVx1_ASAP7_75t_SL g156 ( .A(n_78), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_31), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_113), .B(n_0), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_113), .B(n_1), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_143), .B(n_1), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_114), .B(n_2), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_114), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_115), .B(n_120), .Y(n_172) );
INVx5_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_121), .B(n_2), .Y(n_176) );
BUFx8_ASAP7_75t_L g177 ( .A(n_121), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_115), .B(n_3), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_136), .B(n_3), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_136), .B(n_4), .Y(n_181) );
AO22x2_ASAP7_75t_L g182 ( .A1(n_176), .A2(n_117), .B1(n_155), .B2(n_148), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_161), .B(n_138), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_176), .A2(n_117), .B1(n_155), .B2(n_148), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_176), .Y(n_186) );
NAND2xp33_ASAP7_75t_SL g187 ( .A(n_163), .B(n_124), .Y(n_187) );
XNOR2xp5_ASAP7_75t_L g188 ( .A(n_161), .B(n_116), .Y(n_188) );
OAI22xp33_ASAP7_75t_SL g189 ( .A1(n_161), .A2(n_150), .B1(n_149), .B2(n_144), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_163), .A2(n_140), .B1(n_131), .B2(n_154), .Y(n_190) );
OAI22xp33_ASAP7_75t_SL g191 ( .A1(n_158), .A2(n_130), .B1(n_127), .B2(n_120), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_163), .A2(n_141), .B1(n_145), .B2(n_151), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_163), .A2(n_141), .B1(n_145), .B2(n_151), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_176), .A2(n_179), .B1(n_181), .B2(n_180), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_170), .B(n_133), .Y(n_197) );
NAND3x1_ASAP7_75t_L g198 ( .A(n_158), .B(n_125), .C(n_129), .Y(n_198) );
OA22x2_ASAP7_75t_L g199 ( .A1(n_170), .A2(n_147), .B1(n_142), .B2(n_125), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_180), .B(n_119), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
BUFx10_ASAP7_75t_L g202 ( .A(n_176), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g203 ( .A1(n_158), .A2(n_157), .B1(n_134), .B2(n_129), .Y(n_203) );
OAI22xp33_ASAP7_75t_R g204 ( .A1(n_164), .A2(n_134), .B1(n_142), .B2(n_147), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_180), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_172), .B(n_133), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_176), .A2(n_137), .B1(n_122), .B2(n_118), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_157), .B1(n_156), .B2(n_146), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_172), .B(n_133), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_171), .B(n_123), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_179), .A2(n_133), .B1(n_157), .B2(n_152), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_172), .B(n_133), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_179), .B(n_157), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_179), .A2(n_133), .B1(n_157), .B2(n_139), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_159), .A2(n_132), .B1(n_128), .B2(n_126), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_179), .A2(n_133), .B1(n_153), .B2(n_7), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_179), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_179), .Y(n_222) );
AO22x2_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g224 ( .A1(n_159), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_181), .B(n_8), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_181), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_181), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_202), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_206), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_188), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_206), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_183), .B(n_165), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_211), .B(n_165), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_215), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_202), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_197), .B(n_165), .Y(n_238) );
XOR2xp5_ASAP7_75t_L g239 ( .A(n_188), .B(n_178), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_186), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_201), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
INVxp33_ASAP7_75t_L g244 ( .A(n_183), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_187), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_225), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_200), .B(n_177), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_202), .Y(n_248) );
XOR2xp5_ASAP7_75t_L g249 ( .A(n_190), .B(n_178), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_197), .B(n_177), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
XOR2xp5_ASAP7_75t_L g252 ( .A(n_189), .B(n_178), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_226), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_215), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_214), .B(n_171), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_214), .B(n_171), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_227), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_199), .Y(n_260) );
INVxp33_ASAP7_75t_L g261 ( .A(n_192), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_229), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_182), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_182), .B(n_14), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_182), .Y(n_266) );
XOR2x2_ASAP7_75t_L g267 ( .A(n_191), .B(n_16), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_182), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_185), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_185), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_218), .B(n_177), .Y(n_271) );
XOR2xp5_ASAP7_75t_L g272 ( .A(n_185), .B(n_17), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_185), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_205), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_205), .B(n_171), .Y(n_276) );
INVxp67_ASAP7_75t_SL g277 ( .A(n_196), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_213), .B(n_177), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_198), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_195), .B(n_18), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_216), .B(n_177), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_223), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_209), .B(n_19), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_223), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_212), .B(n_177), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_203), .B(n_177), .Y(n_288) );
INVxp33_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_223), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_219), .B(n_171), .Y(n_291) );
XOR2xp5_ASAP7_75t_L g292 ( .A(n_208), .B(n_19), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_198), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_204), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_208), .B(n_169), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_251), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_235), .B(n_169), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_235), .B(n_169), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_241), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_238), .B(n_224), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_238), .B(n_20), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_295), .B(n_184), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_230), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_251), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_238), .B(n_184), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_234), .B(n_20), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_265), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_236), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_234), .B(n_21), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_230), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_291), .A2(n_220), .B(n_217), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_237), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_236), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_231), .B(n_21), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_233), .B(n_193), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_240), .B(n_22), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_277), .B(n_193), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_265), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_295), .B(n_22), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_295), .B(n_23), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_262), .B(n_24), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_256), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_241), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_256), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_254), .Y(n_329) );
AND2x2_ASAP7_75t_SL g330 ( .A(n_264), .B(n_164), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_257), .B(n_25), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_242), .A2(n_220), .B(n_217), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g333 ( .A1(n_255), .A2(n_210), .B(n_207), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_257), .B(n_25), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_275), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_274), .B(n_26), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_242), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_243), .A2(n_210), .B(n_207), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_274), .B(n_27), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_243), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_255), .B(n_194), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_237), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_258), .B(n_246), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_244), .B(n_28), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_248), .Y(n_345) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_266), .B(n_164), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_258), .B(n_194), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_294), .B(n_28), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_246), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
INVx6_ASAP7_75t_SL g351 ( .A(n_303), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_297), .B(n_278), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_303), .B(n_268), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_342), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_303), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_337), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_297), .B(n_298), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_297), .B(n_259), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_337), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_349), .Y(n_364) );
AND2x6_ASAP7_75t_L g365 ( .A(n_303), .B(n_283), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_310), .B(n_263), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_310), .B(n_275), .Y(n_368) );
INVx5_ASAP7_75t_L g369 ( .A(n_296), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_297), .B(n_269), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_300), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_298), .B(n_270), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_298), .B(n_260), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_296), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
OR2x6_ASAP7_75t_L g376 ( .A(n_303), .B(n_273), .Y(n_376) );
NOR2xp67_ASAP7_75t_L g377 ( .A(n_303), .B(n_283), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_298), .B(n_253), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_300), .B(n_253), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_300), .B(n_261), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_309), .B(n_272), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_303), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_326), .B(n_249), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_303), .B(n_285), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_383), .B(n_239), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_353), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_369), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
BUFx2_ASAP7_75t_R g391 ( .A(n_383), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_369), .B(n_349), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_369), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_361), .B(n_326), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
BUFx12f_ASAP7_75t_L g398 ( .A(n_356), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_381), .B(n_310), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_369), .Y(n_400) );
BUFx2_ASAP7_75t_SL g401 ( .A(n_369), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_378), .B(n_326), .Y(n_402) );
BUFx2_ASAP7_75t_SL g403 ( .A(n_369), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_351), .Y(n_405) );
INVx8_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_351), .Y(n_407) );
INVx3_ASAP7_75t_SL g408 ( .A(n_356), .Y(n_408) );
CKINVDCx8_ASAP7_75t_R g409 ( .A(n_365), .Y(n_409) );
BUFx12f_ASAP7_75t_L g410 ( .A(n_356), .Y(n_410) );
BUFx5_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_356), .B(n_349), .Y(n_412) );
INVx8_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_353), .Y(n_414) );
CKINVDCx11_ASAP7_75t_R g415 ( .A(n_409), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_387), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_409), .A2(n_272), .B1(n_292), .B2(n_381), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_393), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_411), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_385), .B(n_381), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_398), .A2(n_321), .B1(n_292), .B2(n_267), .Y(n_422) );
INVx6_ASAP7_75t_L g423 ( .A(n_398), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_398), .A2(n_321), .B1(n_267), .B2(n_368), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_406), .A2(n_321), .B1(n_356), .B2(n_335), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_392), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_411), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_406), .A2(n_335), .B1(n_365), .B2(n_348), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_376), .B1(n_410), .B2(n_368), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_411), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_386), .B(n_360), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_411), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_395), .A2(n_289), .B(n_252), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_406), .A2(n_365), .B1(n_348), .B2(n_382), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_411), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_399), .B(n_361), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_408), .A2(n_376), .B1(n_354), .B2(n_382), .Y(n_445) );
BUFx2_ASAP7_75t_SL g446 ( .A(n_411), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_411), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_406), .A2(n_365), .B1(n_348), .B2(n_232), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
INVx8_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_410), .A2(n_368), .B1(n_351), .B2(n_361), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_388), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_399), .B(n_348), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_392), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_410), .A2(n_351), .B1(n_366), .B2(n_239), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_388), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_413), .A2(n_365), .B1(n_232), .B2(n_354), .Y(n_457) );
BUFx12f_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_414), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_423), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_417), .A2(n_344), .B1(n_245), .B2(n_312), .C1(n_309), .C2(n_380), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_416), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_453), .B(n_402), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_458), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_432), .A2(n_351), .B1(n_413), .B2(n_402), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_439), .A2(n_376), .B1(n_354), .B2(n_408), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g467 ( .A1(n_458), .A2(n_413), .B1(n_401), .B2(n_403), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_426), .A2(n_413), .B1(n_402), .B2(n_365), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_448), .A2(n_413), .B1(n_402), .B2(n_365), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_458), .A2(n_376), .B1(n_412), .B2(n_354), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_430), .A2(n_376), .B1(n_412), .B2(n_354), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_422), .A2(n_365), .B1(n_366), .B2(n_378), .Y(n_474) );
OAI222xp33_ASAP7_75t_L g475 ( .A1(n_433), .A2(n_389), .B1(n_394), .B2(n_323), .C1(n_322), .C2(n_366), .Y(n_475) );
BUFx4f_ASAP7_75t_SL g476 ( .A(n_430), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_427), .A2(n_365), .B1(n_378), .B2(n_322), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_457), .A2(n_391), .B1(n_377), .B2(n_323), .Y(n_479) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_455), .A2(n_323), .B(n_322), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_421), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_420), .A2(n_365), .B1(n_378), .B2(n_322), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_424), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_434), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_425), .A2(n_365), .B1(n_378), .B2(n_323), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_424), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_446), .A2(n_401), .B1(n_403), .B2(n_386), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_425), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_437), .A2(n_252), .B(n_336), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_442), .B(n_360), .Y(n_493) );
BUFx8_ASAP7_75t_SL g494 ( .A(n_449), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_446), .A2(n_378), .B1(n_370), .B2(n_372), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_423), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_430), .A2(n_370), .B1(n_372), .B2(n_317), .Y(n_497) );
OAI21xp5_ASAP7_75t_SL g498 ( .A1(n_451), .A2(n_312), .B(n_309), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_423), .A2(n_391), .B1(n_377), .B2(n_395), .Y(n_499) );
BUFx12f_ASAP7_75t_L g500 ( .A(n_423), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_449), .B(n_249), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_436), .A2(n_372), .B1(n_370), .B2(n_317), .Y(n_503) );
OR2x2_ASAP7_75t_SL g504 ( .A(n_436), .B(n_393), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_440), .A2(n_372), .B1(n_370), .B2(n_317), .Y(n_505) );
INVx5_ASAP7_75t_SL g506 ( .A(n_440), .Y(n_506) );
OAI222xp33_ASAP7_75t_L g507 ( .A1(n_419), .A2(n_389), .B1(n_394), .B2(n_405), .C1(n_407), .C2(n_390), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_440), .A2(n_372), .B1(n_370), .B2(n_317), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_447), .B(n_414), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_447), .A2(n_372), .B1(n_370), .B2(n_317), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_419), .A2(n_317), .B1(n_336), .B2(n_339), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_429), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_445), .A2(n_380), .B1(n_386), .B2(n_400), .Y(n_514) );
OAI21xp5_ASAP7_75t_SL g515 ( .A1(n_429), .A2(n_312), .B(n_309), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_443), .A2(n_400), .B1(n_353), .B2(n_357), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_443), .A2(n_400), .B1(n_353), .B2(n_357), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_428), .B(n_357), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_444), .Y(n_519) );
OAI21xp33_ASAP7_75t_L g520 ( .A1(n_444), .A2(n_287), .B(n_285), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_450), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_450), .A2(n_317), .B1(n_339), .B2(n_336), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_438), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_438), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_441), .B(n_357), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_418), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_435), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_441), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_450), .A2(n_407), .B1(n_405), .B2(n_390), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_452), .B(n_414), .Y(n_530) );
BUFx4f_ASAP7_75t_SL g531 ( .A(n_429), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_454), .A2(n_312), .B1(n_339), .B2(n_352), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_429), .B(n_363), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_461), .A2(n_450), .B1(n_415), .B2(n_384), .Y(n_534) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_476), .A2(n_450), .B1(n_435), .B2(n_393), .Y(n_535) );
BUFx2_ASAP7_75t_L g536 ( .A(n_504), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_477), .A2(n_435), .B1(n_245), .B2(n_287), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_480), .A2(n_317), .B1(n_290), .B2(n_384), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_479), .A2(n_384), .B1(n_290), .B2(n_358), .Y(n_539) );
OAI211xp5_ASAP7_75t_L g540 ( .A1(n_480), .A2(n_284), .B(n_281), .C(n_344), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_466), .A2(n_384), .B1(n_358), .B2(n_293), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_502), .A2(n_384), .B1(n_358), .B2(n_280), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_492), .A2(n_384), .B1(n_358), .B2(n_346), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_489), .B(n_452), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_462), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_462), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_472), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_472), .B(n_456), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_478), .Y(n_549) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_510), .A2(n_452), .B(n_456), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_471), .B(n_459), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_474), .A2(n_344), .B1(n_281), .B2(n_324), .C(n_352), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_464), .A2(n_396), .B1(n_393), .B2(n_418), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_464), .A2(n_396), .B1(n_393), .B2(n_418), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_468), .A2(n_346), .B1(n_330), .B2(n_331), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_469), .A2(n_396), .B1(n_363), .B2(n_364), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_478), .B(n_459), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_531), .A2(n_396), .B1(n_431), .B2(n_418), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_499), .A2(n_346), .B1(n_330), .B2(n_331), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_489), .A2(n_396), .B1(n_431), .B2(n_418), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_465), .A2(n_346), .B1(n_330), .B2(n_331), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_467), .A2(n_396), .B1(n_364), .B2(n_375), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_470), .A2(n_363), .B1(n_364), .B2(n_375), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_495), .A2(n_346), .B1(n_330), .B2(n_331), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_485), .A2(n_346), .B1(n_330), .B2(n_334), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_515), .A2(n_364), .B1(n_363), .B2(n_375), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_475), .A2(n_488), .B(n_529), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_482), .A2(n_330), .B1(n_334), .B2(n_344), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_481), .B(n_414), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_489), .A2(n_431), .B1(n_418), .B2(n_319), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_498), .B(n_284), .C(n_324), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_500), .A2(n_375), .B1(n_431), .B2(n_371), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_497), .A2(n_371), .B1(n_301), .B2(n_431), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_471), .B(n_431), .Y(n_574) );
OAI222xp33_ASAP7_75t_L g575 ( .A1(n_496), .A2(n_319), .B1(n_334), .B2(n_301), .C1(n_379), .C2(n_304), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_514), .A2(n_334), .B1(n_319), .B2(n_304), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_481), .B(n_319), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_463), .A2(n_324), .B1(n_349), .B2(n_328), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_473), .A2(n_325), .B1(n_328), .B2(n_340), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_483), .A2(n_301), .B1(n_373), .B2(n_362), .C(n_164), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_521), .A2(n_496), .B1(n_503), .B2(n_511), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_504), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_483), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_486), .B(n_379), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_522), .A2(n_325), .B1(n_328), .B2(n_340), .Y(n_585) );
OA222x2_ASAP7_75t_L g586 ( .A1(n_513), .A2(n_343), .B1(n_373), .B2(n_362), .C1(n_340), .C2(n_374), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_486), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_521), .A2(n_343), .B1(n_374), .B2(n_355), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_505), .A2(n_325), .B1(n_328), .B2(n_343), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_508), .A2(n_325), .B1(n_328), .B2(n_316), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_532), .A2(n_325), .B1(n_328), .B2(n_316), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g592 ( .A1(n_491), .A2(n_276), .B1(n_374), .B2(n_320), .C1(n_341), .C2(n_347), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_501), .B(n_29), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_532), .A2(n_325), .B1(n_328), .B2(n_316), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_500), .A2(n_325), .B1(n_328), .B2(n_316), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_484), .B(n_164), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_512), .A2(n_325), .B1(n_328), .B2(n_316), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_501), .B(n_29), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_519), .A2(n_325), .B1(n_328), .B2(n_306), .Y(n_599) );
OAI211xp5_ASAP7_75t_SL g600 ( .A1(n_460), .A2(n_174), .B(n_333), .C(n_341), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_527), .A2(n_374), .B1(n_367), .B2(n_355), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_519), .A2(n_325), .B1(n_328), .B2(n_306), .Y(n_602) );
OA21x2_ASAP7_75t_L g603 ( .A1(n_523), .A2(n_333), .B(n_174), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_523), .B(n_30), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_494), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_493), .A2(n_276), .B1(n_320), .B2(n_333), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_513), .A2(n_528), .B1(n_524), .B2(n_516), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_484), .B(n_174), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_520), .A2(n_174), .B1(n_271), .B2(n_320), .C(n_347), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_520), .A2(n_174), .B1(n_347), .B2(n_341), .C(n_314), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_524), .B(n_30), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_487), .B(n_167), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_528), .A2(n_306), .B1(n_311), .B2(n_374), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_506), .A2(n_367), .B1(n_355), .B2(n_318), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_487), .B(n_167), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_490), .B(n_31), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_517), .A2(n_306), .B1(n_311), .B2(n_315), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_490), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_518), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_506), .A2(n_367), .B1(n_355), .B2(n_315), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_509), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_533), .B(n_167), .C(n_166), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_525), .B(n_32), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_509), .B(n_32), .Y(n_624) );
AOI221xp5_ASAP7_75t_SL g625 ( .A1(n_507), .A2(n_167), .B1(n_314), .B2(n_36), .C(n_37), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_506), .A2(n_306), .B1(n_311), .B2(n_315), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_506), .A2(n_367), .B1(n_355), .B2(n_315), .Y(n_627) );
OAI21xp5_ASAP7_75t_SL g628 ( .A1(n_530), .A2(n_288), .B(n_282), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_530), .A2(n_367), .B1(n_355), .B2(n_315), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_526), .A2(n_311), .B1(n_315), .B2(n_355), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_526), .A2(n_311), .B1(n_315), .B2(n_355), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_526), .B(n_167), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_526), .A2(n_367), .B1(n_314), .B2(n_329), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_526), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_461), .A2(n_367), .B1(n_327), .B2(n_329), .Y(n_635) );
OA21x2_ASAP7_75t_L g636 ( .A1(n_510), .A2(n_338), .B(n_332), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_621), .B(n_167), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_574), .B(n_167), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_625), .A2(n_167), .B1(n_166), .B2(n_160), .C(n_168), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_619), .B(n_33), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_574), .B(n_167), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_567), .B(n_167), .C(n_166), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_551), .B(n_167), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_592), .A2(n_160), .B(n_166), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_570), .B(n_160), .C(n_166), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_593), .B(n_160), .C(n_166), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_571), .A2(n_302), .B1(n_299), .B2(n_307), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_544), .B(n_367), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_534), .A2(n_302), .B1(n_299), .B2(n_307), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_598), .B(n_160), .C(n_166), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_544), .B(n_160), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_551), .B(n_160), .Y(n_652) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_540), .A2(n_538), .B1(n_635), .B2(n_541), .C(n_543), .Y(n_653) );
AOI21xp5_ASAP7_75t_SL g654 ( .A1(n_605), .A2(n_33), .B(n_34), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_538), .A2(n_318), .B1(n_345), .B2(n_313), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_619), .B(n_34), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_607), .A2(n_299), .B(n_302), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_604), .B(n_160), .C(n_166), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_545), .B(n_160), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_581), .A2(n_318), .B1(n_327), .B2(n_329), .C(n_307), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_545), .B(n_160), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_536), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_535), .B(n_160), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_582), .B(n_37), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_611), .B(n_307), .C(n_302), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_582), .A2(n_38), .B(n_39), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_546), .B(n_39), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_546), .B(n_40), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_553), .B(n_160), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_547), .B(n_40), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_559), .A2(n_305), .B1(n_345), .B2(n_313), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_547), .B(n_166), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_539), .A2(n_302), .B1(n_299), .B2(n_307), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_623), .B(n_42), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_605), .A2(n_299), .B(n_332), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_537), .A2(n_307), .B1(n_327), .B2(n_329), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g677 ( .A1(n_542), .A2(n_329), .B1(n_327), .B2(n_308), .C(n_307), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_624), .A2(n_327), .B1(n_166), .B2(n_168), .C(n_175), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_549), .B(n_166), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_549), .B(n_166), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_618), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_583), .B(n_175), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_552), .A2(n_168), .B1(n_175), .B2(n_173), .C(n_338), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_583), .B(n_175), .Y(n_684) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_575), .A2(n_338), .B(n_332), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_587), .B(n_175), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_587), .B(n_175), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_618), .B(n_175), .Y(n_688) );
NOR2xp33_ASAP7_75t_R g689 ( .A(n_586), .B(n_43), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_554), .B(n_168), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_586), .B(n_175), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_558), .A2(n_168), .B(n_175), .C(n_173), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_548), .B(n_175), .Y(n_693) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_566), .A2(n_250), .B(n_345), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_616), .B(n_308), .C(n_313), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_577), .B(n_44), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_557), .B(n_175), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_622), .B(n_168), .C(n_175), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_584), .B(n_168), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_573), .A2(n_296), .B1(n_342), .B2(n_350), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_622), .B(n_168), .C(n_173), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_600), .B(n_168), .C(n_173), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_569), .B(n_168), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_560), .A2(n_305), .B(n_345), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_579), .B(n_168), .C(n_173), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_572), .B(n_563), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_555), .A2(n_296), .B1(n_342), .B2(n_350), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_596), .B(n_168), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_596), .B(n_173), .Y(n_709) );
OAI21xp33_ASAP7_75t_L g710 ( .A1(n_608), .A2(n_296), .B(n_247), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_620), .B(n_173), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_608), .B(n_173), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_634), .B(n_173), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_550), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_628), .B(n_173), .C(n_296), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g716 ( .A1(n_562), .A2(n_308), .B(n_345), .C(n_313), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_636), .B(n_173), .Y(n_717) );
AOI21xp5_ASAP7_75t_SL g718 ( .A1(n_550), .A2(n_313), .B(n_305), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_588), .B(n_350), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_550), .B(n_46), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_636), .B(n_47), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_636), .B(n_48), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_634), .B(n_49), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_636), .B(n_50), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_606), .B(n_51), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_561), .A2(n_305), .B1(n_342), .B2(n_350), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_629), .B(n_296), .C(n_342), .Y(n_727) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_632), .A2(n_279), .B(n_305), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g729 ( .A1(n_627), .A2(n_350), .B(n_342), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_606), .B(n_54), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_576), .B(n_56), .Y(n_731) );
OAI21xp33_ASAP7_75t_SL g732 ( .A1(n_599), .A2(n_602), .B(n_594), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_612), .B(n_57), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_556), .B(n_59), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_612), .B(n_60), .Y(n_735) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_578), .A2(n_296), .B1(n_342), .B2(n_350), .C(n_286), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_595), .B(n_296), .C(n_342), .Y(n_737) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_589), .A2(n_296), .B1(n_350), .B2(n_342), .C(n_66), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_564), .A2(n_350), .B1(n_342), .B2(n_296), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_614), .B(n_350), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_615), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_681), .B(n_615), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_642), .B(n_609), .C(n_580), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_662), .B(n_632), .Y(n_744) );
NAND4xp75_ASAP7_75t_L g745 ( .A(n_691), .B(n_603), .C(n_591), .D(n_597), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_741), .B(n_603), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_638), .B(n_603), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_638), .B(n_633), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_666), .B(n_617), .C(n_585), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_639), .B(n_613), .C(n_626), .Y(n_750) );
NAND3xp33_ASAP7_75t_SL g751 ( .A(n_689), .B(n_565), .C(n_568), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_643), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_641), .B(n_601), .Y(n_753) );
INVx2_ASAP7_75t_SL g754 ( .A(n_637), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_664), .B(n_590), .Y(n_755) );
OR2x2_ASAP7_75t_L g756 ( .A(n_641), .B(n_610), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_689), .B(n_631), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_714), .B(n_630), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_643), .B(n_61), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_684), .A2(n_350), .B1(n_67), .B2(n_68), .Y(n_760) );
INVx1_ASAP7_75t_SL g761 ( .A(n_652), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_720), .B(n_64), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_720), .B(n_69), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_637), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_653), .B(n_70), .C(n_73), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_684), .B(n_74), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_684), .B(n_75), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_651), .B(n_350), .Y(n_768) );
NAND4xp75_ASAP7_75t_L g769 ( .A(n_663), .B(n_76), .C(n_77), .D(n_79), .Y(n_769) );
NAND4xp75_ASAP7_75t_L g770 ( .A(n_663), .B(n_80), .C(n_81), .D(n_83), .Y(n_770) );
OR2x2_ASAP7_75t_L g771 ( .A(n_672), .B(n_85), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_652), .B(n_86), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_679), .B(n_89), .Y(n_773) );
OAI211xp5_ASAP7_75t_SL g774 ( .A1(n_654), .A2(n_94), .B(n_95), .C(n_96), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_667), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_688), .B(n_98), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_644), .A2(n_100), .B(n_101), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_688), .B(n_102), .Y(n_778) );
INVx2_ASAP7_75t_SL g779 ( .A(n_648), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_704), .A2(n_105), .B1(n_106), .B2(n_107), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_680), .B(n_108), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_668), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_682), .B(n_109), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_686), .B(n_111), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_670), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_651), .B(n_648), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_687), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_677), .A2(n_112), .B1(n_716), .B2(n_729), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_706), .B(n_675), .C(n_715), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_640), .A2(n_656), .B1(n_660), .B2(n_646), .C(n_650), .Y(n_790) );
OAI211xp5_ASAP7_75t_SL g791 ( .A1(n_732), .A2(n_706), .B(n_647), .C(n_678), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_728), .B(n_718), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_728), .B(n_740), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_659), .B(n_661), .Y(n_794) );
INVx3_ASAP7_75t_L g795 ( .A(n_728), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_669), .B(n_690), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_723), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_659), .B(n_661), .Y(n_798) );
NAND4xp75_ASAP7_75t_L g799 ( .A(n_669), .B(n_690), .C(n_711), .D(n_740), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_717), .B(n_697), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_693), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_694), .A2(n_658), .B1(n_674), .B2(n_665), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_721), .B(n_722), .Y(n_803) );
AO21x2_ASAP7_75t_L g804 ( .A1(n_724), .A2(n_703), .B(n_723), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_695), .A2(n_683), .B1(n_655), .B2(n_674), .Y(n_805) );
INVx3_ASAP7_75t_L g806 ( .A(n_713), .Y(n_806) );
OAI211xp5_ASAP7_75t_SL g807 ( .A1(n_649), .A2(n_699), .B(n_685), .C(n_657), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_733), .B(n_712), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_727), .B(n_737), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_698), .B(n_701), .C(n_645), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_696), .A2(n_705), .B1(n_725), .B2(n_730), .Y(n_811) );
NAND4xp75_ASAP7_75t_L g812 ( .A(n_711), .B(n_733), .C(n_734), .D(n_696), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_710), .A2(n_735), .B(n_731), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_708), .B(n_709), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_700), .B(n_719), .Y(n_815) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_692), .B(n_702), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_739), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_707), .B(n_734), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_736), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_738), .B(n_676), .C(n_726), .Y(n_820) );
NAND4xp25_ASAP7_75t_L g821 ( .A(n_673), .B(n_642), .C(n_653), .D(n_654), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_671), .B(n_662), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_691), .B(n_642), .C(n_666), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_681), .Y(n_824) );
AO21x2_ASAP7_75t_L g825 ( .A1(n_717), .A2(n_722), .B(n_721), .Y(n_825) );
XOR2x2_ASAP7_75t_L g826 ( .A(n_812), .B(n_823), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_775), .B(n_782), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_744), .B(n_824), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_785), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_744), .B(n_742), .Y(n_830) );
OR2x2_ASAP7_75t_L g831 ( .A(n_742), .B(n_752), .Y(n_831) );
NAND4xp75_ASAP7_75t_L g832 ( .A(n_757), .B(n_796), .C(n_816), .D(n_792), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_792), .B(n_747), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_808), .B(n_751), .Y(n_834) );
INVx1_ASAP7_75t_SL g835 ( .A(n_761), .Y(n_835) );
XNOR2xp5_ASAP7_75t_L g836 ( .A(n_808), .B(n_821), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_817), .B(n_801), .Y(n_837) );
AO22x2_ASAP7_75t_L g838 ( .A1(n_795), .A2(n_779), .B1(n_793), .B2(n_789), .Y(n_838) );
XOR2x2_ASAP7_75t_L g839 ( .A(n_765), .B(n_757), .Y(n_839) );
XNOR2xp5_ASAP7_75t_L g840 ( .A(n_745), .B(n_802), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_747), .B(n_797), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_796), .A2(n_799), .B(n_788), .Y(n_842) );
XOR2x2_ASAP7_75t_L g843 ( .A(n_749), .B(n_769), .Y(n_843) );
XNOR2x2_ASAP7_75t_L g844 ( .A(n_809), .B(n_790), .Y(n_844) );
NAND4xp75_ASAP7_75t_L g845 ( .A(n_822), .B(n_819), .C(n_818), .D(n_815), .Y(n_845) );
NAND4xp75_ASAP7_75t_L g846 ( .A(n_818), .B(n_815), .C(n_763), .D(n_762), .Y(n_846) );
NAND2xp33_ASAP7_75t_R g847 ( .A(n_786), .B(n_795), .Y(n_847) );
INVx1_ASAP7_75t_SL g848 ( .A(n_759), .Y(n_848) );
BUFx12f_ASAP7_75t_L g849 ( .A(n_771), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_786), .Y(n_850) );
NAND2x1_ASAP7_75t_L g851 ( .A(n_786), .B(n_795), .Y(n_851) );
XOR2xp5_ASAP7_75t_L g852 ( .A(n_814), .B(n_755), .Y(n_852) );
INVxp67_ASAP7_75t_L g853 ( .A(n_756), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_791), .A2(n_807), .B1(n_764), .B2(n_754), .Y(n_854) );
INVx1_ASAP7_75t_SL g855 ( .A(n_759), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_787), .B(n_804), .Y(n_856) );
INVx1_ASAP7_75t_SL g857 ( .A(n_754), .Y(n_857) );
INVxp67_ASAP7_75t_SL g858 ( .A(n_768), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_806), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_800), .Y(n_860) );
INVx3_ASAP7_75t_L g861 ( .A(n_797), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_800), .Y(n_862) );
NAND4xp75_ASAP7_75t_SL g863 ( .A(n_762), .B(n_763), .C(n_767), .D(n_766), .Y(n_863) );
INVx5_ASAP7_75t_L g864 ( .A(n_766), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_797), .B(n_804), .Y(n_865) );
NAND4xp75_ASAP7_75t_L g866 ( .A(n_748), .B(n_803), .C(n_777), .D(n_758), .Y(n_866) );
INVxp67_ASAP7_75t_L g867 ( .A(n_748), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_798), .Y(n_868) );
NAND4xp75_ASAP7_75t_L g869 ( .A(n_758), .B(n_772), .C(n_753), .D(n_768), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_825), .B(n_798), .Y(n_870) );
OR2x2_ASAP7_75t_L g871 ( .A(n_746), .B(n_825), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_806), .B(n_813), .Y(n_872) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_813), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_794), .B(n_811), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_840), .B(n_810), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_837), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_829), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_871), .B(n_820), .Y(n_878) );
OAI22xp33_ASAP7_75t_SL g879 ( .A1(n_851), .A2(n_780), .B1(n_783), .B2(n_760), .Y(n_879) );
INVx1_ASAP7_75t_SL g880 ( .A(n_835), .Y(n_880) );
XOR2x2_ASAP7_75t_L g881 ( .A(n_826), .B(n_770), .Y(n_881) );
BUFx3_ASAP7_75t_L g882 ( .A(n_859), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_868), .Y(n_883) );
XOR2x2_ASAP7_75t_L g884 ( .A(n_826), .B(n_805), .Y(n_884) );
INVx1_ASAP7_75t_SL g885 ( .A(n_857), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_827), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_853), .B(n_811), .Y(n_887) );
XNOR2xp5_ASAP7_75t_L g888 ( .A(n_845), .B(n_805), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_831), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_860), .Y(n_890) );
INVx2_ASAP7_75t_SL g891 ( .A(n_859), .Y(n_891) );
XNOR2x2_ASAP7_75t_L g892 ( .A(n_844), .B(n_750), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_862), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_828), .Y(n_894) );
NOR2x1_ASAP7_75t_L g895 ( .A(n_832), .B(n_774), .Y(n_895) );
XOR2x2_ASAP7_75t_L g896 ( .A(n_844), .B(n_743), .Y(n_896) );
BUFx2_ASAP7_75t_L g897 ( .A(n_833), .Y(n_897) );
XOR2x2_ASAP7_75t_L g898 ( .A(n_836), .B(n_776), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_839), .A2(n_778), .B1(n_773), .B2(n_781), .Y(n_899) );
XNOR2xp5_ASAP7_75t_L g900 ( .A(n_839), .B(n_784), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_833), .B(n_870), .Y(n_901) );
INVxp67_ASAP7_75t_L g902 ( .A(n_873), .Y(n_902) );
AO22x2_ASAP7_75t_L g903 ( .A1(n_878), .A2(n_872), .B1(n_850), .B2(n_846), .Y(n_903) );
NAND2xp5_ASAP7_75t_SL g904 ( .A(n_879), .B(n_854), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_896), .A2(n_842), .B1(n_843), .B2(n_834), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_876), .B(n_867), .Y(n_906) );
OA22x2_ASAP7_75t_L g907 ( .A1(n_888), .A2(n_850), .B1(n_852), .B2(n_872), .Y(n_907) );
AO22x2_ASAP7_75t_L g908 ( .A1(n_891), .A2(n_874), .B1(n_869), .B2(n_866), .Y(n_908) );
AO22x1_ASAP7_75t_L g909 ( .A1(n_895), .A2(n_864), .B1(n_858), .B2(n_865), .Y(n_909) );
OA22x2_ASAP7_75t_L g910 ( .A1(n_900), .A2(n_865), .B1(n_870), .B2(n_873), .Y(n_910) );
AOI22x1_ASAP7_75t_L g911 ( .A1(n_892), .A2(n_838), .B1(n_847), .B2(n_861), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_896), .A2(n_843), .B1(n_847), .B2(n_838), .Y(n_912) );
OA22x2_ASAP7_75t_L g913 ( .A1(n_892), .A2(n_899), .B1(n_887), .B2(n_880), .Y(n_913) );
OA22x2_ASAP7_75t_L g914 ( .A1(n_897), .A2(n_885), .B1(n_901), .B2(n_884), .Y(n_914) );
INVx3_ASAP7_75t_L g915 ( .A(n_882), .Y(n_915) );
AO22x2_ASAP7_75t_L g916 ( .A1(n_891), .A2(n_863), .B1(n_838), .B2(n_871), .Y(n_916) );
AOI22x1_ASAP7_75t_SL g917 ( .A1(n_884), .A2(n_848), .B1(n_855), .B2(n_861), .Y(n_917) );
AO22x1_ASAP7_75t_L g918 ( .A1(n_875), .A2(n_864), .B1(n_861), .B2(n_856), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_906), .Y(n_919) );
OAI22xp5_ASAP7_75t_SL g920 ( .A1(n_905), .A2(n_875), .B1(n_898), .B2(n_849), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_915), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_911), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_916), .Y(n_923) );
AOI322xp5_ASAP7_75t_L g924 ( .A1(n_904), .A2(n_902), .A3(n_894), .B1(n_889), .B2(n_886), .C1(n_841), .C2(n_830), .Y(n_924) );
INVx2_ASAP7_75t_SL g925 ( .A(n_916), .Y(n_925) );
INVx1_ASAP7_75t_SL g926 ( .A(n_917), .Y(n_926) );
HB1xp67_ASAP7_75t_SL g927 ( .A(n_913), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_920), .A2(n_912), .B1(n_914), .B2(n_907), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_921), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_921), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_919), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_925), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_929), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_928), .A2(n_927), .B1(n_926), .B2(n_908), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_930), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_934), .A2(n_922), .B1(n_925), .B2(n_932), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_933), .A2(n_922), .B1(n_932), .B2(n_881), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_935), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_938), .Y(n_939) );
BUFx2_ASAP7_75t_L g940 ( .A(n_937), .Y(n_940) );
INVxp67_ASAP7_75t_L g941 ( .A(n_939), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_940), .A2(n_936), .B1(n_931), .B2(n_923), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_941), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_942), .Y(n_944) );
OAI22x1_ASAP7_75t_L g945 ( .A1(n_944), .A2(n_923), .B1(n_902), .B2(n_924), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_945), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_946), .A2(n_943), .B1(n_881), .B2(n_910), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_947), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_948), .A2(n_903), .B1(n_882), .B2(n_890), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_949), .Y(n_950) );
AOI221x1_ASAP7_75t_L g951 ( .A1(n_950), .A2(n_903), .B1(n_877), .B2(n_898), .C(n_893), .Y(n_951) );
AOI211xp5_ASAP7_75t_L g952 ( .A1(n_951), .A2(n_909), .B(n_918), .C(n_883), .Y(n_952) );
endmodule