module real_jpeg_23769_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_173;
wire n_40;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_0),
.A2(n_44),
.B1(n_61),
.B2(n_62),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_69),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_27),
.C(n_39),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_108),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_115),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_5),
.A2(n_24),
.B1(n_126),
.B2(n_213),
.Y(n_216)
);

INVx8_ASAP7_75t_SL g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_71),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_10),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_81)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_11),
.B(n_61),
.C(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_79),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_12),
.A2(n_67),
.B1(n_79),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_79),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_119),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_119),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_119),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_15),
.Y(n_126)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_15),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_149),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_20),
.B(n_121),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_96),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_21),
.B(n_82),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_22),
.B(n_52),
.C(n_72),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_23),
.B(n_36),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_24),
.A2(n_89),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_24),
.A2(n_85),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_24),
.A2(n_206),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_24),
.A2(n_33),
.B(n_89),
.Y(n_232)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_25),
.B(n_34),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_25),
.A2(n_31),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_25),
.A2(n_173),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_26),
.B(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_28),
.Y(n_214)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_45),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_37),
.B(n_50),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_37),
.A2(n_47),
.B1(n_192),
.B2(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_37),
.B(n_108),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_40),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_42),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_41),
.A2(n_76),
.B(n_228),
.C(n_230),
.Y(n_227)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_42),
.B(n_188),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g230 ( 
.A(n_42),
.B(n_61),
.C(n_75),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_46),
.A2(n_130),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_46),
.A2(n_93),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_46),
.A2(n_93),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_47),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_47),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_72),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_69),
.B2(n_70),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_53),
.Y(n_120)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_54),
.B(n_108),
.CON(n_107),
.SN(n_107)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_57),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_69),
.B1(n_107),
.B2(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_65),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_62),
.B(n_107),
.C(n_109),
.Y(n_106)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g229 ( 
.A(n_62),
.B(n_108),
.CON(n_229),
.SN(n_229)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_69),
.B(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_70),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B(n_80),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_73),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_73),
.A2(n_112),
.B1(n_115),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_73),
.A2(n_115),
.B1(n_178),
.B2(n_229),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_77),
.A2(n_113),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_78),
.B(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_91),
.B2(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_95),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_90),
.A2(n_102),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_93),
.B(n_157),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_96),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_110),
.C(n_116),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_97),
.A2(n_98),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_106),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_108),
.B(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_110),
.B(n_116),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_118),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_148),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_132),
.B1(n_146),
.B2(n_147),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_140),
.B1(n_141),
.B2(n_145),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_180),
.B(n_262),
.C(n_266),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_165),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_152),
.B(n_165),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_154),
.B(n_155),
.C(n_162),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_170),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_166),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_168),
.B(n_170),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_176),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_171),
.A2(n_174),
.B1(n_175),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_261),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_256),
.B(n_260),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_240),
.B(n_255),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_223),
.B(n_239),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_202),
.B(n_222),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_189),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_197),
.C(n_200),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_209),
.B(n_221),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_208),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_215),
.B(n_220),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_238),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_233),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_234),
.C(n_235),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_242),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_250),
.C(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);


endmodule