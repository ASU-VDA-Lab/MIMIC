module fake_netlist_6_1640_n_1545 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1545);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1545;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_77),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_31),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_53),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_42),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_49),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_55),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_70),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_106),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_75),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_59),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_1),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_71),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_68),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_130),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_62),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_81),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_97),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_13),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_44),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_37),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_14),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_84),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_22),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_0),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_94),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_27),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_8),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_98),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_37),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_24),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_40),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_18),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_140),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_133),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_38),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_147),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_56),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_33),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_100),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_45),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_39),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_42),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_28),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_91),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_114),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_54),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_17),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_85),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_112),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_73),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_11),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_58),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_88),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_113),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_27),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_115),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_104),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_123),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_43),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_36),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_26),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_87),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_44),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_93),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_125),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_105),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_2),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_124),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_119),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_82),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_96),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_111),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_16),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_90),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_107),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_11),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_9),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_34),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_32),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_51),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_24),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_63),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_65),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_53),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_83),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_2),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_121),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_131),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_10),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_136),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_66),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_151),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_163),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_161),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_153),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_153),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_186),
.B(n_5),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_164),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_197),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_171),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_214),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_154),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_154),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_170),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_296),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_170),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_173),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_174),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_175),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_205),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_180),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_167),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_179),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_157),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_275),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_251),
.B(n_7),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_156),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_181),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_179),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_275),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_188),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_190),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_186),
.B(n_212),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_258),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_200),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_251),
.B(n_12),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_162),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_209),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_216),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_219),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_159),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_189),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_206),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_225),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_159),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_228),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_206),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_236),
.Y(n_358)
);

BUFx6f_ASAP7_75t_SL g359 ( 
.A(n_205),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_192),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_166),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_240),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_242),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_166),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_249),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_250),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_176),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_176),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_253),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_196),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_178),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_178),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_182),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_259),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_182),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_264),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_323),
.B(n_212),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_305),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_306),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_325),
.Y(n_385)
);

BUFx8_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_310),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_313),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_241),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_268),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_320),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_322),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_325),
.B(n_168),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_324),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_241),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_335),
.B(n_206),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_312),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_311),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_309),
.B(n_298),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_333),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_314),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_315),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_205),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_316),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_371),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_298),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_337),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_316),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_317),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_317),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_318),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_319),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_319),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_326),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_326),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_364),
.B(n_158),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_334),
.B(n_235),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_338),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_343),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_348),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_342),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_338),
.B(n_235),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_328),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

BUFx4f_ASAP7_75t_L g450 ( 
.A(n_391),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_335),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_403),
.A2(n_307),
.B1(n_346),
.B2(n_331),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_350),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_382),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_332),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_406),
.B(n_360),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_409),
.A2(n_327),
.B1(n_308),
.B2(n_287),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_407),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_416),
.B(n_235),
.Y(n_462)
);

AND3x2_ASAP7_75t_L g463 ( 
.A(n_381),
.B(n_327),
.C(n_247),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_358),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_390),
.B(n_365),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_444),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_377),
.B(n_366),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_380),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_383),
.B(n_374),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_390),
.B(n_376),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_391),
.B(n_353),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_391),
.B(n_357),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

NOR2x1p5_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_185),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_387),
.B(n_349),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_445),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_341),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_391),
.A2(n_194),
.B1(n_287),
.B2(n_269),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_391),
.B(n_184),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_381),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_L g488 ( 
.A1(n_439),
.A2(n_203),
.B1(n_301),
.B2(n_297),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_391),
.B(n_303),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_389),
.B(n_354),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_441),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_439),
.B(n_194),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_419),
.B(n_152),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_392),
.B(n_344),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_393),
.B(n_369),
.Y(n_495)
);

BUFx4f_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_392),
.B(n_344),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_379),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_395),
.B(n_363),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_441),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_416),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_441),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_384),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_386),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_379),
.B(n_270),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_388),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_385),
.B(n_345),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_400),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_396),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_445),
.B(n_345),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_445),
.A2(n_239),
.B1(n_269),
.B2(n_213),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_L g522 ( 
.A(n_398),
.B(n_268),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_401),
.B(n_412),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_397),
.B(n_272),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_402),
.B(n_273),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_402),
.B(n_404),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_404),
.B(n_274),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_411),
.A2(n_213),
.B1(n_278),
.B2(n_239),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_423),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_415),
.A2(n_260),
.B1(n_195),
.B2(n_243),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_415),
.B(n_152),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_418),
.B(n_276),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_418),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_420),
.B(n_289),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_421),
.B(n_268),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_155),
.Y(n_541)
);

BUFx8_ASAP7_75t_SL g542 ( 
.A(n_408),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_424),
.B(n_356),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_155),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_386),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

INVx3_ASAP7_75t_R g547 ( 
.A(n_432),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_442),
.B(n_362),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_413),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_425),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_427),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_443),
.B(n_291),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_429),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_429),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_430),
.B(n_299),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_426),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_427),
.B(n_405),
.Y(n_560)
);

BUFx4f_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

CKINVDCx11_ASAP7_75t_R g562 ( 
.A(n_433),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_385),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_434),
.B(n_302),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_423),
.A2(n_207),
.B1(n_278),
.B2(n_260),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_438),
.B(n_160),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_434),
.B(n_160),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_434),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_434),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_386),
.B(n_288),
.Y(n_574)
);

BUFx4f_ASAP7_75t_L g575 ( 
.A(n_414),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_419),
.B(n_359),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_419),
.B(n_288),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_414),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_419),
.Y(n_579)
);

AND3x2_ASAP7_75t_L g580 ( 
.A(n_414),
.B(n_233),
.C(n_247),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_428),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_428),
.Y(n_582)
);

AND3x4_ASAP7_75t_L g583 ( 
.A(n_428),
.B(n_208),
.C(n_221),
.Y(n_583)
);

AND2x4_ASAP7_75t_SL g584 ( 
.A(n_482),
.B(n_288),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_499),
.B(n_165),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_457),
.B(n_288),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_458),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_558),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_482),
.A2(n_233),
.B1(n_257),
.B2(n_266),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_450),
.B(n_268),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_469),
.Y(n_591)
);

BUFx5_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

AND2x6_ASAP7_75t_SL g593 ( 
.A(n_481),
.B(n_185),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_512),
.B(n_199),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_578),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_450),
.B(n_268),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_169),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_581),
.B(n_169),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_455),
.B(n_172),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_496),
.B(n_257),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_512),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_506),
.B(n_266),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_465),
.B(n_201),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_496),
.B(n_177),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_506),
.A2(n_237),
.B1(n_183),
.B2(n_295),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_476),
.B(n_177),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_578),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_464),
.B(n_202),
.Y(n_611)
);

NOR2x1p5_ASAP7_75t_L g612 ( 
.A(n_451),
.B(n_211),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_485),
.B(n_183),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_502),
.A2(n_462),
.B1(n_452),
.B2(n_467),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_510),
.B(n_191),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_460),
.B(n_187),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_462),
.A2(n_191),
.B1(n_204),
.B2(n_217),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_471),
.B(n_215),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_505),
.B(n_218),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_480),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_505),
.B(n_220),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_460),
.B(n_245),
.Y(n_624)
);

OAI221xp5_ASAP7_75t_L g625 ( 
.A1(n_567),
.A2(n_210),
.B1(n_195),
.B2(n_198),
.C(n_207),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_582),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_511),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_519),
.B(n_223),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_583),
.A2(n_252),
.B1(n_292),
.B2(n_294),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_519),
.B(n_223),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_446),
.B(n_222),
.Y(n_632)
);

NOR2xp67_ASAP7_75t_L g633 ( 
.A(n_543),
.B(n_431),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_513),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_519),
.B(n_237),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_487),
.B(n_224),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_513),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_519),
.B(n_571),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_514),
.B(n_267),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_462),
.A2(n_293),
.B1(n_279),
.B2(n_277),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_560),
.A2(n_480),
.B1(n_462),
.B2(n_524),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

OAI221xp5_ASAP7_75t_L g643 ( 
.A1(n_520),
.A2(n_198),
.B1(n_210),
.B2(n_243),
.C(n_244),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_492),
.A2(n_277),
.B1(n_279),
.B2(n_281),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_516),
.A2(n_295),
.B1(n_293),
.B2(n_281),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_517),
.B(n_431),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_494),
.B(n_435),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_521),
.B(n_528),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_SL g649 ( 
.A(n_509),
.B(n_244),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_475),
.B(n_226),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_525),
.A2(n_359),
.B1(n_436),
.B2(n_435),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_546),
.Y(n_653)
);

BUFx6f_ASAP7_75t_SL g654 ( 
.A(n_566),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_489),
.B(n_493),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_534),
.B(n_227),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_537),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_497),
.B(n_229),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_542),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_537),
.B(n_230),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_539),
.A2(n_255),
.B1(n_290),
.B2(n_286),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_451),
.B(n_284),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_477),
.A2(n_256),
.B1(n_280),
.B2(n_271),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_550),
.B(n_282),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_527),
.A2(n_265),
.B1(n_263),
.B2(n_262),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_553),
.B(n_261),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_535),
.B(n_538),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_557),
.B(n_254),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_483),
.A2(n_248),
.B1(n_246),
.B2(n_238),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_550),
.A2(n_232),
.B1(n_231),
.B2(n_234),
.Y(n_670)
);

INVxp67_ASAP7_75t_R g671 ( 
.A(n_547),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_551),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_551),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_673)
);

NAND2x1_ASAP7_75t_L g674 ( 
.A(n_448),
.B(n_67),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_566),
.B(n_21),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_497),
.B(n_23),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_534),
.B(n_69),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_554),
.B(n_78),
.Y(n_678)
);

NAND2x1_ASAP7_75t_L g679 ( 
.A(n_448),
.B(n_60),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_556),
.B(n_86),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_492),
.B(n_25),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_534),
.B(n_148),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_565),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_546),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_572),
.B(n_143),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_526),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_563),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_565),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_568),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_518),
.B(n_141),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_568),
.B(n_518),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_564),
.B(n_139),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_533),
.B(n_128),
.Y(n_694)
);

BUFx12f_ASAP7_75t_L g695 ( 
.A(n_562),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_533),
.B(n_127),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_484),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_558),
.B(n_126),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_558),
.B(n_122),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_558),
.B(n_117),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_541),
.B(n_102),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_558),
.B(n_101),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_541),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_559),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_544),
.B(n_569),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_504),
.B(n_29),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_575),
.B(n_30),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_575),
.B(n_38),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_559),
.B(n_54),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_40),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_522),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_449),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_488),
.A2(n_569),
.B(n_540),
.C(n_570),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_575),
.B(n_41),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_478),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_561),
.B(n_47),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_461),
.B(n_48),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_706),
.B(n_523),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_591),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_606),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_653),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_706),
.B(n_459),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_641),
.A2(n_545),
.B1(n_509),
.B2(n_493),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_706),
.B(n_493),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_461),
.Y(n_726)
);

INVx5_ASAP7_75t_L g727 ( 
.A(n_691),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_703),
.B(n_604),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_684),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_655),
.A2(n_579),
.B(n_447),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_588),
.A2(n_603),
.B(n_701),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_602),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_591),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_603),
.A2(n_447),
.B(n_448),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_587),
.B(n_500),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_708),
.A2(n_709),
.B(n_717),
.C(n_711),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_701),
.A2(n_448),
.B(n_472),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_632),
.B(n_495),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_602),
.B(n_490),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_688),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_619),
.B(n_548),
.Y(n_741)
);

O2A1O1Ixp5_ASAP7_75t_L g742 ( 
.A1(n_601),
.A2(n_616),
.B(n_600),
.C(n_609),
.Y(n_742)
);

AOI21x1_ASAP7_75t_L g743 ( 
.A1(n_646),
.A2(n_456),
.B(n_454),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_636),
.B(n_529),
.C(n_463),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_586),
.B(n_508),
.Y(n_745)
);

OAI321xp33_ASAP7_75t_L g746 ( 
.A1(n_686),
.A2(n_574),
.A3(n_530),
.B1(n_532),
.B2(n_577),
.C(n_573),
.Y(n_746)
);

OAI21xp33_ASAP7_75t_L g747 ( 
.A1(n_681),
.A2(n_549),
.B(n_508),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_633),
.B(n_573),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_617),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_692),
.B(n_507),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_659),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_648),
.A2(n_473),
.B(n_479),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_594),
.B(n_583),
.Y(n_753)
);

AO32x2_ASAP7_75t_L g754 ( 
.A1(n_630),
.A2(n_583),
.A3(n_580),
.B1(n_547),
.B2(n_50),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_647),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_709),
.A2(n_491),
.B(n_503),
.C(n_501),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_607),
.A2(n_470),
.B(n_479),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_651),
.A2(n_549),
.B(n_466),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_695),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_607),
.A2(n_470),
.B(n_473),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_615),
.A2(n_545),
.B1(n_509),
.B2(n_576),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_695),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_614),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_662),
.B(n_466),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_717),
.A2(n_491),
.B(n_501),
.C(n_507),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_668),
.B(n_628),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_694),
.A2(n_545),
.B1(n_509),
.B2(n_468),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_657),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_498),
.B1(n_468),
.B2(n_472),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_713),
.A2(n_498),
.B(n_50),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_676),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_596),
.A2(n_696),
.B(n_694),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_624),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_696),
.A2(n_51),
.B1(n_498),
.B2(n_691),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_696),
.A2(n_693),
.B(n_585),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_658),
.B(n_584),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_642),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_629),
.A2(n_631),
.B(n_635),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_584),
.B(n_621),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_666),
.B(n_665),
.C(n_670),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_691),
.B(n_592),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_683),
.B(n_689),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_690),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_716),
.B(n_712),
.C(n_672),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_656),
.A2(n_678),
.B(n_680),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_650),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_677),
.A2(n_685),
.B(n_682),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_677),
.A2(n_685),
.B(n_682),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_597),
.B(n_598),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_SL g790 ( 
.A1(n_675),
.A2(n_715),
.B(n_613),
.C(n_623),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_599),
.A2(n_605),
.B1(n_622),
.B2(n_613),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_622),
.Y(n_792)
);

AOI21x1_ASAP7_75t_L g793 ( 
.A1(n_704),
.A2(n_705),
.B(n_627),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_660),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_589),
.A2(n_640),
.B1(n_618),
.B2(n_608),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_707),
.B(n_644),
.C(n_625),
.Y(n_796)
);

NAND2x1_ASAP7_75t_L g797 ( 
.A(n_687),
.B(n_627),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_592),
.B(n_664),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_669),
.B(n_652),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_592),
.B(n_620),
.Y(n_800)
);

AOI22x1_ASAP7_75t_L g801 ( 
.A1(n_595),
.A2(n_626),
.B1(n_610),
.B2(n_612),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_673),
.A2(n_643),
.B1(n_592),
.B2(n_698),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_671),
.B(n_661),
.Y(n_803)
);

NOR2x1_ASAP7_75t_L g804 ( 
.A(n_698),
.B(n_699),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_674),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_639),
.B(n_663),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_700),
.A2(n_702),
.B(n_718),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_710),
.A2(n_645),
.B(n_679),
.C(n_654),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_654),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_593),
.B(n_649),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_621),
.B(n_650),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_708),
.A2(n_709),
.B(n_717),
.C(n_711),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_714),
.A2(n_601),
.B(n_590),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_653),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_706),
.B(n_633),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_587),
.B(n_632),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_714),
.A2(n_601),
.B(n_590),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_713),
.A2(n_637),
.B(n_634),
.Y(n_820)
);

INVx11_ASAP7_75t_L g821 ( 
.A(n_695),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_641),
.A2(n_615),
.B1(n_703),
.B2(n_706),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_641),
.A2(n_615),
.B1(n_703),
.B2(n_706),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_653),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_714),
.A2(n_601),
.B(n_590),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_606),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_688),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_591),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_632),
.A2(n_667),
.B1(n_641),
.B2(n_611),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_591),
.Y(n_835)
);

OAI321xp33_ASAP7_75t_L g836 ( 
.A1(n_686),
.A2(n_452),
.A3(n_331),
.B1(n_346),
.B2(n_632),
.C(n_488),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_653),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_606),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_839)
);

BUFx4f_ASAP7_75t_L g840 ( 
.A(n_695),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_SL g841 ( 
.A(n_708),
.B(n_509),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_587),
.B(n_632),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_695),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_706),
.B(n_633),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_586),
.B(n_457),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_653),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_706),
.B(n_531),
.Y(n_849)
);

NOR2x1p5_ASAP7_75t_SL g850 ( 
.A(n_592),
.B(n_486),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_638),
.A2(n_561),
.B(n_655),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_833),
.A2(n_812),
.B(n_736),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_720),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_729),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_737),
.A2(n_793),
.B(n_734),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_813),
.A2(n_827),
.B(n_819),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_847),
.B(n_789),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_742),
.A2(n_788),
.B(n_787),
.Y(n_858)
);

OAI21xp33_ASAP7_75t_L g859 ( 
.A1(n_741),
.A2(n_738),
.B(n_816),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_752),
.A2(n_760),
.B(n_757),
.Y(n_860)
);

INVx4_ASAP7_75t_SL g861 ( 
.A(n_720),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_837),
.Y(n_862)
);

AOI221xp5_ASAP7_75t_SL g863 ( 
.A1(n_822),
.A2(n_823),
.B1(n_755),
.B2(n_774),
.C(n_795),
.Y(n_863)
);

AO221x2_ASAP7_75t_L g864 ( 
.A1(n_780),
.A2(n_744),
.B1(n_836),
.B2(n_754),
.C(n_723),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_814),
.Y(n_865)
);

AND2x6_ASAP7_75t_L g866 ( 
.A(n_804),
.B(n_798),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_SL g867 ( 
.A1(n_741),
.A2(n_738),
.B1(n_816),
.B2(n_842),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_745),
.B(n_773),
.Y(n_868)
);

OAI22x1_ASAP7_75t_L g869 ( 
.A1(n_842),
.A2(n_753),
.B1(n_735),
.B2(n_764),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_825),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_755),
.B(n_794),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_794),
.B(n_849),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_749),
.B(n_773),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_766),
.B(n_728),
.Y(n_874)
);

AO31x2_ASAP7_75t_L g875 ( 
.A1(n_807),
.A2(n_851),
.A3(n_846),
.B(n_844),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_753),
.A2(n_796),
.B(n_799),
.C(n_735),
.Y(n_876)
);

AOI21x1_ASAP7_75t_SL g877 ( 
.A1(n_725),
.A2(n_800),
.B(n_782),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_727),
.B(n_726),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_727),
.B(n_750),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_756),
.A2(n_839),
.B(n_834),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_727),
.B(n_721),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_824),
.A2(n_828),
.B(n_829),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_776),
.A2(n_739),
.B1(n_845),
.B2(n_815),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_777),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_765),
.A2(n_801),
.B(n_797),
.Y(n_886)
);

AOI21xp33_ASAP7_75t_L g887 ( 
.A1(n_746),
.A2(n_790),
.B(n_802),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_739),
.B(n_720),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_785),
.A2(n_770),
.B(n_778),
.Y(n_889)
);

BUFx8_ASAP7_75t_L g890 ( 
.A(n_759),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_832),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_832),
.B(n_786),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_837),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_767),
.A2(n_769),
.B(n_719),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_769),
.A2(n_724),
.B(n_790),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_841),
.A2(n_806),
.B(n_761),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_808),
.A2(n_802),
.B(n_805),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_796),
.A2(n_784),
.B(n_792),
.C(n_838),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_763),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_748),
.A2(n_783),
.B(n_768),
.C(n_830),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_733),
.B(n_792),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_791),
.A2(n_850),
.B(n_784),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_771),
.A2(n_764),
.B(n_803),
.C(n_747),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_732),
.B(n_832),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_835),
.B(n_832),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_732),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_805),
.A2(n_786),
.B(n_811),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_809),
.A2(n_779),
.B(n_805),
.Y(n_908)
);

NAND2x1_ASAP7_75t_L g909 ( 
.A(n_835),
.B(n_811),
.Y(n_909)
);

OAI21x1_ASAP7_75t_L g910 ( 
.A1(n_810),
.A2(n_754),
.B(n_740),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_848),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_740),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_751),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_754),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_754),
.Y(n_915)
);

AOI211x1_ASAP7_75t_L g916 ( 
.A1(n_758),
.A2(n_831),
.B(n_826),
.C(n_840),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_831),
.B(n_762),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_826),
.B(n_840),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_843),
.B(n_821),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_843),
.B(n_786),
.Y(n_920)
);

AO21x1_ASAP7_75t_L g921 ( 
.A1(n_833),
.A2(n_812),
.B(n_736),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_775),
.A2(n_638),
.B(n_496),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_847),
.B(n_833),
.Y(n_923)
);

AO31x2_ASAP7_75t_L g924 ( 
.A1(n_822),
.A2(n_823),
.A3(n_731),
.B(n_807),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_727),
.B(n_781),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_847),
.B(n_745),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_847),
.B(n_833),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_847),
.B(n_833),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_847),
.B(n_833),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_847),
.B(n_745),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_847),
.B(n_833),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_833),
.A2(n_741),
.B1(n_802),
.B2(n_769),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_833),
.B(n_738),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_751),
.Y(n_934)
);

INVx4_ASAP7_75t_SL g935 ( 
.A(n_720),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_814),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_775),
.A2(n_638),
.B(n_496),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_847),
.B(n_833),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_833),
.A2(n_738),
.B(n_741),
.C(n_772),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_727),
.B(n_781),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_809),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_777),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_775),
.A2(n_638),
.B(n_496),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_814),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_814),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_749),
.B(n_602),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_820),
.A2(n_743),
.B(n_730),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_833),
.B(n_738),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_727),
.B(n_781),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_847),
.B(n_833),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_813),
.A2(n_827),
.B(n_819),
.Y(n_951)
);

BUFx12f_ASAP7_75t_L g952 ( 
.A(n_814),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_833),
.A2(n_741),
.B1(n_802),
.B2(n_769),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_847),
.B(n_833),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_833),
.A2(n_812),
.B(n_736),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_817),
.A2(n_824),
.B(n_818),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_817),
.A2(n_824),
.B(n_818),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_775),
.A2(n_772),
.B(n_731),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_944),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_865),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_926),
.B(n_930),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_907),
.B(n_920),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_945),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_920),
.B(n_892),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_873),
.B(n_874),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_861),
.B(n_935),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_890),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_864),
.A2(n_932),
.B1(n_953),
.B2(n_869),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_857),
.B(n_874),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_953),
.A2(n_868),
.B1(n_955),
.B2(n_852),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_891),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_891),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_876),
.B(n_872),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_891),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_891),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_854),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_857),
.B(n_872),
.Y(n_977)
);

NOR2xp67_ASAP7_75t_L g978 ( 
.A(n_913),
.B(n_934),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_921),
.A2(n_950),
.B1(n_938),
.B2(n_931),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_854),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_923),
.B(n_927),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_856),
.A2(n_951),
.B1(n_923),
.B2(n_927),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_928),
.B(n_929),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_952),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_906),
.B(n_865),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_913),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_870),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_958),
.A2(n_943),
.B(n_937),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_854),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_928),
.B(n_929),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_871),
.B(n_912),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_941),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_936),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_SL g995 ( 
.A1(n_887),
.A2(n_898),
.B(n_903),
.C(n_954),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_L g996 ( 
.A(n_911),
.B(n_946),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_931),
.A2(n_938),
.B1(n_950),
.B2(n_915),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_887),
.A2(n_894),
.B(n_897),
.C(n_884),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_853),
.B(n_880),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_893),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_871),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_917),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_861),
.B(n_935),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_885),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_862),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_941),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_910),
.B(n_904),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_888),
.B(n_942),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_901),
.B(n_882),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_919),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_863),
.B(n_901),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_905),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_882),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_918),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_863),
.B(n_914),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_909),
.B(n_908),
.Y(n_1016)
);

INVx3_ASAP7_75t_SL g1017 ( 
.A(n_866),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_915),
.A2(n_895),
.B1(n_949),
.B2(n_940),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_915),
.B(n_878),
.Y(n_1019)
);

INVx6_ASAP7_75t_L g1020 ( 
.A(n_918),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_902),
.B(n_924),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_855),
.A2(n_883),
.B(n_879),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_905),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_879),
.A2(n_881),
.B(n_889),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_900),
.B(n_949),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_866),
.B(n_924),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_925),
.A2(n_940),
.B1(n_916),
.B2(n_896),
.Y(n_1027)
);

OR2x6_ASAP7_75t_SL g1028 ( 
.A(n_877),
.B(n_866),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_866),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_875),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_886),
.B(n_947),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_875),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_957),
.A2(n_867),
.B1(n_953),
.B2(n_932),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_956),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_860),
.B(n_859),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_853),
.Y(n_1036)
);

OAI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_867),
.A2(n_859),
.B(n_741),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_933),
.A2(n_948),
.B1(n_859),
.B2(n_867),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_859),
.B(n_741),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_933),
.A2(n_948),
.B1(n_859),
.B2(n_867),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_907),
.B(n_920),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_944),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_944),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_L g1044 ( 
.A(n_913),
.B(n_934),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_859),
.B(n_933),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_891),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_958),
.A2(n_775),
.B(n_922),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_958),
.A2(n_775),
.B(n_922),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_944),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_907),
.B(n_920),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_944),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_934),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_873),
.B(n_874),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_920),
.B(n_786),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_873),
.B(n_874),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_890),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_859),
.B(n_933),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_L g1058 ( 
.A(n_867),
.B(n_741),
.C(n_632),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_859),
.B(n_741),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_944),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_958),
.A2(n_775),
.B(n_922),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_899),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_859),
.A2(n_741),
.B(n_948),
.C(n_933),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_920),
.B(n_786),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_859),
.B(n_933),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_926),
.B(n_930),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_926),
.B(n_930),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_858),
.A2(n_741),
.B(n_738),
.C(n_632),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_939),
.A2(n_833),
.B(n_741),
.C(n_738),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_920),
.B(n_786),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_865),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_926),
.B(n_930),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1019),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1047),
.A2(n_1061),
.B(n_1048),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_1052),
.Y(n_1075)
);

BUFx2_ASAP7_75t_R g1076 ( 
.A(n_984),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_973),
.B(n_1038),
.Y(n_1077)
);

INVx6_ASAP7_75t_L g1078 ( 
.A(n_971),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_967),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_962),
.B(n_1041),
.Y(n_1080)
);

BUFx8_ASAP7_75t_L g1081 ( 
.A(n_985),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1062),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1022),
.A2(n_1024),
.B(n_989),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1039),
.B(n_1066),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1058),
.A2(n_1037),
.B1(n_1040),
.B2(n_1038),
.Y(n_1085)
);

INVx11_ASAP7_75t_L g1086 ( 
.A(n_1056),
.Y(n_1086)
);

AO21x1_ASAP7_75t_SL g1087 ( 
.A1(n_1026),
.A2(n_968),
.B(n_1040),
.Y(n_1087)
);

CKINVDCx10_ASAP7_75t_R g1088 ( 
.A(n_962),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_988),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_1042),
.Y(n_1090)
);

INVx3_ASAP7_75t_SL g1091 ( 
.A(n_987),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_972),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_976),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1007),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1019),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1069),
.A2(n_1063),
.B(n_1068),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1030),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_993),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1071),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1035),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_960),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1045),
.A2(n_1057),
.B1(n_1065),
.B2(n_1033),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1001),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1004),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_994),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1045),
.A2(n_1065),
.B1(n_1057),
.B2(n_1059),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1008),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_960),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_961),
.A2(n_1014),
.B1(n_1072),
.B2(n_1067),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_972),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_992),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_977),
.A2(n_969),
.B1(n_991),
.B2(n_983),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_986),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_997),
.B(n_982),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_965),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1053),
.Y(n_1116)
);

AO21x1_ASAP7_75t_SL g1117 ( 
.A1(n_1026),
.A2(n_979),
.B(n_970),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1055),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_981),
.A2(n_983),
.B1(n_997),
.B2(n_982),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_974),
.Y(n_1120)
);

BUFx2_ASAP7_75t_R g1121 ( 
.A(n_1049),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_998),
.A2(n_1015),
.B(n_1034),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1013),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_R g1124 ( 
.A1(n_1005),
.A2(n_1009),
.B1(n_1043),
.B2(n_995),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1000),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_969),
.B(n_981),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_996),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1015),
.Y(n_1128)
);

CKINVDCx11_ASAP7_75t_R g1129 ( 
.A(n_993),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1031),
.A2(n_1027),
.B(n_1018),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1002),
.A2(n_1020),
.B1(n_976),
.B2(n_1041),
.Y(n_1131)
);

OA21x2_ASAP7_75t_L g1132 ( 
.A1(n_1011),
.A2(n_1021),
.B(n_1025),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1020),
.A2(n_976),
.B1(n_1050),
.B2(n_964),
.Y(n_1133)
);

BUFx2_ASAP7_75t_SL g1134 ( 
.A(n_966),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1012),
.Y(n_1135)
);

OAI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1050),
.A2(n_1044),
.B1(n_978),
.B2(n_993),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1028),
.Y(n_1137)
);

INVxp67_ASAP7_75t_SL g1138 ( 
.A(n_975),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1054),
.B(n_1064),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_1010),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1054),
.A2(n_1070),
.B1(n_1064),
.B2(n_959),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_975),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1060),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1051),
.Y(n_1144)
);

CKINVDCx11_ASAP7_75t_R g1145 ( 
.A(n_963),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1023),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1006),
.A2(n_980),
.B1(n_990),
.B2(n_1017),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_1029),
.B(n_1016),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_980),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1070),
.B(n_966),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1029),
.B(n_1036),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_980),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1029),
.B(n_1036),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_SL g1154 ( 
.A1(n_990),
.A2(n_975),
.B1(n_1046),
.B2(n_1003),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1046),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_999),
.A2(n_1003),
.B(n_990),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1071),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_973),
.B(n_1038),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_988),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1058),
.A2(n_741),
.B1(n_948),
.B2(n_933),
.Y(n_1160)
);

BUFx2_ASAP7_75t_R g1161 ( 
.A(n_1052),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1029),
.B(n_973),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1058),
.A2(n_741),
.B1(n_948),
.B2(n_933),
.Y(n_1163)
);

BUFx2_ASAP7_75t_R g1164 ( 
.A(n_1052),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1029),
.B(n_973),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_973),
.B(n_1038),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1032),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1042),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1032),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_967),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_SL g1171 ( 
.A(n_1161),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1094),
.B(n_1132),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1094),
.B(n_1132),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1126),
.B(n_1073),
.Y(n_1174)
);

BUFx2_ASAP7_75t_SL g1175 ( 
.A(n_1093),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1162),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_1159),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1080),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1080),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1167),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1169),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1132),
.B(n_1100),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1162),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1080),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1101),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1097),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1074),
.A2(n_1083),
.B(n_1096),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1165),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1085),
.A2(n_1112),
.B(n_1114),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1122),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1122),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1165),
.B(n_1130),
.Y(n_1193)
);

BUFx2_ASAP7_75t_SL g1194 ( 
.A(n_1093),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1073),
.B(n_1095),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1077),
.B(n_1158),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1158),
.B(n_1166),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1084),
.B(n_1113),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1114),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1166),
.B(n_1087),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1087),
.B(n_1095),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1127),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1148),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1137),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1088),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1119),
.A2(n_1102),
.B(n_1133),
.Y(n_1206)
);

AOI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1131),
.A2(n_1151),
.B(n_1153),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1106),
.B(n_1128),
.Y(n_1208)
);

NOR2x1_ASAP7_75t_SL g1209 ( 
.A(n_1117),
.B(n_1128),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1117),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1099),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1151),
.B(n_1153),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1134),
.B(n_1156),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1123),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1103),
.B(n_1115),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1116),
.B(n_1118),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1104),
.A2(n_1137),
.B(n_1107),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1111),
.B(n_1082),
.Y(n_1218)
);

INVx4_ASAP7_75t_SL g1219 ( 
.A(n_1078),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1172),
.B(n_1157),
.Y(n_1220)
);

OAI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1190),
.A2(n_1109),
.B1(n_1198),
.B2(n_1141),
.C(n_1208),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1172),
.B(n_1108),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1172),
.B(n_1135),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1202),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1173),
.B(n_1146),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1173),
.B(n_1105),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1173),
.B(n_1155),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1182),
.B(n_1155),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1182),
.B(n_1180),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1182),
.B(n_1152),
.Y(n_1230)
);

OAI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1208),
.A2(n_1143),
.B1(n_1154),
.B2(n_1125),
.C(n_1147),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1177),
.B(n_1089),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1181),
.Y(n_1233)
);

OAI221xp5_ASAP7_75t_L g1234 ( 
.A1(n_1185),
.A2(n_1091),
.B1(n_1144),
.B2(n_1124),
.C(n_1089),
.Y(n_1234)
);

INVx5_ASAP7_75t_L g1235 ( 
.A(n_1193),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1171),
.A2(n_1124),
.B1(n_1149),
.B2(n_1121),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1195),
.B(n_1090),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1174),
.B(n_1136),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1174),
.B(n_1199),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1171),
.B(n_1091),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1202),
.Y(n_1241)
);

NOR2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1210),
.B(n_1079),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1199),
.B(n_1138),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_1193),
.B(n_1134),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1195),
.B(n_1092),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1214),
.B(n_1092),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1186),
.B(n_1149),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1186),
.B(n_1168),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1193),
.B(n_1078),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1204),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1217),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1191),
.B(n_1110),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1217),
.Y(n_1253)
);

OAI221xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1234),
.A2(n_1200),
.B1(n_1213),
.B2(n_1193),
.C(n_1185),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1236),
.B(n_1221),
.C(n_1234),
.Y(n_1255)
);

NOR3xp33_ASAP7_75t_L g1256 ( 
.A(n_1236),
.B(n_1207),
.C(n_1206),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1229),
.B(n_1196),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1245),
.B(n_1211),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1229),
.B(n_1196),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1233),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1221),
.A2(n_1210),
.B1(n_1205),
.B2(n_1213),
.Y(n_1261)
);

NOR3xp33_ASAP7_75t_L g1262 ( 
.A(n_1231),
.B(n_1207),
.C(n_1206),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1229),
.B(n_1196),
.Y(n_1263)
);

NAND4xp25_ASAP7_75t_L g1264 ( 
.A(n_1238),
.B(n_1216),
.C(n_1215),
.D(n_1218),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1238),
.B(n_1210),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1231),
.A2(n_1210),
.B1(n_1242),
.B2(n_1205),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1251),
.B(n_1187),
.C(n_1201),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1242),
.A2(n_1209),
.B(n_1210),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1239),
.A2(n_1189),
.B1(n_1197),
.B2(n_1215),
.C(n_1243),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1233),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1220),
.B(n_1197),
.Y(n_1271)
);

NOR3xp33_ASAP7_75t_L g1272 ( 
.A(n_1237),
.B(n_1206),
.C(n_1203),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1251),
.B(n_1187),
.C(n_1201),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1253),
.B(n_1187),
.C(n_1201),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1227),
.B(n_1197),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1220),
.B(n_1189),
.Y(n_1276)
);

AND2x2_ASAP7_75t_SL g1277 ( 
.A(n_1250),
.B(n_1210),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1227),
.B(n_1200),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1220),
.B(n_1178),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1222),
.B(n_1178),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1222),
.B(n_1178),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1222),
.B(n_1179),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1239),
.B(n_1179),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1253),
.B(n_1237),
.C(n_1243),
.Y(n_1284)
);

OAI221xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1247),
.A2(n_1200),
.B1(n_1213),
.B2(n_1193),
.C(n_1216),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1230),
.B(n_1184),
.Y(n_1286)
);

OA211x2_ASAP7_75t_L g1287 ( 
.A1(n_1240),
.A2(n_1219),
.B(n_1175),
.C(n_1194),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1227),
.B(n_1193),
.Y(n_1288)
);

OAI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1232),
.A2(n_1205),
.B1(n_1213),
.B2(n_1210),
.C(n_1183),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1246),
.B(n_1187),
.C(n_1214),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1226),
.B(n_1184),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1228),
.B(n_1192),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1247),
.B(n_1075),
.Y(n_1293)
);

OAI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1224),
.A2(n_1213),
.B1(n_1176),
.B2(n_1188),
.C(n_1183),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1224),
.A2(n_1139),
.B(n_1150),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1233),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_1246),
.B(n_1187),
.C(n_1192),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1296),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1257),
.B(n_1235),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1259),
.B(n_1235),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1259),
.B(n_1235),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1263),
.B(n_1278),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1260),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1288),
.B(n_1235),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1260),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1263),
.B(n_1235),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1255),
.A2(n_1204),
.B1(n_1212),
.B2(n_1139),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1277),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1270),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1278),
.B(n_1275),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1270),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1275),
.B(n_1235),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1296),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1292),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1276),
.B(n_1223),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1292),
.Y(n_1316)
);

INVxp67_ASAP7_75t_SL g1317 ( 
.A(n_1284),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1288),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1271),
.B(n_1235),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1277),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1280),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1267),
.B(n_1244),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1281),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1282),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1268),
.B(n_1244),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1272),
.B(n_1228),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1291),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1283),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1279),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1297),
.B(n_1252),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1273),
.B(n_1252),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1290),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1321),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1298),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1309),
.Y(n_1335)
);

OAI33xp33_ASAP7_75t_L g1336 ( 
.A1(n_1332),
.A2(n_1258),
.A3(n_1264),
.B1(n_1265),
.B2(n_1248),
.B3(n_1266),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1298),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1309),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1308),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1303),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1303),
.Y(n_1341)
);

NOR3x1_ASAP7_75t_L g1342 ( 
.A(n_1320),
.B(n_1289),
.C(n_1294),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1331),
.B(n_1286),
.Y(n_1343)
);

NOR2x1_ASAP7_75t_SL g1344 ( 
.A(n_1308),
.B(n_1244),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1299),
.B(n_1244),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1303),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1328),
.B(n_1269),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1305),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1298),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1308),
.A2(n_1256),
.B1(n_1262),
.B2(n_1261),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1328),
.B(n_1265),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1305),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1308),
.B(n_1241),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1331),
.B(n_1274),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1305),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1311),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1304),
.B(n_1244),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1332),
.B(n_1254),
.C(n_1285),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1311),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1328),
.B(n_1225),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1304),
.B(n_1249),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1299),
.B(n_1249),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1299),
.B(n_1249),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1311),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1314),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1314),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1313),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1331),
.B(n_1252),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1314),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1298),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1347),
.B(n_1317),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1354),
.B(n_1332),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1340),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1344),
.B(n_1302),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1334),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1339),
.B(n_1241),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1333),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1344),
.B(n_1339),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1358),
.A2(n_1317),
.B(n_1322),
.C(n_1320),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1354),
.B(n_1330),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1334),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1340),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1351),
.B(n_1321),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1343),
.B(n_1330),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1353),
.B(n_1302),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1336),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1342),
.B(n_1326),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1353),
.B(n_1302),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1350),
.B(n_1326),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1341),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1353),
.B(n_1362),
.Y(n_1391)
);

NAND2x1_ASAP7_75t_L g1392 ( 
.A(n_1357),
.B(n_1320),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1338),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1341),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1357),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1346),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1346),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1343),
.B(n_1326),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1368),
.B(n_1330),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1360),
.B(n_1327),
.Y(n_1401)
);

AOI322xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1345),
.A2(n_1316),
.A3(n_1310),
.B1(n_1312),
.B2(n_1300),
.C1(n_1301),
.C2(n_1306),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1337),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1348),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1368),
.B(n_1327),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1337),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1348),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1364),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1364),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1363),
.B(n_1327),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1338),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1345),
.B(n_1304),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1352),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1396),
.B(n_1357),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1376),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1396),
.B(n_1361),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1386),
.A2(n_1307),
.B1(n_1325),
.B2(n_1295),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1372),
.B(n_1335),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1392),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1372),
.B(n_1365),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1380),
.B(n_1366),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1371),
.B(n_1318),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1380),
.B(n_1399),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1376),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1374),
.B(n_1361),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1373),
.Y(n_1426)
);

CKINVDCx16_ASAP7_75t_R g1427 ( 
.A(n_1377),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1361),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1373),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1391),
.B(n_1310),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1392),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1379),
.A2(n_1307),
.B1(n_1325),
.B2(n_1322),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1376),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1393),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1384),
.B(n_1383),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1382),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1378),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1384),
.B(n_1369),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1378),
.B(n_1322),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1395),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1389),
.A2(n_1325),
.B1(n_1315),
.B2(n_1249),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1385),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1395),
.Y(n_1443)
);

AOI222xp33_ASAP7_75t_L g1444 ( 
.A1(n_1387),
.A2(n_1322),
.B1(n_1324),
.B2(n_1323),
.C1(n_1329),
.C2(n_1319),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1382),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1385),
.A2(n_1325),
.B1(n_1322),
.B2(n_1315),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1391),
.A2(n_1322),
.B1(n_1325),
.B2(n_1388),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1410),
.B(n_1318),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1412),
.B(n_1310),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1432),
.A2(n_1402),
.B1(n_1388),
.B2(n_1413),
.C(n_1409),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1427),
.B(n_1411),
.Y(n_1451)
);

NAND2xp67_ASAP7_75t_L g1452 ( 
.A(n_1415),
.B(n_1412),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1434),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1427),
.A2(n_1417),
.B1(n_1437),
.B2(n_1440),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1443),
.A2(n_1439),
.B1(n_1428),
.B2(n_1425),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1426),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1418),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1430),
.B(n_1449),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1444),
.A2(n_1447),
.B(n_1441),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1435),
.B(n_1170),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1442),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1435),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1430),
.B(n_1401),
.Y(n_1463)
);

AOI31xp33_ASAP7_75t_L g1464 ( 
.A1(n_1419),
.A2(n_1164),
.A3(n_1402),
.B(n_1400),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1442),
.Y(n_1465)
);

AOI222xp33_ASAP7_75t_L g1466 ( 
.A1(n_1422),
.A2(n_1405),
.B1(n_1413),
.B2(n_1293),
.C1(n_1408),
.C2(n_1404),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1419),
.A2(n_1400),
.B(n_1394),
.Y(n_1467)
);

AOI211xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1446),
.A2(n_1268),
.B(n_1408),
.C(n_1390),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1423),
.Y(n_1469)
);

NAND2xp67_ASAP7_75t_L g1470 ( 
.A(n_1415),
.B(n_1375),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1423),
.B(n_1170),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1449),
.B(n_1318),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1418),
.B(n_1390),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1425),
.B(n_1394),
.Y(n_1474)
);

NAND2x1_ASAP7_75t_L g1475 ( 
.A(n_1461),
.B(n_1431),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1457),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1448),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1457),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1462),
.B(n_1416),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1456),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1453),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1469),
.B(n_1416),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1458),
.B(n_1421),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1454),
.B(n_1414),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1473),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1461),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1471),
.B(n_1414),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1471),
.B(n_1428),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1465),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1450),
.B(n_1474),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1463),
.B(n_1421),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1464),
.A2(n_1459),
.B1(n_1455),
.B2(n_1460),
.Y(n_1493)
);

OAI211xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1491),
.A2(n_1476),
.B(n_1489),
.C(n_1488),
.Y(n_1494)
);

AOI21xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1491),
.A2(n_1466),
.B(n_1431),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1493),
.A2(n_1467),
.B1(n_1465),
.B2(n_1474),
.C(n_1429),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1493),
.A2(n_1439),
.B1(n_1433),
.B2(n_1424),
.Y(n_1497)
);

AOI211xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1477),
.A2(n_1439),
.B(n_1426),
.C(n_1436),
.Y(n_1498)
);

OAI32xp33_ASAP7_75t_L g1499 ( 
.A1(n_1485),
.A2(n_1424),
.A3(n_1433),
.B1(n_1468),
.B2(n_1420),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1480),
.A2(n_1439),
.B1(n_1472),
.B2(n_1420),
.Y(n_1500)
);

AOI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1482),
.A2(n_1429),
.B1(n_1445),
.B2(n_1436),
.C(n_1438),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1483),
.A2(n_1445),
.B(n_1438),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1486),
.B(n_1452),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1475),
.A2(n_1479),
.B(n_1478),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1494),
.B(n_1487),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1503),
.Y(n_1506)
);

NOR4xp25_ASAP7_75t_L g1507 ( 
.A(n_1496),
.B(n_1490),
.C(n_1481),
.D(n_1484),
.Y(n_1507)
);

NOR3xp33_ASAP7_75t_SL g1508 ( 
.A(n_1499),
.B(n_1492),
.C(n_1081),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1509)
);

NOR2x1_ASAP7_75t_L g1510 ( 
.A(n_1504),
.B(n_1159),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1498),
.B(n_1409),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1500),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1497),
.B(n_1145),
.C(n_1129),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1502),
.B(n_1168),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_SL g1515 ( 
.A(n_1507),
.B(n_1501),
.C(n_1140),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1511),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1505),
.A2(n_1398),
.B(n_1397),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1506),
.Y(n_1518)
);

NOR3xp33_ASAP7_75t_L g1519 ( 
.A(n_1510),
.B(n_1145),
.C(n_1129),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1518),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1515),
.A2(n_1513),
.B1(n_1512),
.B2(n_1509),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1519),
.B(n_1514),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1516),
.A2(n_1508),
.B1(n_1079),
.B2(n_1407),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1517),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1515),
.A2(n_1407),
.B1(n_1404),
.B2(n_1397),
.Y(n_1525)
);

OAI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1521),
.A2(n_1381),
.B1(n_1403),
.B2(n_1398),
.C(n_1406),
.Y(n_1526)
);

XNOR2x1_ASAP7_75t_L g1527 ( 
.A(n_1523),
.B(n_1081),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1520),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1524),
.B(n_1375),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1522),
.B(n_1075),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_L g1531 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1527),
.B(n_1081),
.Y(n_1532)
);

NOR3xp33_ASAP7_75t_L g1533 ( 
.A(n_1529),
.B(n_1525),
.C(n_1086),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1531),
.Y(n_1534)
);

NAND4xp25_ASAP7_75t_SL g1535 ( 
.A(n_1534),
.B(n_1533),
.C(n_1526),
.D(n_1532),
.Y(n_1535)
);

OA22x2_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_1381),
.B1(n_1403),
.B2(n_1406),
.Y(n_1536)
);

AO21x2_ASAP7_75t_L g1537 ( 
.A1(n_1535),
.A2(n_1403),
.B(n_1381),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1536),
.A2(n_1086),
.B1(n_1076),
.B2(n_1140),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1537),
.A2(n_1355),
.B1(n_1356),
.B2(n_1359),
.C(n_1367),
.Y(n_1539)
);

XOR2xp5_ASAP7_75t_L g1540 ( 
.A(n_1538),
.B(n_1075),
.Y(n_1540)
);

XNOR2xp5_ASAP7_75t_L g1541 ( 
.A(n_1539),
.B(n_1287),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1540),
.Y(n_1542)
);

AOI222xp33_ASAP7_75t_L g1543 ( 
.A1(n_1542),
.A2(n_1541),
.B1(n_1367),
.B2(n_1349),
.C1(n_1370),
.C2(n_1098),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_R g1544 ( 
.A1(n_1543),
.A2(n_1287),
.B1(n_1098),
.B2(n_1370),
.C(n_1349),
.Y(n_1544)
);

AOI211xp5_ASAP7_75t_L g1545 ( 
.A1(n_1544),
.A2(n_1142),
.B(n_1120),
.C(n_1110),
.Y(n_1545)
);


endmodule