module real_jpeg_18451_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_0),
.B(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

OR2x4_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_19),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_3),
.B(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_3),
.B(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_4),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_14),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NAND4xp25_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_25),
.C(n_36),
.D(n_41),
.Y(n_6)
);

AOI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_18),
.B(n_21),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_9),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g11 ( 
.A1(n_12),
.A2(n_15),
.B(n_16),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_31),
.B(n_33),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_17),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_25)
);

AND2x4_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

OR2x4_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_44),
.B(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);


endmodule