module fake_jpeg_23710_n_45 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_1),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_10),
.B1(n_20),
.B2(n_19),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.C(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_36),
.B1(n_34),
.B2(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_24),
.B1(n_13),
.B2(n_6),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_3),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_33),
.C(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B1(n_38),
.B2(n_25),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_44)
);

AOI221xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_45)
);


endmodule