module fake_jpeg_15652_n_354 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_354);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_45),
.Y(n_64)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_20),
.Y(n_75)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_45),
.B1(n_30),
.B2(n_34),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_43),
.B1(n_55),
.B2(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_77),
.A2(n_95),
.B1(n_48),
.B2(n_51),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_55),
.B1(n_54),
.B2(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_48),
.B1(n_51),
.B2(n_56),
.Y(n_131)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_97),
.Y(n_115)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_55),
.B1(n_53),
.B2(n_42),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_50),
.B1(n_44),
.B2(n_48),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_112),
.B1(n_113),
.B2(n_44),
.Y(n_124)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_68),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_64),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_114),
.Y(n_139)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_69),
.C(n_59),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_127),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_84),
.A2(n_42),
.B1(n_34),
.B2(n_33),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_80),
.C(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_112),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_137),
.B1(n_145),
.B2(n_85),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_25),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_143),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_32),
.B1(n_28),
.B2(n_35),
.Y(n_145)
);

INVxp67_ASAP7_75t_R g147 ( 
.A(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_52),
.B1(n_87),
.B2(n_90),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_131),
.C(n_51),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_74),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_157),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_78),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_115),
.B(n_28),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_32),
.Y(n_175)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_91),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_127),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_168),
.B1(n_170),
.B2(n_141),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_82),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_83),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_51),
.B1(n_49),
.B2(n_24),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_79),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_175),
.B(n_27),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_195),
.C(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_116),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_41),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_181),
.Y(n_218)
);

NAND2x1_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_134),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_188),
.B(n_197),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_119),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_139),
.C(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_139),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_143),
.B(n_142),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_169),
.B1(n_168),
.B2(n_149),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_140),
.A3(n_31),
.B1(n_21),
.B2(n_40),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_188),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_141),
.B(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_170),
.B(n_166),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_162),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_230),
.C(n_231),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_210),
.B1(n_180),
.B2(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_213),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_200),
.B1(n_181),
.B2(n_183),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_160),
.B1(n_123),
.B2(n_125),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_125),
.B1(n_136),
.B2(n_153),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_215),
.B1(n_193),
.B2(n_194),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_184),
.Y(n_213)
);

FAx1_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_117),
.CI(n_135),
.CON(n_214),
.SN(n_214)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_216),
.B(n_197),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_173),
.B1(n_123),
.B2(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_156),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_27),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_41),
.Y(n_226)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_41),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_175),
.B(n_21),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_174),
.C(n_187),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_47),
.C(n_46),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_47),
.C(n_46),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_29),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_235),
.A2(n_209),
.B1(n_232),
.B2(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_219),
.B(n_214),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_212),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_193),
.B(n_174),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_249),
.B1(n_250),
.B2(n_255),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_194),
.C(n_198),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_252),
.C(n_257),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_187),
.B(n_192),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_220),
.B1(n_203),
.B2(n_205),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_199),
.C(n_182),
.Y(n_252)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_199),
.B1(n_182),
.B2(n_152),
.Y(n_256)
);

AO22x1_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_29),
.B1(n_26),
.B2(n_39),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_183),
.C(n_135),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_240),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_264),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_274),
.B1(n_275),
.B2(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_207),
.Y(n_267)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_233),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_273),
.B(n_236),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_203),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_276),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_233),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_246),
.A2(n_219),
.B1(n_226),
.B2(n_230),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_29),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_29),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.Y(n_288)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_258),
.B1(n_247),
.B2(n_234),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_257),
.B1(n_258),
.B2(n_241),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_286),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_249),
.B1(n_244),
.B2(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_292),
.C(n_297),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_256),
.B1(n_250),
.B2(n_237),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_243),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_26),
.C(n_254),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_299),
.C(n_291),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_263),
.B(n_26),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_26),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_17),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_299),
.C(n_296),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_1),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_302),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_260),
.A3(n_265),
.B1(n_272),
.B2(n_266),
.C1(n_278),
.C2(n_276),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_304),
.A2(n_313),
.B(n_5),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_321)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_274),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_6),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_312),
.C(n_36),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_262),
.C(n_275),
.Y(n_312)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_285),
.A2(n_275),
.B(n_36),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_318),
.C(n_323),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_294),
.B1(n_297),
.B2(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_325),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_25),
.B1(n_23),
.B2(n_33),
.Y(n_319)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_301),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_318),
.B(n_316),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_23),
.B1(n_16),
.B2(n_8),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_6),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_311),
.A2(n_306),
.B1(n_312),
.B2(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_6),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_328),
.B(n_332),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_324),
.B1(n_315),
.B2(n_9),
.Y(n_337)
);

FAx1_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_309),
.CI(n_7),
.CON(n_332),
.SN(n_332)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_335),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_7),
.C(n_10),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_338),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_332),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_340),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_15),
.B(n_11),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_10),
.Y(n_342)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_330),
.A3(n_329),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_11),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g347 ( 
.A1(n_343),
.A2(n_337),
.B(n_341),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_15),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_346),
.B(n_10),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_349),
.B(n_344),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_345),
.B1(n_348),
.B2(n_14),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_11),
.B(n_12),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_352),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_353),
.B(n_12),
.Y(n_354)
);


endmodule