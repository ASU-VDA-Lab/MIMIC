module fake_jpeg_8678_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_16),
.B1(n_24),
.B2(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_16),
.B1(n_15),
.B2(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_45),
.B1(n_24),
.B2(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_63),
.B1(n_12),
.B2(n_17),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_33),
.B(n_34),
.C(n_32),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_64),
.Y(n_77)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_14),
.B1(n_25),
.B2(n_23),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_2),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_2),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_48),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_R g68 ( 
.A(n_62),
.B(n_58),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_52),
.B(n_64),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_65),
.B(n_23),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_55),
.C(n_57),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_86),
.C(n_77),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_70),
.C(n_84),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_88),
.C(n_80),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_101),
.C(n_91),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_68),
.B1(n_77),
.B2(n_81),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.C(n_105),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_91),
.A3(n_90),
.B1(n_70),
.B2(n_89),
.C1(n_60),
.C2(n_61),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_72),
.A3(n_21),
.B1(n_20),
.B2(n_51),
.C1(n_34),
.C2(n_37),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_7),
.B(n_8),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_108),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_21),
.C(n_20),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_106),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_37),
.B(n_46),
.C(n_11),
.D(n_8),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_51),
.B(n_7),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_112),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_3),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_59),
.Y(n_115)
);


endmodule