module fake_jpeg_6967_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_21),
.B1(n_32),
.B2(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_58),
.B1(n_18),
.B2(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_21),
.B1(n_17),
.B2(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_37),
.B1(n_26),
.B2(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_40),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_57),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_60),
.B1(n_57),
.B2(n_51),
.Y(n_107)
);

NAND2x1_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_41),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_70),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_47),
.B1(n_59),
.B2(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_72),
.B1(n_38),
.B2(n_39),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_80),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_35),
.B1(n_39),
.B2(n_30),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_85),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_35),
.C(n_33),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_56),
.C(n_19),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_35),
.B(n_1),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_28),
.B(n_35),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_19),
.B(n_25),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_0),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_38),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_63),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_25),
.C(n_24),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_109),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_53),
.B1(n_42),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_81),
.B1(n_67),
.B2(n_76),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_75),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_72),
.B1(n_66),
.B2(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_74),
.B1(n_75),
.B2(n_86),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_121),
.B1(n_126),
.B2(n_95),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_84),
.B(n_69),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_87),
.B(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_84),
.B1(n_69),
.B2(n_23),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_127),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_31),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_92),
.B(n_8),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_130),
.B1(n_134),
.B2(n_6),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_23),
.B1(n_51),
.B2(n_24),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_25),
.C(n_2),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_93),
.B1(n_98),
.B2(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_4),
.C(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_5),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_133),
.B(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_117),
.B(n_115),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_151),
.B1(n_157),
.B2(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_103),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_92),
.C(n_8),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_155),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_161),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_92),
.B(n_9),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_154),
.B(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_9),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_9),
.B(n_10),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_102),
.B1(n_96),
.B2(n_12),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_96),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_167),
.B1(n_152),
.B2(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_124),
.B1(n_130),
.B2(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_171),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_140),
.B(n_141),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_177),
.B(n_178),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_123),
.C(n_122),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_138),
.C(n_142),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_188),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_142),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_144),
.B1(n_154),
.B2(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_196),
.B1(n_202),
.B2(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_173),
.C(n_177),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_182),
.Y(n_194)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_155),
.B1(n_150),
.B2(n_145),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_190),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_170),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_201),
.B(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_156),
.B1(n_127),
.B2(n_153),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_199),
.B(n_172),
.C(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_209),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_172),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_178),
.C(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_221),
.C(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_184),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_189),
.B1(n_196),
.B2(n_191),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_227),
.B1(n_209),
.B2(n_203),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_174),
.B1(n_165),
.B2(n_176),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_235),
.B(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_227),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_210),
.C(n_208),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_219),
.B(n_217),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_208),
.C(n_211),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_225),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_242),
.B(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_229),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_216),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_198),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_233),
.A3(n_228),
.B1(n_216),
.B2(n_204),
.C1(n_165),
.C2(n_197),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_244),
.B(n_228),
.C(n_129),
.Y(n_252)
);

OAI31xp67_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_248),
.A3(n_11),
.B(n_12),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_251),
.B1(n_14),
.B2(n_15),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_10),
.Y(n_256)
);


endmodule