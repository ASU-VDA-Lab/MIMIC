module fake_netlist_1_12451_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NAND2xp33_ASAP7_75t_SL g3 ( .A(n_0), .B(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
NOR2xp33_ASAP7_75t_L g5 ( .A(n_4), .B(n_0), .Y(n_5) );
NOR2x1_ASAP7_75t_R g6 ( .A(n_5), .B(n_4), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_0), .Y(n_7) );
OR2x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_3), .Y(n_8) );
NOR4xp75_ASAP7_75t_L g9 ( .A(n_8), .B(n_7), .C(n_1), .D(n_2), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_1), .Y(n_11) );
endmodule