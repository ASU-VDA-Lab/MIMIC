module fake_netlist_5_2313_n_1315 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1315);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1315;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1292;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_370;
wire n_976;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1309;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_1286;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_577;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_384;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_163),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_223),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_194),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_6),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_329),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_64),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_120),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_286),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_266),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_336),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_281),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_278),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_295),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_129),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_165),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_121),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_258),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_112),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_199),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_301),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_122),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_188),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_288),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_136),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_97),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_154),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_108),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_61),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_106),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_169),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_184),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_245),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_284),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_343),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_81),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_207),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_0),
.B(n_77),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_271),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_44),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_299),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_305),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_267),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_53),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_283),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_304),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_259),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_124),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_174),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_236),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_319),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_264),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_87),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_119),
.B(n_317),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_75),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_202),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_71),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_220),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_263),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_134),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_161),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_231),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_221),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_337),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_252),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_279),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_206),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_172),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_201),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_162),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_262),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_67),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_29),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_282),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_179),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_42),
.Y(n_423)
);

BUFx2_ASAP7_75t_SL g424 ( 
.A(n_212),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_224),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_18),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_100),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_190),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_38),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_101),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_62),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_138),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_67),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_34),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_46),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_155),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_33),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_254),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_18),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_92),
.Y(n_441)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_325),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_99),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_131),
.B(n_222),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_79),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_105),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_102),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_321),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_123),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_315),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_81),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_260),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_256),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_113),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_248),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_208),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_32),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_320),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_226),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_116),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_291),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_183),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_16),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_318),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_94),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_200),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_273),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_331),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_209),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_65),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_251),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_79),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_335),
.Y(n_473)
);

BUFx5_ASAP7_75t_L g474 ( 
.A(n_125),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_12),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_55),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_88),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_242),
.Y(n_478)
);

BUFx8_ASAP7_75t_SL g479 ( 
.A(n_130),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_211),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_227),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_98),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_287),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_180),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_232),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_17),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_68),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_14),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_310),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_244),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_268),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_170),
.Y(n_492)
);

BUFx5_ASAP7_75t_L g493 ( 
.A(n_225),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_285),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_322),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_217),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_93),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_3),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_141),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_139),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_41),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_0),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_358),
.Y(n_504)
);

BUFx8_ASAP7_75t_SL g505 ( 
.A(n_479),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_476),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_498),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_1),
.Y(n_509)
);

BUFx8_ASAP7_75t_SL g510 ( 
.A(n_423),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_358),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_1),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_463),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_395),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_361),
.A2(n_364),
.B(n_362),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_487),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

BUFx8_ASAP7_75t_SL g528 ( 
.A(n_426),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_347),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_351),
.B(n_4),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_354),
.B(n_5),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_383),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_489),
.B(n_5),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_393),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_7),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_350),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_410),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_386),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_402),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_413),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_419),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_352),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_375),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_433),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_349),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_422),
.B(n_8),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_449),
.B(n_8),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_453),
.A2(n_90),
.B(n_89),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_441),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

CKINVDCx6p67_ASAP7_75t_R g557 ( 
.A(n_391),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_451),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_462),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_480),
.B(n_9),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_501),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_442),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_382),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_470),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_390),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_403),
.Y(n_571)
);

OAI22x1_ASAP7_75t_SL g572 ( 
.A1(n_436),
.A2(n_475),
.B1(n_435),
.B2(n_438),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_353),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_491),
.B(n_10),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_365),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_366),
.A2(n_95),
.B(n_91),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_460),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_368),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_369),
.B(n_10),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_370),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_503),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_505),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_511),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_516),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_519),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_510),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_506),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_507),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_551),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_528),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_523),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_573),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_513),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_557),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_513),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_513),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_537),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_529),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_514),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_514),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_529),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_536),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_571),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_514),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_525),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_548),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_546),
.B(n_471),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_548),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_525),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_548),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_525),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_563),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_567),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_544),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_566),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_532),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_567),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_577),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_577),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_569),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_546),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_522),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_526),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_520),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_504),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_597),
.B(n_533),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_627),
.B(n_530),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_552),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_622),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_610),
.B(n_512),
.Y(n_637)
);

INVx8_ASAP7_75t_L g638 ( 
.A(n_596),
.Y(n_638)
);

BUFx5_ASAP7_75t_L g639 ( 
.A(n_591),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_594),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_588),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_603),
.B(n_518),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_626),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_598),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_608),
.B(n_518),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_614),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_601),
.B(n_518),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_588),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_604),
.B(n_502),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_380),
.B1(n_381),
.B2(n_348),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_632),
.B(n_555),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_589),
.B(n_531),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_588),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_587),
.B(n_531),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_607),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_592),
.B(n_521),
.C(n_553),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_619),
.B(n_585),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_593),
.B(n_535),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_602),
.B(n_502),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_606),
.B(n_550),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_631),
.B(n_445),
.C(n_568),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_595),
.B(n_535),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_612),
.B(n_509),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_595),
.B(n_509),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_609),
.B(n_611),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_628),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_582),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_581),
.A2(n_561),
.B1(n_574),
.B2(n_579),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_613),
.B(n_508),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_623),
.B(n_579),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_615),
.B(n_355),
.Y(n_672)
);

BUFx4_ASAP7_75t_L g673 ( 
.A(n_586),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_629),
.B(n_580),
.C(n_575),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_616),
.B(n_517),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_621),
.B(n_578),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_630),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_583),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_584),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_624),
.B(n_561),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_600),
.B(n_524),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_617),
.B(n_578),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_618),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_590),
.B(n_384),
.C(n_372),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_622),
.B(n_574),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_597),
.B(n_578),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_SL g688 ( 
.A(n_626),
.B(n_440),
.C(n_429),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_620),
.B(n_524),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_622),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_620),
.B(n_532),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_534),
.Y(n_692)
);

NAND2x1_ASAP7_75t_L g693 ( 
.A(n_588),
.B(n_374),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_627),
.B(n_405),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_SL g695 ( 
.A(n_651),
.B(n_407),
.C(n_406),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_636),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_633),
.B(n_409),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_661),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_689),
.A2(n_424),
.B1(n_377),
.B2(n_378),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_686),
.B(n_539),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_679),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_686),
.B(n_539),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_684),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_678),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_687),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_683),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_641),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_668),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_690),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_640),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_649),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_682),
.A2(n_576),
.B(n_554),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_686),
.B(n_539),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_665),
.A2(n_448),
.B1(n_454),
.B2(n_443),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_658),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_660),
.B(n_540),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_670),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_641),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_SL g719 ( 
.A(n_657),
.B(n_472),
.C(n_457),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_677),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_638),
.B(n_558),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_664),
.A2(n_545),
.B(n_527),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_667),
.B(n_644),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_647),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_655),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_663),
.A2(n_478),
.B1(n_447),
.B2(n_444),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_634),
.A2(n_357),
.B1(n_359),
.B2(n_356),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_638),
.B(n_558),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_SL g729 ( 
.A(n_659),
.B(n_408),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_653),
.B(n_572),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_671),
.B(n_656),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_654),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_680),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_SL g734 ( 
.A(n_694),
.B(n_488),
.C(n_363),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_669),
.B(n_540),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_681),
.B(n_538),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_688),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_639),
.B(n_547),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_692),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_675),
.A2(n_367),
.B1(n_371),
.B2(n_360),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_674),
.B(n_541),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_R g742 ( 
.A(n_666),
.B(n_373),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_639),
.B(n_547),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_693),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_652),
.B(n_376),
.Y(n_745)
);

CKINVDCx8_ASAP7_75t_R g746 ( 
.A(n_673),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_648),
.A2(n_400),
.B(n_450),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_645),
.B(n_559),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_662),
.B(n_543),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_676),
.B(n_379),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_637),
.A2(n_455),
.B1(n_456),
.B2(n_452),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_672),
.B(n_549),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_685),
.B(n_562),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_562),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_642),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_385),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_635),
.B(n_564),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_SL g758 ( 
.A1(n_651),
.A2(n_570),
.B1(n_388),
.B2(n_389),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_635),
.B(n_564),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_679),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_661),
.B(n_570),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_635),
.B(n_564),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_678),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_635),
.B(n_459),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_668),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_635),
.B(n_465),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_678),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_633),
.B(n_387),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_650),
.B(n_392),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_678),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_691),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_661),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_678),
.Y(n_773)
);

NOR2x1_ASAP7_75t_R g774 ( 
.A(n_668),
.B(n_394),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_633),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_650),
.B(n_404),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_635),
.B(n_483),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_661),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_635),
.B(n_490),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_678),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_668),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_668),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_697),
.A2(n_494),
.B1(n_495),
.B2(n_492),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_771),
.A2(n_497),
.B(n_496),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_768),
.B(n_499),
.Y(n_785)
);

O2A1O1Ixp5_ASAP7_75t_L g786 ( 
.A1(n_747),
.A2(n_500),
.B(n_560),
.C(n_556),
.Y(n_786)
);

OR2x6_ASAP7_75t_SL g787 ( 
.A(n_708),
.B(n_411),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_764),
.A2(n_565),
.B(n_412),
.C(n_414),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_696),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_SL g790 ( 
.A(n_765),
.B(n_415),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_782),
.Y(n_791)
);

OAI22x1_ASAP7_75t_L g792 ( 
.A1(n_730),
.A2(n_417),
.B1(n_418),
.B2(n_416),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_746),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_698),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_706),
.B(n_421),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_739),
.B(n_705),
.Y(n_796)
);

OAI22x1_ASAP7_75t_L g797 ( 
.A1(n_772),
.A2(n_778),
.B1(n_714),
.B2(n_715),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_731),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_725),
.B(n_428),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_726),
.A2(n_766),
.B(n_779),
.C(n_777),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_699),
.A2(n_437),
.B1(n_439),
.B2(n_430),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_733),
.A2(n_458),
.B1(n_466),
.B2(n_461),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_703),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_757),
.B(n_467),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_717),
.B(n_468),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_709),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_759),
.A2(n_473),
.B(n_469),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_SL g808 ( 
.A(n_718),
.B(n_477),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_710),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_762),
.A2(n_485),
.B(n_482),
.Y(n_810)
);

AO21x1_ASAP7_75t_L g811 ( 
.A1(n_700),
.A2(n_713),
.B(n_702),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_745),
.A2(n_493),
.B(n_474),
.C(n_12),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_SL g813 ( 
.A(n_775),
.B(n_493),
.C(n_474),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_781),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_736),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_753),
.B(n_721),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_753),
.B(n_11),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_720),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_736),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_723),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_755),
.A2(n_493),
.B(n_14),
.C(n_11),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_731),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_719),
.A2(n_16),
.B(n_13),
.C(n_15),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_723),
.B(n_96),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_721),
.B(n_728),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_704),
.A2(n_19),
.B(n_15),
.C(n_17),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_728),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_738),
.A2(n_748),
.B(n_743),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_758),
.B(n_19),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_769),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_752),
.B(n_103),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_756),
.B(n_104),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_749),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_SL g834 ( 
.A(n_718),
.B(n_20),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_741),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_776),
.B(n_21),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_716),
.B(n_22),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_774),
.B(n_23),
.Y(n_838)
);

OAI21x1_ASAP7_75t_L g839 ( 
.A1(n_744),
.A2(n_109),
.B(n_107),
.Y(n_839)
);

OA21x2_ASAP7_75t_L g840 ( 
.A1(n_722),
.A2(n_111),
.B(n_110),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_763),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_751),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_767),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_770),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_773),
.B(n_27),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_707),
.A2(n_115),
.B(n_114),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_727),
.B(n_28),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_780),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_734),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_718),
.A2(n_118),
.B(n_117),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_724),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_754),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_701),
.Y(n_853)
);

CKINVDCx10_ASAP7_75t_R g854 ( 
.A(n_737),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_741),
.A2(n_34),
.B(n_35),
.Y(n_856)
);

BUFx4f_ASAP7_75t_L g857 ( 
.A(n_754),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_740),
.B(n_35),
.Y(n_858)
);

BUFx12f_ASAP7_75t_L g859 ( 
.A(n_729),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_742),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_732),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_750),
.B(n_36),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_711),
.B(n_37),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_744),
.B(n_39),
.C(n_40),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_698),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_768),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_768),
.B(n_43),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_697),
.A2(n_127),
.B1(n_128),
.B2(n_126),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_698),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_771),
.A2(n_133),
.B(n_132),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_768),
.B(n_44),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_SL g872 ( 
.A(n_695),
.B(n_45),
.C(n_46),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_697),
.B(n_45),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_696),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_696),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_768),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_725),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_706),
.B(n_135),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_708),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_768),
.B(n_50),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_698),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_708),
.B(n_137),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_768),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_746),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_696),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_768),
.B(n_51),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_698),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_746),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_768),
.B(n_52),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_746),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_SL g891 ( 
.A(n_708),
.B(n_140),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_697),
.A2(n_143),
.B1(n_144),
.B2(n_142),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_771),
.A2(n_146),
.B(n_145),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_761),
.B(n_53),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_768),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_697),
.B(n_54),
.C(n_56),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_746),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_746),
.Y(n_898)
);

OAI21xp33_ASAP7_75t_SL g899 ( 
.A1(n_735),
.A2(n_57),
.B(n_58),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_SL g900 ( 
.A1(n_712),
.A2(n_148),
.B(n_149),
.C(n_147),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_746),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_L g902 ( 
.A1(n_697),
.A2(n_57),
.B(n_58),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_696),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_771),
.A2(n_151),
.B(n_150),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_SL g905 ( 
.A(n_697),
.B(n_59),
.C(n_60),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_747),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_696),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_800),
.A2(n_153),
.B(n_152),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_828),
.A2(n_157),
.B(n_156),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_814),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_811),
.A2(n_159),
.B(n_158),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_873),
.A2(n_858),
.B1(n_871),
.B2(n_867),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_798),
.B(n_160),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_869),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_833),
.B(n_63),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_839),
.A2(n_166),
.B(n_164),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_789),
.Y(n_917)
);

AO21x2_ASAP7_75t_L g918 ( 
.A1(n_813),
.A2(n_785),
.B(n_880),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_803),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_894),
.B(n_64),
.Y(n_920)
);

AO21x2_ASAP7_75t_L g921 ( 
.A1(n_886),
.A2(n_168),
.B(n_167),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_794),
.B(n_65),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_875),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_791),
.Y(n_924)
);

OR2x6_ASAP7_75t_SL g925 ( 
.A(n_879),
.B(n_66),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_819),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_870),
.A2(n_173),
.B(n_171),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_793),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_847),
.B(n_69),
.C(n_70),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_835),
.B(n_175),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_793),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_877),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_884),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_815),
.B(n_820),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_822),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_822),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_893),
.A2(n_177),
.B(n_176),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_874),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_885),
.Y(n_940)
);

OAI21x1_ASAP7_75t_SL g941 ( 
.A1(n_906),
.A2(n_830),
.B(n_904),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_824),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_903),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_907),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_809),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_825),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_786),
.A2(n_181),
.B(n_178),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_796),
.B(n_71),
.Y(n_948)
);

BUFx12f_ASAP7_75t_L g949 ( 
.A(n_884),
.Y(n_949)
);

AOI22x1_ASAP7_75t_L g950 ( 
.A1(n_792),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_889),
.A2(n_250),
.B1(n_345),
.B2(n_344),
.Y(n_951)
);

BUFx6f_ASAP7_75t_SL g952 ( 
.A(n_888),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_900),
.A2(n_185),
.B(n_182),
.Y(n_953)
);

BUFx12f_ASAP7_75t_L g954 ( 
.A(n_888),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_890),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_806),
.Y(n_956)
);

AO21x2_ASAP7_75t_L g957 ( 
.A1(n_837),
.A2(n_187),
.B(n_186),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_860),
.B(n_72),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_881),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_825),
.B(n_73),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_824),
.B(n_818),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_857),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_784),
.A2(n_191),
.B(n_189),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_812),
.A2(n_193),
.B(n_192),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_887),
.Y(n_965)
);

OAI21x1_ASAP7_75t_SL g966 ( 
.A1(n_842),
.A2(n_196),
.B(n_195),
.Y(n_966)
);

OA21x2_ASAP7_75t_L g967 ( 
.A1(n_863),
.A2(n_198),
.B(n_197),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_816),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_795),
.B(n_74),
.Y(n_969)
);

INVx4_ASAP7_75t_SL g970 ( 
.A(n_890),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_844),
.Y(n_971)
);

BUFx2_ASAP7_75t_SL g972 ( 
.A(n_882),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_848),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_851),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_862),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_975)
);

AO21x2_ASAP7_75t_L g976 ( 
.A1(n_804),
.A2(n_269),
.B(n_340),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_846),
.A2(n_265),
.B(n_339),
.Y(n_977)
);

AO21x1_ASAP7_75t_SL g978 ( 
.A1(n_866),
.A2(n_261),
.B(n_338),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_897),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_855),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_853),
.B(n_203),
.Y(n_981)
);

AO22x2_ASAP7_75t_L g982 ( 
.A1(n_905),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_799),
.B(n_82),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_861),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_845),
.Y(n_985)
);

OAI21x1_ASAP7_75t_SL g986 ( 
.A1(n_843),
.A2(n_272),
.B(n_334),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_827),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_821),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_898),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_788),
.A2(n_270),
.B(n_333),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_827),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_840),
.A2(n_257),
.B(n_332),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_805),
.B(n_83),
.Y(n_993)
);

AO21x2_ASAP7_75t_L g994 ( 
.A1(n_832),
.A2(n_255),
.B(n_330),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_856),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_901),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_840),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_859),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_817),
.B(n_204),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_850),
.A2(n_274),
.B(n_328),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_831),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_901),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_797),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_878),
.B(n_83),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_891),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_829),
.B(n_84),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_787),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_836),
.Y(n_1008)
);

AO21x2_ASAP7_75t_L g1009 ( 
.A1(n_807),
.A2(n_253),
.B(n_327),
.Y(n_1009)
);

AO21x2_ASAP7_75t_L g1010 ( 
.A1(n_810),
.A2(n_249),
.B(n_326),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_790),
.B(n_84),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_899),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_872),
.B(n_85),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_854),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_838),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_849),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_868),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_892),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_783),
.Y(n_1019)
);

OA21x2_ASAP7_75t_L g1020 ( 
.A1(n_876),
.A2(n_275),
.B(n_324),
.Y(n_1020)
);

NOR2x1_ASAP7_75t_R g1021 ( 
.A(n_834),
.B(n_85),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_802),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_808),
.Y(n_1023)
);

INVx5_ASAP7_75t_L g1024 ( 
.A(n_864),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_823),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_801),
.A2(n_247),
.B(n_316),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_902),
.B(n_86),
.Y(n_1027)
);

AO21x2_ASAP7_75t_L g1028 ( 
.A1(n_883),
.A2(n_246),
.B(n_314),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_895),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_896),
.B(n_205),
.Y(n_1030)
);

BUFx10_ASAP7_75t_L g1031 ( 
.A(n_826),
.Y(n_1031)
);

CKINVDCx8_ASAP7_75t_R g1032 ( 
.A(n_852),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_841),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_798),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_798),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1008),
.B(n_86),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_936),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_912),
.B(n_87),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_983),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_919),
.Y(n_1040)
);

OAI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_1032),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_917),
.Y(n_1042)
);

INVx8_ASAP7_75t_L g1043 ( 
.A(n_928),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_959),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_942),
.B(n_219),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_956),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_L g1047 ( 
.A(n_933),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_914),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_956),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_970),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_940),
.Y(n_1051)
);

INVxp33_ASAP7_75t_L g1052 ( 
.A(n_991),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_935),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_SL g1054 ( 
.A1(n_1006),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1015),
.B(n_346),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_965),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_952),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_943),
.Y(n_1058)
);

BUFx2_ASAP7_75t_R g1059 ( 
.A(n_931),
.Y(n_1059)
);

BUFx2_ASAP7_75t_R g1060 ( 
.A(n_955),
.Y(n_1060)
);

CKINVDCx11_ASAP7_75t_R g1061 ( 
.A(n_1014),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_932),
.Y(n_1062)
);

INVxp33_ASAP7_75t_L g1063 ( 
.A(n_984),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1004),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_968),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_926),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_SL g1067 ( 
.A1(n_1006),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_939),
.Y(n_1069)
);

AO21x1_ASAP7_75t_SL g1070 ( 
.A1(n_908),
.A2(n_240),
.B(n_241),
.Y(n_1070)
);

BUFx4f_ASAP7_75t_SL g1071 ( 
.A(n_949),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_971),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1013),
.B(n_243),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1004),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_1074)
);

INVx3_ASAP7_75t_SL g1075 ( 
.A(n_970),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_973),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_974),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_910),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_935),
.Y(n_1079)
);

NOR2x1_ASAP7_75t_R g1080 ( 
.A(n_954),
.B(n_289),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1029),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_979),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_923),
.Y(n_1083)
);

INVx8_ASAP7_75t_L g1084 ( 
.A(n_989),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_1005),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_997),
.A2(n_298),
.B(n_300),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_920),
.B(n_302),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_969),
.A2(n_303),
.B1(n_306),
.B2(n_307),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_988),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_SL g1090 ( 
.A1(n_1030),
.A2(n_308),
.B1(n_309),
.B2(n_311),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1017),
.A2(n_312),
.B1(n_313),
.B2(n_1018),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_985),
.A2(n_1001),
.B(n_1012),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_924),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_980),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1030),
.A2(n_1016),
.B1(n_993),
.B2(n_1025),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_987),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_980),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_935),
.Y(n_1098)
);

CKINVDCx11_ASAP7_75t_R g1099 ( 
.A(n_925),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_941),
.A2(n_992),
.B(n_990),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_948),
.B(n_999),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_999),
.B(n_1011),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_961),
.B(n_915),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_SL g1104 ( 
.A1(n_1025),
.A2(n_950),
.B1(n_1022),
.B2(n_929),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1001),
.A2(n_1012),
.B(n_995),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_909),
.A2(n_992),
.B(n_941),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_945),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_996),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1002),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1003),
.A2(n_995),
.B1(n_1019),
.B2(n_975),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_922),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_987),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1034),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_962),
.B(n_942),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1033),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_987),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_981),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_981),
.Y(n_1118)
);

AO21x1_ASAP7_75t_L g1119 ( 
.A1(n_951),
.A2(n_1026),
.B(n_938),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1034),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1027),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1020),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1031),
.A2(n_950),
.B1(n_1024),
.B2(n_978),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_934),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_934),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_916),
.A2(n_927),
.B(n_977),
.Y(n_1126)
);

INVx6_ASAP7_75t_L g1127 ( 
.A(n_946),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1035),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_1035),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_942),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_962),
.B(n_958),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_946),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1061),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1040),
.B(n_962),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_1108),
.B(n_1035),
.Y(n_1135)
);

OR2x2_ASAP7_75t_SL g1136 ( 
.A(n_1038),
.B(n_998),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1121),
.B(n_1024),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1076),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1057),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_1043),
.B(n_960),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1037),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1055),
.B(n_930),
.C(n_1007),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1044),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_1043),
.B(n_960),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1050),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1101),
.B(n_937),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1050),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1102),
.B(n_1103),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1036),
.B(n_982),
.C(n_1021),
.Y(n_1149)
);

NAND2xp33_ASAP7_75t_R g1150 ( 
.A(n_1131),
.B(n_967),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1073),
.B(n_982),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_1127),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1119),
.A2(n_953),
.A3(n_911),
.B(n_918),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1111),
.B(n_1023),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1095),
.B(n_1031),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1110),
.B(n_972),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1048),
.B(n_1023),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1056),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_1093),
.B(n_998),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1057),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1065),
.B(n_1023),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1062),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_R g1163 ( 
.A(n_1075),
.B(n_998),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1077),
.Y(n_1164)
);

AOI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1104),
.A2(n_966),
.B1(n_986),
.B2(n_964),
.C(n_1028),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1082),
.B(n_1109),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1087),
.B(n_913),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1096),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1122),
.A2(n_963),
.A3(n_947),
.B(n_921),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1063),
.B(n_994),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1122),
.A2(n_947),
.A3(n_1009),
.B(n_957),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1114),
.B(n_1009),
.C(n_976),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1069),
.B(n_1010),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1046),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1084),
.B(n_1000),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_1112),
.Y(n_1176)
);

BUFx10_ASAP7_75t_L g1177 ( 
.A(n_1127),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1066),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1049),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1123),
.B(n_1074),
.C(n_1064),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1117),
.A2(n_1118),
.B1(n_1092),
.B2(n_1115),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1084),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1051),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1058),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1072),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_R g1186 ( 
.A(n_1047),
.B(n_1071),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1047),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_SL g1188 ( 
.A(n_1041),
.B(n_1088),
.C(n_1130),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1132),
.B(n_1120),
.Y(n_1189)
);

NAND4xp25_ASAP7_75t_L g1190 ( 
.A(n_1124),
.B(n_1125),
.C(n_1107),
.D(n_1083),
.Y(n_1190)
);

CKINVDCx16_ASAP7_75t_R g1191 ( 
.A(n_1078),
.Y(n_1191)
);

NOR2x1p5_ASAP7_75t_L g1192 ( 
.A(n_1045),
.B(n_1079),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1116),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1042),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1099),
.Y(n_1195)
);

CKINVDCx8_ASAP7_75t_R g1196 ( 
.A(n_1053),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_R g1197 ( 
.A(n_1053),
.B(n_1098),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1068),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1105),
.B(n_1094),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1138),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1141),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1143),
.B(n_1097),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1180),
.A2(n_1090),
.B(n_1067),
.C(n_1054),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1151),
.B(n_1089),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1164),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1149),
.A2(n_1039),
.B1(n_1091),
.B2(n_1081),
.C(n_1052),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1194),
.B(n_1100),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1198),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1197),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1158),
.B(n_1059),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1174),
.B(n_1106),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1179),
.B(n_1070),
.Y(n_1213)
);

BUFx4f_ASAP7_75t_SL g1214 ( 
.A(n_1187),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1166),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1185),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1173),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1196),
.Y(n_1218)
);

INVx4_ASAP7_75t_R g1219 ( 
.A(n_1145),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1155),
.A2(n_1156),
.B1(n_1137),
.B2(n_1190),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1157),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1183),
.B(n_1184),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1152),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1148),
.B(n_1060),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1162),
.B(n_1128),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1168),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1181),
.B(n_1085),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1192),
.B(n_1086),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1146),
.B(n_1113),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1161),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1177),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1175),
.B(n_1126),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1170),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1233),
.B(n_1172),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1200),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1205),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1209),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1230),
.B(n_1154),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1203),
.B(n_1165),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1207),
.B(n_1153),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1201),
.B(n_1176),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1226),
.B(n_1167),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1207),
.B(n_1171),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1204),
.B(n_1212),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1221),
.B(n_1142),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1221),
.B(n_1204),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1212),
.B(n_1169),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1202),
.B(n_1191),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1217),
.B(n_1136),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1213),
.B(n_1189),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1203),
.B(n_1188),
.C(n_1150),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1222),
.B(n_1178),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1228),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1244),
.B(n_1215),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1235),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1236),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1250),
.B(n_1213),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1247),
.B(n_1208),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1237),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1246),
.B(n_1232),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1253),
.B(n_1232),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1234),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1242),
.B(n_1216),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1263),
.B(n_1234),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1255),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1260),
.B(n_1239),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1258),
.B(n_1238),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1254),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1256),
.A2(n_1239),
.B1(n_1251),
.B2(n_1227),
.C(n_1241),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1259),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1257),
.B(n_1243),
.Y(n_1271)
);

NOR2x1_ASAP7_75t_R g1272 ( 
.A(n_1262),
.B(n_1133),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1261),
.B(n_1240),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1269),
.A2(n_1227),
.B(n_1245),
.Y(n_1274)
);

NOR2x1_ASAP7_75t_SL g1275 ( 
.A(n_1271),
.B(n_1262),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1269),
.B(n_1206),
.C(n_1220),
.Y(n_1276)
);

AND2x2_ASAP7_75t_SL g1277 ( 
.A(n_1266),
.B(n_1249),
.Y(n_1277)
);

XNOR2x1_ASAP7_75t_L g1278 ( 
.A(n_1268),
.B(n_1139),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1265),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1266),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1264),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1280),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1279),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1277),
.B(n_1273),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1281),
.B(n_1267),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1276),
.A2(n_1274),
.B1(n_1262),
.B2(n_1278),
.Y(n_1286)
);

XOR2x2_ASAP7_75t_L g1287 ( 
.A(n_1286),
.B(n_1276),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1282),
.A2(n_1272),
.B(n_1275),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1285),
.B(n_1270),
.Y(n_1289)
);

AND3x1_ASAP7_75t_L g1290 ( 
.A(n_1284),
.B(n_1211),
.C(n_1223),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1283),
.B(n_1160),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1283),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1292),
.Y(n_1293)
);

NOR3x1_ASAP7_75t_L g1294 ( 
.A(n_1287),
.B(n_1223),
.C(n_1210),
.Y(n_1294)
);

OAI211xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1288),
.A2(n_1291),
.B(n_1289),
.C(n_1252),
.Y(n_1295)
);

OAI321xp33_ASAP7_75t_L g1296 ( 
.A1(n_1295),
.A2(n_1290),
.A3(n_1144),
.B1(n_1140),
.B2(n_1248),
.C(n_1224),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_SL g1297 ( 
.A(n_1293),
.B(n_1159),
.C(n_1195),
.Y(n_1297)
);

NOR2x1_ASAP7_75t_L g1298 ( 
.A(n_1297),
.B(n_1182),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1298),
.A2(n_1294),
.B1(n_1296),
.B2(n_1225),
.C(n_1229),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_R g1300 ( 
.A(n_1299),
.B(n_1214),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1299),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1301),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1300),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1302),
.Y(n_1304)
);

OAI22x1_ASAP7_75t_L g1305 ( 
.A1(n_1303),
.A2(n_1134),
.B1(n_1163),
.B2(n_1135),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1304),
.Y(n_1306)
);

OAI22x1_ASAP7_75t_L g1307 ( 
.A1(n_1305),
.A2(n_1186),
.B1(n_1262),
.B2(n_1129),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1306),
.B(n_1231),
.Y(n_1308)
);

INVxp33_ASAP7_75t_SL g1309 ( 
.A(n_1307),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1309),
.A2(n_1231),
.B1(n_1144),
.B2(n_1140),
.Y(n_1310)
);

XNOR2xp5_ASAP7_75t_L g1311 ( 
.A(n_1308),
.B(n_1147),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1311),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1310),
.A2(n_1218),
.B1(n_1080),
.B2(n_1219),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1312),
.B(n_1218),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1314),
.A2(n_1313),
.B1(n_1193),
.B2(n_1113),
.Y(n_1315)
);


endmodule