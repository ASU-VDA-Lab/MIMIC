module real_jpeg_5399_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g133 ( 
.A(n_0),
.Y(n_133)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_179),
.B1(n_181),
.B2(n_185),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_2),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_2),
.A2(n_128),
.B1(n_185),
.B2(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_2),
.A2(n_185),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_3),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_4),
.A2(n_43),
.B1(n_183),
.B2(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_65),
.C(n_177),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_4),
.B(n_129),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_4),
.B(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_4),
.B(n_187),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_4),
.B(n_370),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_5),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_5),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_5),
.A2(n_74),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_6),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_6),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_6),
.A2(n_46),
.B1(n_144),
.B2(n_238),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_6),
.A2(n_144),
.B1(n_197),
.B2(n_306),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_6),
.A2(n_144),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_8),
.Y(n_120)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_9),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_9),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_9),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_10),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_10),
.A2(n_85),
.B1(n_145),
.B2(n_218),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_10),
.A2(n_85),
.B1(n_193),
.B2(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_10),
.A2(n_85),
.B1(n_334),
.B2(n_337),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_13),
.A2(n_61),
.B1(n_76),
.B2(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_14),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_14),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_14),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_15),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_15),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_15),
.A2(n_100),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_15),
.A2(n_100),
.B1(n_182),
.B2(n_209),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_15),
.A2(n_100),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_16),
.A2(n_60),
.B1(n_64),
.B2(n_67),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_16),
.A2(n_67),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_259),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_258),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_221),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_21),
.B(n_221),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_154),
.C(n_205),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_22),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_23),
.B(n_80),
.C(n_113),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_47),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_24),
.A2(n_47),
.B1(n_48),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_24),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.A3(n_33),
.B1(n_36),
.B2(n_42),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_28),
.Y(n_143)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_28),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_29),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_29),
.Y(n_370)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_38),
.A2(n_91),
.B1(n_93),
.B2(n_96),
.Y(n_90)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_42),
.A2(n_43),
.B(n_86),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_43),
.B(n_88),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_43),
.A2(n_49),
.B(n_308),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_SL g366 ( 
.A1(n_43),
.A2(n_367),
.B(n_368),
.Y(n_366)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_58),
.B1(n_68),
.B2(n_72),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_49),
.A2(n_196),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_49),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_50),
.A2(n_73),
.B1(n_195),
.B2(n_202),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_50),
.A2(n_59),
.B1(n_273),
.B2(n_279),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_50),
.B(n_311),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_50),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_56),
.Y(n_201)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_56),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_57),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_62),
.Y(n_313)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_66),
.Y(n_336)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_71),
.Y(n_253)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_71),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_77),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_78),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_112),
.B2(n_113),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_88),
.B(n_98),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_82),
.A2(n_88),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_89),
.B(n_99),
.Y(n_215)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_101),
.Y(n_238)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_104),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_104),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_140),
.B(n_149),
.Y(n_113)
);

AOI22x1_ASAP7_75t_L g227 ( 
.A1(n_114),
.A2(n_129),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_114),
.B(n_228),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_114),
.A2(n_149),
.B(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_115),
.A2(n_141),
.B1(n_153),
.B2(n_217),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_129),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_125),
.B2(n_127),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_124),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_124),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_SL g383 ( 
.A(n_125),
.B(n_384),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_129),
.Y(n_153)
);

AO22x2_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_137),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g319 ( 
.A(n_131),
.Y(n_319)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_133),
.Y(n_301)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_133),
.Y(n_384)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_139),
.Y(n_382)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_150),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_153),
.A2(n_217),
.B(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_154),
.A2(n_155),
.B1(n_205),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_194),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_156),
.B(n_194),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_178),
.B1(n_186),
.B2(n_188),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_157),
.A2(n_292),
.B(n_297),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_157),
.A2(n_186),
.B1(n_318),
.B2(n_360),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_157),
.A2(n_297),
.B(n_360),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_158),
.A2(n_187),
.B1(n_189),
.B2(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_163),
.B1(n_166),
.B2(n_168),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_SL g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_169),
.A2(n_207),
.B(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_174),
.B2(n_176),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_172),
.Y(n_314)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_175),
.Y(n_338)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_186),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_187),
.B(n_208),
.Y(n_297)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_193),
.Y(n_363)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_204),
.Y(n_340)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_216),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_206),
.B(n_216),
.Y(n_264)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_210),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_212),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_241),
.B1(n_256),
.B2(n_257),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_235),
.B1(n_239),
.B2(n_240),
.Y(n_226)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.Y(n_241)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_285),
.B(n_403),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_282),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_262),
.B(n_282),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_269),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_263),
.B(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_269),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.C(n_281),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_270),
.B(n_394),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_272),
.B(n_281),
.Y(n_394)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_277),
.Y(n_307)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_397),
.B(n_402),
.Y(n_285)
);

AO21x1_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_386),
.B(n_396),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_354),
.B(n_385),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_322),
.B(n_353),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_303),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_290),
.B(n_303),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_291),
.A2(n_298),
.B1(n_299),
.B2(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_296),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_315),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_316),
.C(n_321),
.Y(n_355)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_344),
.B(n_352),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_331),
.B(n_343),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_342),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_342),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_339),
.B(n_341),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_350),
.Y(n_352)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_356),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_371),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_364),
.B2(n_365),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_364),
.C(n_371),
.Y(n_387)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

AOI32xp33_ASAP7_75t_L g375 ( 
.A1(n_369),
.A2(n_376),
.A3(n_377),
.B1(n_380),
.B2(n_383),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_375),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_387),
.B(n_388),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_393),
.B2(n_395),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_392),
.C(n_395),
.Y(n_398)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_398),
.B(n_399),
.Y(n_402)
);


endmodule