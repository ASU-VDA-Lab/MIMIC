module fake_ariane_529_n_2099 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2099);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2099;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_274;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_246;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx10_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_26),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_138),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_8),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_105),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_21),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_38),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_143),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_1),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_29),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_99),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_93),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_42),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_80),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_169),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_109),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_62),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_12),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_124),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_134),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_205),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_59),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_115),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_196),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_144),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_38),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_179),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_211),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_85),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_141),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_117),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_81),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_201),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_83),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_104),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_113),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_57),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_33),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_154),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_98),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_63),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_187),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_70),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_67),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_155),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_135),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_175),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_61),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_176),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_123),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_73),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_84),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_198),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_114),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_191),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_20),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_188),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_75),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_46),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_153),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_181),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_63),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_193),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_90),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_132),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_53),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_19),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_116),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_186),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_67),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_53),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_152),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_190),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_164),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_166),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_47),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_3),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_130),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_34),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_110),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_78),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_18),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_70),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_103),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_54),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_150),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_146),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_145),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_28),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_33),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_156),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_10),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_22),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_64),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_58),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_96),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_58),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_180),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_34),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_87),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_64),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_136),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_161),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_28),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_13),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_71),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_22),
.Y(n_350)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_41),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_62),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_168),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_18),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_5),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_17),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_24),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_160),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_91),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_3),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_56),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_208),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_101),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_126),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_69),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_73),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_19),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_184),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_44),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_131),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_54),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_35),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_192),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_69),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_40),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_25),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_119),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_43),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_178),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_167),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_125),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_23),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_68),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_165),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_122),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_36),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_151),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_0),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_7),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_72),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_17),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_142),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_14),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_47),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_74),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_56),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_173),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_162),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_12),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_200),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_41),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_183),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_49),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_182),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_195),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_52),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_68),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_72),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_55),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_36),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_16),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_11),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_159),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_52),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_14),
.Y(n_416)
);

BUFx8_ASAP7_75t_SL g417 ( 
.A(n_120),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_417),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_220),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_259),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_278),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_311),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_217),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_217),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_230),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_381),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_290),
.B(n_0),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_398),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_R g430 ( 
.A(n_238),
.B(n_76),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_408),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_230),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_232),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_215),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_222),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_226),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_232),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_410),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_229),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_233),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_238),
.B(n_5),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_233),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_235),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_250),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_220),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_250),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_253),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_252),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_256),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_290),
.B(n_6),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_252),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_261),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_266),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_266),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_277),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_277),
.B(n_7),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_315),
.B(n_9),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_264),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_282),
.B(n_9),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_262),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_275),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_279),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_282),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_295),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_R g466 ( 
.A(n_301),
.B(n_77),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_218),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_401),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_280),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_212),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_281),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_295),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_225),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_302),
.B(n_10),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_284),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_288),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_297),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_302),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_305),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_218),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_304),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_213),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_212),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_308),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_309),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_212),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_320),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_214),
.B(n_79),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_320),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_313),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_305),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_306),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_319),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_306),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_323),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_307),
.B(n_11),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_307),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_325),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_326),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_316),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_320),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_332),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_340),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_316),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_342),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_406),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_406),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_225),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_324),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_324),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_327),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_406),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_239),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_351),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_327),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_329),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_329),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_213),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_353),
.B(n_15),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_237),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_344),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_353),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_365),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_494),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_467),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_423),
.B(n_382),
.Y(n_532)
);

BUFx8_ASAP7_75t_L g533 ( 
.A(n_482),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_494),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_513),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_423),
.B(n_365),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_424),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_424),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_426),
.B(n_300),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_420),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_437),
.B(n_300),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_374),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_444),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_444),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_446),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_448),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_448),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_451),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_453),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_455),
.B(n_456),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_456),
.B(n_337),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_464),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_465),
.B(n_374),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_472),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_421),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_472),
.B(n_337),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_478),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_479),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_378),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_493),
.B(n_350),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_496),
.A2(n_290),
.B(n_224),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_482),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_499),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_499),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_506),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_506),
.Y(n_585)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_511),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_511),
.A2(n_380),
.B(n_378),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_466),
.B(n_223),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_517),
.B(n_350),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_517),
.B(n_518),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_518),
.B(n_392),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_519),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_380),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_524),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_524),
.B(n_525),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_525),
.B(n_419),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_428),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_520),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_428),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_520),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_450),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_450),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_457),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_460),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_474),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_458),
.B(n_445),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_498),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_509),
.B(n_228),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_SL g613 ( 
.A(n_612),
.B(n_436),
.C(n_435),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_533),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_607),
.A2(n_441),
.B1(n_521),
.B2(n_491),
.Y(n_615)
);

NOR2x1p5_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_418),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_538),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_542),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_530),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_538),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_530),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_509),
.Y(n_623)
);

INVx4_ASAP7_75t_SL g624 ( 
.A(n_586),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_538),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_530),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_530),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_530),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_544),
.Y(n_629)
);

INVx8_ASAP7_75t_L g630 ( 
.A(n_599),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_610),
.B(n_514),
.Y(n_631)
);

BUFx10_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_607),
.B(n_514),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_589),
.A2(n_430),
.B1(n_443),
.B2(n_439),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_530),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_607),
.B(n_447),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_544),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_607),
.B(n_608),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_608),
.B(n_449),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_593),
.B(n_473),
.Y(n_641)
);

AND3x2_ASAP7_75t_L g642 ( 
.A(n_612),
.B(n_548),
.C(n_531),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_544),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_586),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_608),
.A2(n_489),
.B1(n_480),
.B2(n_522),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_608),
.B(n_452),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_541),
.B(n_461),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_586),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_549),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_549),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_551),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_548),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_548),
.B(n_488),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_599),
.B(n_351),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_609),
.B(n_462),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_530),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_551),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_551),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_530),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_553),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_553),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_609),
.B(n_463),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_553),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_541),
.B(n_469),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_541),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_536),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_542),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_609),
.B(n_471),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_611),
.B(n_475),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_541),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_541),
.B(n_558),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_531),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_593),
.B(n_385),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_586),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_533),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_532),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_611),
.A2(n_392),
.B1(n_515),
.B2(n_510),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_554),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_593),
.B(n_599),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_541),
.B(n_558),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_532),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_556),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_611),
.B(n_601),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_601),
.A2(n_390),
.B1(n_260),
.B2(n_476),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_550),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_601),
.B(n_603),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_603),
.A2(n_242),
.B1(n_247),
.B2(n_239),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_586),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_558),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_558),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_556),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_556),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_606),
.B(n_477),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_536),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_589),
.A2(n_484),
.B1(n_485),
.B2(n_481),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_536),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_536),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_533),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_603),
.A2(n_495),
.B1(n_497),
.B2(n_492),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_R g704 ( 
.A(n_588),
.B(n_422),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_558),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_536),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_558),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_560),
.Y(n_708)
);

BUFx4f_ASAP7_75t_L g709 ( 
.A(n_588),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_560),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_540),
.Y(n_711)
);

BUFx4f_ASAP7_75t_L g712 ( 
.A(n_588),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_540),
.B(n_500),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_536),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_605),
.B(n_501),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_605),
.B(n_504),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_533),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_540),
.Y(n_718)
);

AND2x2_ASAP7_75t_SL g719 ( 
.A(n_588),
.B(n_223),
.Y(n_719)
);

INVx6_ASAP7_75t_L g720 ( 
.A(n_586),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_564),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_558),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_536),
.Y(n_724)
);

NOR2x1p5_ASAP7_75t_L g725 ( 
.A(n_561),
.B(n_505),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_588),
.B(n_224),
.Y(n_726)
);

INVxp33_ASAP7_75t_SL g727 ( 
.A(n_545),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_545),
.B(n_507),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_586),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_536),
.Y(n_731)
);

BUFx8_ASAP7_75t_SL g732 ( 
.A(n_594),
.Y(n_732)
);

INVx5_ASAP7_75t_L g733 ( 
.A(n_558),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_564),
.Y(n_734)
);

NOR2x1p5_ASAP7_75t_L g735 ( 
.A(n_561),
.B(n_523),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_564),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_605),
.B(n_242),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_528),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_559),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_545),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_606),
.B(n_243),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_580),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_528),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_606),
.A2(n_588),
.B1(n_594),
.B2(n_579),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_533),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_598),
.B(n_348),
.C(n_347),
.Y(n_746)
);

INVx5_ASAP7_75t_L g747 ( 
.A(n_559),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_563),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_563),
.B(n_247),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_537),
.A2(n_292),
.B1(n_416),
.B2(n_415),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_559),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_600),
.B(n_602),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_555),
.Y(n_753)
);

BUFx4f_ASAP7_75t_L g754 ( 
.A(n_559),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_600),
.B(n_385),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_571),
.B(n_459),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_528),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_559),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_559),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_563),
.B(n_228),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_559),
.B(n_388),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_580),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_594),
.A2(n_352),
.B1(n_416),
.B2(n_415),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_738),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_617),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_688),
.B(n_555),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_620),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_633),
.B(n_555),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_656),
.B(n_555),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_625),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_678),
.B(n_425),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_649),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_618),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_671),
.B(n_555),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_686),
.B(n_555),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_682),
.B(n_623),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_682),
.B(n_562),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_629),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_682),
.B(n_562),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_709),
.Y(n_780)
);

INVx8_ASAP7_75t_L g781 ( 
.A(n_630),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_682),
.A2(n_468),
.B1(n_572),
.B2(n_571),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_649),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_738),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_653),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_743),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_618),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_638),
.Y(n_788)
);

AND2x2_ASAP7_75t_SL g789 ( 
.A(n_744),
.B(n_537),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_682),
.B(n_562),
.Y(n_790)
);

NOR2x1p5_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_631),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_743),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_757),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_639),
.A2(n_598),
.B(n_577),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_669),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_682),
.B(n_562),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_669),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_664),
.B(n_562),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_713),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_630),
.B(n_562),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_675),
.B(n_559),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_630),
.B(n_565),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_630),
.B(n_565),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_753),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_670),
.B(n_565),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_757),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_684),
.B(n_427),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_709),
.B(n_559),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_646),
.B(n_429),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_697),
.B(n_565),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_643),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_709),
.B(n_574),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_655),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_650),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_637),
.B(n_640),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_615),
.A2(n_597),
.B1(n_565),
.B2(n_585),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_651),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_652),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_637),
.B(n_565),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_658),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_659),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_712),
.A2(n_639),
.B(n_641),
.C(n_740),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_661),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_727),
.B(n_597),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_675),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_675),
.A2(n_572),
.B1(n_585),
.B2(n_580),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_640),
.B(n_597),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_642),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_SL g830 ( 
.A(n_616),
.B(n_585),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_655),
.B(n_570),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_712),
.B(n_574),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_727),
.B(n_597),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_647),
.B(n_597),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_647),
.B(n_597),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_632),
.B(n_587),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_712),
.B(n_574),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_663),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_665),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_753),
.B(n_574),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_648),
.A2(n_577),
.B(n_575),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_753),
.B(n_574),
.Y(n_842)
);

CKINVDCx16_ASAP7_75t_R g843 ( 
.A(n_654),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_760),
.B(n_470),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_681),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_641),
.B(n_587),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_711),
.B(n_587),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_632),
.B(n_590),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_654),
.B(n_291),
.C(n_283),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_756),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_685),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_SL g852 ( 
.A(n_614),
.B(n_248),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_632),
.B(n_574),
.Y(n_853)
);

INVxp67_ASAP7_75t_SL g854 ( 
.A(n_677),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_689),
.B(n_760),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_695),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_696),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_741),
.B(n_590),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_675),
.A2(n_595),
.B1(n_590),
.B2(n_594),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_675),
.B(n_595),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_715),
.B(n_716),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_675),
.B(n_595),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_634),
.B(n_533),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_713),
.B(n_276),
.C(n_248),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_728),
.B(n_579),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_708),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_728),
.B(n_579),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_655),
.B(n_570),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_710),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_655),
.A2(n_594),
.B1(n_570),
.B2(n_592),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_719),
.B(n_574),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_720),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_750),
.A2(n_690),
.B1(n_726),
.B2(n_719),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_721),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_750),
.A2(n_529),
.B1(n_535),
.B2(n_528),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_726),
.B(n_574),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_737),
.B(n_579),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_722),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_734),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_736),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_742),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_703),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_748),
.B(n_600),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_729),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_762),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_600),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_752),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_622),
.Y(n_888)
);

NOR2x2_ASAP7_75t_L g889 ( 
.A(n_749),
.B(n_431),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_737),
.B(n_579),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_737),
.B(n_602),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_739),
.B(n_574),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_679),
.B(n_602),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_699),
.B(n_602),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_755),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_749),
.B(n_604),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_704),
.A2(n_594),
.B1(n_592),
.B2(n_576),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_619),
.Y(n_898)
);

AOI221xp5_ASAP7_75t_L g899 ( 
.A1(n_687),
.A2(n_400),
.B1(n_276),
.B2(n_292),
.C(n_303),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_739),
.B(n_578),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_761),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_725),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_739),
.B(n_578),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_749),
.B(n_604),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_749),
.B(n_604),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_729),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_739),
.B(n_578),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_604),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_648),
.A2(n_575),
.B1(n_596),
.B2(n_567),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_763),
.B(n_539),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_690),
.A2(n_576),
.B1(n_592),
.B2(n_567),
.Y(n_911)
);

AND2x6_ASAP7_75t_SL g912 ( 
.A(n_674),
.B(n_303),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_622),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_L g914 ( 
.A(n_746),
.B(n_582),
.C(n_578),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_666),
.B(n_596),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_619),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_674),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_666),
.B(n_539),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_614),
.B(n_539),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_761),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_717),
.B(n_539),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_690),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_622),
.B(n_543),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_717),
.B(n_543),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_662),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_662),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_745),
.B(n_543),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_751),
.B(n_578),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_745),
.B(n_543),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_662),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_667),
.B(n_546),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_667),
.B(n_546),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_794),
.A2(n_754),
.B(n_683),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_818),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_773),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_825),
.B(n_750),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_818),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_825),
.B(n_576),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_797),
.B(n_438),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_833),
.B(n_702),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_808),
.A2(n_754),
.B(n_683),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_764),
.Y(n_942)
);

AOI21xp33_ASAP7_75t_L g943 ( 
.A1(n_809),
.A2(n_702),
.B(n_486),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_841),
.A2(n_754),
.B(n_673),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_799),
.B(n_454),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_833),
.A2(n_354),
.B(n_349),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_861),
.A2(n_547),
.B(n_552),
.C(n_546),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_808),
.A2(n_673),
.B(n_667),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_836),
.A2(n_547),
.B(n_552),
.C(n_546),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_771),
.B(n_483),
.Y(n_950)
);

O2A1O1Ixp5_ASAP7_75t_L g951 ( 
.A1(n_861),
.A2(n_694),
.B(n_705),
.C(n_693),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_766),
.B(n_487),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_781),
.Y(n_953)
);

CKINVDCx10_ASAP7_75t_R g954 ( 
.A(n_843),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_812),
.A2(n_694),
.B(n_693),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_801),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_776),
.B(n_751),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_812),
.A2(n_694),
.B(n_693),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_819),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_764),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_871),
.A2(n_627),
.B(n_626),
.Y(n_961)
);

NOR2x1_ASAP7_75t_L g962 ( 
.A(n_855),
.B(n_547),
.Y(n_962)
);

AOI33xp33_ASAP7_75t_L g963 ( 
.A1(n_899),
.A2(n_336),
.A3(n_312),
.B1(n_318),
.B2(n_321),
.B3(n_328),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_882),
.A2(n_503),
.B1(n_508),
.B2(n_490),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_SL g965 ( 
.A(n_787),
.B(n_732),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_915),
.A2(n_388),
.B(n_526),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_781),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_766),
.B(n_547),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_836),
.B(n_552),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_848),
.B(n_552),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_871),
.A2(n_876),
.B(n_798),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_769),
.A2(n_707),
.B1(n_723),
.B2(n_705),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_848),
.B(n_557),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_832),
.A2(n_707),
.B(n_705),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_876),
.A2(n_627),
.B(n_626),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_846),
.B(n_557),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_847),
.B(n_557),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_804),
.B(n_751),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_798),
.A2(n_635),
.B(n_628),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_804),
.B(n_751),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_774),
.B(n_557),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_786),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_858),
.B(n_566),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_795),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_831),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_918),
.A2(n_635),
.B(n_628),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_816),
.B(n_782),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_886),
.B(n_566),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_886),
.B(n_566),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_831),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_831),
.B(n_624),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_786),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_832),
.A2(n_723),
.B(n_707),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_917),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_810),
.A2(n_730),
.B1(n_723),
.B2(n_759),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_834),
.B(n_835),
.C(n_828),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_837),
.A2(n_759),
.B(n_730),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_918),
.A2(n_657),
.B(n_636),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_777),
.B(n_758),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_837),
.A2(n_759),
.B(n_730),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_781),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_915),
.A2(n_357),
.B(n_355),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_859),
.A2(n_676),
.B1(n_692),
.B2(n_644),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_813),
.B(n_732),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_897),
.B(n_566),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_840),
.A2(n_842),
.B(n_805),
.Y(n_1006)
);

AOI221x1_ASAP7_75t_L g1007 ( 
.A1(n_823),
.A2(n_527),
.B1(n_534),
.B2(n_526),
.C(n_731),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_931),
.A2(n_676),
.B(n_644),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_807),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_772),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_900),
.A2(n_657),
.B(n_636),
.Y(n_1011)
);

OAI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_768),
.A2(n_362),
.B(n_361),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_883),
.B(n_568),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_850),
.B(n_720),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_873),
.A2(n_535),
.B1(n_529),
.B2(n_527),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_840),
.A2(n_676),
.B(n_644),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_842),
.A2(n_692),
.B(n_668),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_838),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_883),
.B(n_568),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_779),
.B(n_790),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_868),
.A2(n_720),
.B1(n_731),
.B2(n_724),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_817),
.A2(n_591),
.B(n_584),
.C(n_581),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_850),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_868),
.B(n_826),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_912),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_864),
.A2(n_591),
.B(n_584),
.C(n_581),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_868),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_923),
.A2(n_668),
.B(n_660),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_911),
.B(n_789),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_789),
.B(n_568),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_775),
.A2(n_692),
.B(n_691),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_853),
.A2(n_691),
.B(n_660),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_870),
.B(n_568),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_838),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_785),
.B(n_573),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_853),
.A2(n_700),
.B(n_698),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_829),
.B(n_624),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_L g1038 ( 
.A(n_826),
.B(n_758),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_873),
.A2(n_700),
.B(n_698),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_844),
.B(n_573),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_823),
.A2(n_581),
.B(n_584),
.C(n_591),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_852),
.A2(n_701),
.B(n_706),
.C(n_714),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_830),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_922),
.A2(n_535),
.B1(n_529),
.B2(n_527),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_800),
.A2(n_803),
.B(n_802),
.Y(n_1045)
);

AO21x1_ASAP7_75t_L g1046 ( 
.A1(n_894),
.A2(n_534),
.B(n_526),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_895),
.B(n_573),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_902),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_796),
.B(n_758),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_908),
.B(n_573),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_865),
.B(n_581),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_888),
.A2(n_706),
.B(n_701),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_792),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_923),
.A2(n_724),
.B(n_714),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_765),
.B(n_767),
.Y(n_1055)
);

OAI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_770),
.A2(n_367),
.B(n_366),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_888),
.A2(n_758),
.B(n_621),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_896),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_778),
.B(n_584),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_L g1060 ( 
.A1(n_900),
.A2(n_577),
.B(n_591),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_826),
.B(n_621),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_854),
.Y(n_1062)
);

INVx11_ASAP7_75t_L g1063 ( 
.A(n_889),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_788),
.B(n_534),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_869),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_904),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_913),
.A2(n_621),
.B(n_672),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_772),
.B(n_672),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_772),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_867),
.B(n_621),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_849),
.B(n_624),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_827),
.B(n_672),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_905),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_SL g1074 ( 
.A1(n_860),
.A2(n_577),
.B(n_318),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_913),
.A2(n_680),
.B(n_672),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_811),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_814),
.B(n_578),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_780),
.B(n_821),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_932),
.A2(n_680),
.B(n_672),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_822),
.B(n_372),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_824),
.B(n_373),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_772),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_791),
.B(n_228),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_L g1084 ( 
.A(n_862),
.B(n_680),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_792),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_815),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_932),
.A2(n_926),
.B(n_925),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_930),
.A2(n_733),
.B(n_680),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_909),
.B(n_845),
.C(n_839),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_903),
.A2(n_733),
.B(n_680),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_869),
.A2(n_400),
.B(n_375),
.C(n_368),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_903),
.A2(n_747),
.B(n_733),
.Y(n_1092)
);

BUFx4f_ASAP7_75t_L g1093 ( 
.A(n_857),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_894),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_866),
.B(n_321),
.C(n_312),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_891),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_907),
.A2(n_928),
.B(n_914),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_874),
.B(n_578),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_878),
.Y(n_1099)
);

AOI22x1_ASAP7_75t_L g1100 ( 
.A1(n_878),
.A2(n_578),
.B1(n_583),
.B2(n_582),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_879),
.B(n_333),
.C(n_328),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_907),
.A2(n_529),
.B(n_535),
.C(n_413),
.Y(n_1102)
);

INVx11_ASAP7_75t_L g1103 ( 
.A(n_875),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_881),
.A2(n_336),
.B(n_375),
.C(n_370),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_910),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_928),
.A2(n_747),
.B(n_733),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_880),
.B(n_376),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_783),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_881),
.A2(n_338),
.B(n_370),
.C(n_384),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_793),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_851),
.B(n_582),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_856),
.B(n_379),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_885),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_793),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_887),
.B(n_582),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_901),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_898),
.A2(n_916),
.B(n_892),
.Y(n_1117)
);

OAI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_885),
.A2(n_389),
.B(n_387),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_887),
.A2(n_747),
.B(n_733),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_783),
.B(n_884),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_920),
.A2(n_356),
.B1(n_293),
.B2(n_289),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1094),
.A2(n_890),
.B1(n_877),
.B2(n_863),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_934),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_952),
.A2(n_384),
.B(n_404),
.C(n_333),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_938),
.B(n_893),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_954),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1103),
.A2(n_875),
.B1(n_394),
.B2(n_335),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_969),
.A2(n_921),
.B(n_919),
.Y(n_1128)
);

OAI22x1_ASAP7_75t_L g1129 ( 
.A1(n_964),
.A2(n_338),
.B1(n_394),
.B2(n_335),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_987),
.A2(n_404),
.B1(n_368),
.B2(n_377),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_970),
.A2(n_927),
.B(n_924),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_950),
.B(n_1009),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_973),
.A2(n_929),
.B(n_806),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_987),
.A2(n_872),
.B1(n_884),
.B2(n_906),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_942),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_SL g1136 ( 
.A(n_953),
.B(n_1001),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_939),
.Y(n_1137)
);

NOR2x1_ASAP7_75t_R g1138 ( 
.A(n_935),
.B(n_395),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_937),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_936),
.A2(n_413),
.B1(n_391),
.B2(n_352),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_940),
.B(n_1076),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1001),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_991),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1024),
.B(n_872),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1025),
.A2(n_411),
.B1(n_397),
.B2(n_407),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1013),
.A2(n_806),
.B(n_783),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1040),
.B(n_784),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_991),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_959),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1023),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1078),
.A2(n_356),
.B(n_293),
.C(n_286),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1029),
.A2(n_377),
.B1(n_391),
.B2(n_783),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1078),
.B(n_582),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1019),
.A2(n_906),
.B(n_884),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1002),
.A2(n_414),
.B(n_241),
.C(n_251),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_1076),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_960),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1055),
.A2(n_906),
.B1(n_884),
.B2(n_582),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_946),
.A2(n_414),
.B(n_241),
.C(n_251),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1058),
.B(n_582),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_945),
.B(n_906),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1001),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1058),
.B(n_582),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_982),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1073),
.B(n_583),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_SL g1166 ( 
.A(n_1095),
.B(n_402),
.C(n_409),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1024),
.B(n_624),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_988),
.A2(n_747),
.B(n_583),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1024),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1001),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1089),
.A2(n_1070),
.B(n_1093),
.C(n_971),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_994),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1062),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1093),
.B(n_583),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1004),
.B(n_268),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_747),
.B(n_583),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_984),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1095),
.A2(n_237),
.B(n_258),
.C(n_268),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1048),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_943),
.A2(n_358),
.B1(n_268),
.B2(n_258),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_SL g1181 ( 
.A(n_953),
.B(n_967),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1069),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_965),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_979),
.A2(n_583),
.B(n_216),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1089),
.A2(n_583),
.B(n_405),
.C(n_403),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1070),
.A2(n_583),
.B(n_399),
.C(n_396),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1030),
.B(n_15),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1018),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1034),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_985),
.B(n_236),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1031),
.A2(n_393),
.B(n_386),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1116),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_985),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_1004),
.B(n_219),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_990),
.B(n_358),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_1043),
.B(n_369),
.C(n_364),
.Y(n_1196)
);

BUFx8_ASAP7_75t_SL g1197 ( 
.A(n_1083),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_990),
.B(n_221),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_992),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_956),
.A2(n_363),
.B1(n_360),
.B2(n_359),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1063),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1027),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1101),
.A2(n_346),
.B(n_345),
.C(n_343),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1101),
.A2(n_341),
.B(n_339),
.C(n_334),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1045),
.A2(n_270),
.B(n_330),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_956),
.A2(n_269),
.B1(n_231),
.B2(n_317),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1065),
.B(n_1099),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_967),
.B(n_227),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1041),
.A2(n_234),
.B(n_240),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1012),
.A2(n_272),
.B(n_244),
.C(n_314),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1113),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1027),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1066),
.B(n_16),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1096),
.B(n_20),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1035),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1105),
.B(n_21),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1080),
.B(n_1081),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1080),
.B(n_25),
.Y(n_1218)
);

BUFx12f_ASAP7_75t_L g1219 ( 
.A(n_1069),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1086),
.B(n_245),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1091),
.A2(n_26),
.B(n_27),
.C(n_29),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_996),
.A2(n_273),
.B(n_246),
.C(n_310),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1064),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_949),
.A2(n_331),
.B(n_322),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1053),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1014),
.B(n_249),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1014),
.B(n_254),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_981),
.A2(n_274),
.B(n_255),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1105),
.B(n_27),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1037),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1069),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1069),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1091),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1081),
.B(n_30),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_976),
.A2(n_285),
.B1(n_257),
.B2(n_299),
.Y(n_1235)
);

BUFx12f_ASAP7_75t_SL g1236 ( 
.A(n_1082),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1107),
.B(n_31),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1008),
.A2(n_287),
.B(n_263),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_SL g1239 ( 
.A1(n_957),
.A2(n_331),
.B(n_322),
.C(n_236),
.Y(n_1239)
);

NOR2x1_ASAP7_75t_L g1240 ( 
.A(n_1010),
.B(n_331),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1107),
.B(n_265),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1085),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1112),
.B(n_32),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1037),
.B(n_35),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_L g1245 ( 
.A1(n_966),
.A2(n_37),
.B(n_40),
.C(n_42),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1028),
.A2(n_294),
.B(n_267),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1054),
.A2(n_298),
.B(n_296),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1082),
.Y(n_1248)
);

OR2x4_ASAP7_75t_L g1249 ( 
.A(n_1112),
.B(n_37),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_968),
.A2(n_271),
.B(n_322),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1082),
.B(n_331),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1119),
.A2(n_331),
.B(n_322),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1110),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1082),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_983),
.A2(n_322),
.B(n_236),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1032),
.A2(n_236),
.B(n_108),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1108),
.B(n_236),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_963),
.B(n_44),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_977),
.B(n_45),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1108),
.Y(n_1260)
);

BUFx2_ASAP7_75t_SL g1261 ( 
.A(n_1108),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1108),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1056),
.B(n_45),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1010),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1033),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1114),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1118),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1020),
.B(n_48),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1104),
.A2(n_50),
.B(n_51),
.C(n_55),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1120),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1044),
.B(n_50),
.Y(n_1271)
);

CKINVDCx8_ASAP7_75t_R g1272 ( 
.A(n_1071),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1036),
.A2(n_127),
.B(n_206),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1088),
.A2(n_121),
.B(n_204),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1104),
.A2(n_51),
.B(n_59),
.C(n_60),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1109),
.B(n_60),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1120),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1044),
.B(n_1047),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_955),
.A2(n_128),
.B(n_202),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1071),
.B(n_65),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1059),
.A2(n_65),
.B1(n_66),
.B2(n_82),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1007),
.A2(n_129),
.B(n_88),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1219),
.Y(n_1283)
);

BUFx12f_ASAP7_75t_L g1284 ( 
.A(n_1126),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1217),
.A2(n_1121),
.B(n_1109),
.C(n_1026),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1169),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1215),
.B(n_1015),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1207),
.Y(n_1288)
);

AO32x2_ASAP7_75t_L g1289 ( 
.A1(n_1140),
.A2(n_995),
.A3(n_972),
.B1(n_1046),
.B2(n_1041),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1141),
.B(n_1192),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1241),
.B(n_962),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1171),
.A2(n_951),
.B(n_948),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1150),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1123),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1280),
.B(n_1061),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1172),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1125),
.A2(n_1005),
.B(n_1061),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1227),
.A2(n_1006),
.B(n_1087),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1147),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1173),
.B(n_1015),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1256),
.A2(n_1011),
.B(n_1060),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1128),
.A2(n_1038),
.B(n_933),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1137),
.B(n_1020),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1223),
.B(n_947),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1132),
.B(n_1021),
.Y(n_1305)
);

OAI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1218),
.A2(n_1077),
.B(n_1098),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1135),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1252),
.A2(n_1117),
.A3(n_941),
.B(n_1115),
.Y(n_1308)
);

OAI22x1_ASAP7_75t_L g1309 ( 
.A1(n_1237),
.A2(n_957),
.B1(n_1049),
.B2(n_999),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1139),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1187),
.A2(n_1097),
.B(n_975),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1183),
.B(n_1049),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1158),
.A2(n_1052),
.A3(n_997),
.B(n_1000),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1273),
.A2(n_944),
.B(n_986),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1131),
.A2(n_1072),
.B(n_1084),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1197),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1231),
.B(n_978),
.Y(n_1317)
);

INVx3_ASAP7_75t_SL g1318 ( 
.A(n_1201),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1207),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1234),
.A2(n_1072),
.B(n_999),
.C(n_1022),
.Y(n_1320)
);

AO32x2_ASAP7_75t_L g1321 ( 
.A1(n_1140),
.A2(n_1003),
.A3(n_1074),
.B1(n_1039),
.B2(n_1051),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1157),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1161),
.B(n_1050),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1255),
.A2(n_998),
.B(n_1042),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1175),
.B(n_1111),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1149),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_SL g1327 ( 
.A(n_1272),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1153),
.A2(n_1133),
.B(n_1158),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1188),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1164),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1185),
.A2(n_958),
.A3(n_974),
.B(n_993),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1169),
.B(n_978),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1280),
.B(n_1068),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1243),
.A2(n_1102),
.B(n_961),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1146),
.A2(n_1100),
.B(n_1057),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1244),
.B(n_1156),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1209),
.A2(n_1075),
.B(n_1067),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1169),
.B(n_980),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1179),
.B(n_980),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1189),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1127),
.B(n_1068),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1177),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1211),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1169),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1199),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1127),
.B(n_1106),
.Y(n_1346)
);

INVxp67_ASAP7_75t_SL g1347 ( 
.A(n_1230),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1154),
.A2(n_1079),
.B(n_1016),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1239),
.A2(n_1017),
.B(n_1092),
.Y(n_1349)
);

AOI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1184),
.A2(n_1090),
.B(n_89),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1225),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1166),
.A2(n_66),
.B(n_94),
.C(n_95),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1186),
.A2(n_100),
.A3(n_102),
.B(n_107),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1242),
.Y(n_1354)
);

NAND3x1_ASAP7_75t_L g1355 ( 
.A(n_1263),
.B(n_111),
.C(n_118),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1202),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1253),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1279),
.A2(n_137),
.B(n_140),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1250),
.A2(n_147),
.B(n_174),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1193),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1266),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1216),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1216),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1168),
.A2(n_177),
.B(n_194),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1176),
.A2(n_197),
.B(n_210),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1274),
.A2(n_1278),
.B(n_1259),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1130),
.B(n_1212),
.Y(n_1367)
);

AOI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1124),
.A2(n_1155),
.B(n_1206),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1240),
.A2(n_1282),
.B(n_1209),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1130),
.A2(n_1268),
.B(n_1229),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1129),
.A2(n_1276),
.B1(n_1180),
.B2(n_1267),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1282),
.A2(n_1257),
.B(n_1251),
.Y(n_1372)
);

AO21x1_ASAP7_75t_L g1373 ( 
.A1(n_1187),
.A2(n_1265),
.B(n_1281),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1143),
.B(n_1148),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1244),
.B(n_1280),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1151),
.A2(n_1204),
.B1(n_1203),
.B2(n_1235),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1265),
.A2(n_1195),
.B1(n_1258),
.B2(n_1198),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1178),
.A2(n_1159),
.B(n_1222),
.C(n_1122),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1160),
.A2(n_1163),
.B(n_1165),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1213),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1246),
.A2(n_1247),
.B(n_1205),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1214),
.B(n_1143),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1248),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1271),
.A2(n_1233),
.B(n_1275),
.C(n_1269),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1224),
.A2(n_1245),
.B(n_1134),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1230),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1148),
.B(n_1220),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1152),
.A2(n_1281),
.A3(n_1210),
.B(n_1235),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1224),
.A2(n_1174),
.B(n_1226),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1152),
.B(n_1190),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1270),
.A2(n_1248),
.B(n_1191),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1145),
.A2(n_1206),
.B1(n_1200),
.B2(n_1194),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1221),
.A2(n_1200),
.B(n_1208),
.C(n_1196),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1277),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1228),
.A2(n_1238),
.B(n_1270),
.C(n_1136),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1254),
.A2(n_1262),
.B(n_1264),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1142),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1190),
.B(n_1144),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1249),
.A2(n_1262),
.A3(n_1254),
.B(n_1190),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1144),
.A2(n_1249),
.B(n_1167),
.C(n_1181),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1182),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1142),
.A2(n_1162),
.B1(n_1170),
.B2(n_1261),
.Y(n_1402)
);

NAND2x1_ASAP7_75t_L g1403 ( 
.A(n_1182),
.B(n_1232),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1167),
.A2(n_1260),
.B(n_1232),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1236),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1217),
.A2(n_773),
.B1(n_669),
.B2(n_618),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1137),
.B(n_945),
.Y(n_1407)
);

NOR4xp25_ASAP7_75t_L g1408 ( 
.A(n_1218),
.B(n_1234),
.C(n_1217),
.D(n_1243),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1217),
.B(n_773),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1207),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_956),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1217),
.A2(n_1094),
.B1(n_1241),
.B2(n_940),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1217),
.A2(n_1241),
.B(n_1218),
.C(n_1234),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1138),
.B(n_773),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1217),
.A2(n_1241),
.B(n_1218),
.C(n_1234),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1135),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1217),
.A2(n_773),
.B1(n_669),
.B2(n_618),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1217),
.A2(n_1241),
.B(n_1218),
.C(n_1234),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1252),
.A2(n_1046),
.A3(n_1007),
.B(n_966),
.Y(n_1419)
);

NAND2x2_ASAP7_75t_L g1420 ( 
.A(n_1126),
.B(n_935),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_956),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1217),
.A2(n_1094),
.B1(n_1241),
.B2(n_940),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1241),
.A2(n_940),
.B(n_1217),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1280),
.B(n_1024),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_956),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1135),
.Y(n_1426)
);

AOI221x1_ASAP7_75t_L g1427 ( 
.A1(n_1265),
.A2(n_1281),
.B1(n_1130),
.B2(n_1171),
.C(n_1234),
.Y(n_1427)
);

AND3x4_ASAP7_75t_L g1428 ( 
.A(n_1196),
.B(n_935),
.C(n_1194),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_SL g1429 ( 
.A1(n_1171),
.A2(n_1141),
.B(n_940),
.C(n_1218),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1207),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1217),
.B(n_678),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_956),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1256),
.A2(n_1011),
.B(n_1060),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1217),
.A2(n_1241),
.B(n_1218),
.C(n_1234),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_956),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1217),
.A2(n_1241),
.B(n_1218),
.C(n_1234),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1135),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1241),
.A2(n_940),
.B(n_1217),
.Y(n_1438)
);

AO21x1_ASAP7_75t_L g1439 ( 
.A1(n_1243),
.A2(n_1234),
.B(n_1218),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1123),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1219),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1249),
.A2(n_773),
.B1(n_669),
.B2(n_618),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1219),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1217),
.B(n_678),
.Y(n_1444)
);

AO31x2_ASAP7_75t_L g1445 ( 
.A1(n_1252),
.A2(n_1046),
.A3(n_1007),
.B(n_966),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1156),
.B(n_618),
.Y(n_1446)
);

AO32x2_ASAP7_75t_L g1447 ( 
.A1(n_1140),
.A2(n_1130),
.A3(n_1265),
.B1(n_1152),
.B2(n_1127),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1123),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1217),
.B(n_678),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1241),
.A2(n_940),
.B(n_1217),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_SL g1451 ( 
.A1(n_1171),
.A2(n_1141),
.B(n_940),
.C(n_1218),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1294),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1288),
.B(n_1319),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1288),
.B(n_1319),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1410),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1296),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1310),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_SL g1458 ( 
.A(n_1284),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1397),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1293),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1371),
.A2(n_1370),
.B1(n_1373),
.B2(n_1439),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1440),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_1316),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1412),
.A2(n_1422),
.B1(n_1450),
.B2(n_1423),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1405),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1392),
.A2(n_1406),
.B1(n_1417),
.B2(n_1438),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1411),
.A2(n_1425),
.B(n_1421),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1318),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1448),
.Y(n_1469)
);

INVx6_ASAP7_75t_L g1470 ( 
.A(n_1443),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1390),
.A2(n_1442),
.B1(n_1305),
.B2(n_1287),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1427),
.A2(n_1346),
.B1(n_1367),
.B2(n_1449),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1368),
.A2(n_1380),
.B1(n_1376),
.B2(n_1363),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1326),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1413),
.A2(n_1418),
.B(n_1415),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1443),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1362),
.A2(n_1407),
.B1(n_1409),
.B2(n_1444),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1431),
.A2(n_1414),
.B1(n_1295),
.B2(n_1424),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1299),
.A2(n_1437),
.B1(n_1330),
.B2(n_1322),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1443),
.Y(n_1480)
);

BUFx10_ASAP7_75t_L g1481 ( 
.A(n_1342),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1307),
.A2(n_1416),
.B1(n_1426),
.B2(n_1291),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1360),
.Y(n_1483)
);

CKINVDCx6p67_ASAP7_75t_R g1484 ( 
.A(n_1283),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1295),
.A2(n_1424),
.B1(n_1387),
.B2(n_1420),
.Y(n_1485)
);

BUFx10_ASAP7_75t_L g1486 ( 
.A(n_1303),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1345),
.A2(n_1354),
.B1(n_1361),
.B2(n_1357),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1283),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1300),
.A2(n_1341),
.B1(n_1333),
.B2(n_1325),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1351),
.A2(n_1430),
.B1(n_1410),
.B2(n_1375),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1430),
.B(n_1408),
.Y(n_1491)
);

BUFx2_ASAP7_75t_R g1492 ( 
.A(n_1336),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1356),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1333),
.A2(n_1382),
.B1(n_1446),
.B2(n_1398),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1329),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1329),
.Y(n_1496)
);

BUFx12f_ASAP7_75t_L g1497 ( 
.A(n_1441),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1327),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1312),
.A2(n_1441),
.B1(n_1377),
.B2(n_1340),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1434),
.A2(n_1436),
.B(n_1393),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1428),
.A2(n_1343),
.B1(n_1323),
.B2(n_1447),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1290),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1383),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1317),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1285),
.A2(n_1384),
.B1(n_1304),
.B2(n_1378),
.Y(n_1505)
);

BUFx4f_ASAP7_75t_SL g1506 ( 
.A(n_1401),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1298),
.A2(n_1366),
.B(n_1320),
.Y(n_1507)
);

BUFx2_ASAP7_75t_SL g1508 ( 
.A(n_1339),
.Y(n_1508)
);

OAI22x1_ASAP7_75t_SL g1509 ( 
.A1(n_1386),
.A2(n_1401),
.B1(n_1447),
.B2(n_1383),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1447),
.A2(n_1385),
.B1(n_1311),
.B2(n_1334),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1429),
.B(n_1451),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1394),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1404),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1404),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1286),
.Y(n_1515)
);

CKINVDCx6p67_ASAP7_75t_R g1516 ( 
.A(n_1374),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1400),
.A2(n_1355),
.B1(n_1389),
.B2(n_1347),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1385),
.A2(n_1306),
.B1(n_1302),
.B2(n_1352),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1286),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1328),
.A2(n_1292),
.B1(n_1435),
.B2(n_1432),
.Y(n_1520)
);

CKINVDCx6p67_ASAP7_75t_R g1521 ( 
.A(n_1309),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1369),
.A2(n_1321),
.B1(n_1388),
.B2(n_1332),
.Y(n_1522)
);

BUFx10_ASAP7_75t_L g1523 ( 
.A(n_1332),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1402),
.Y(n_1524)
);

INVx11_ASAP7_75t_L g1525 ( 
.A(n_1403),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1338),
.A2(n_1344),
.B1(n_1337),
.B2(n_1396),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1344),
.B(n_1391),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1399),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1315),
.A2(n_1348),
.B(n_1314),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1388),
.B(n_1344),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1395),
.A2(n_1297),
.B1(n_1381),
.B2(n_1365),
.Y(n_1531)
);

INVx6_ASAP7_75t_L g1532 ( 
.A(n_1388),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1364),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1289),
.A2(n_1350),
.B1(n_1324),
.B2(n_1321),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1379),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1324),
.A2(n_1372),
.B1(n_1358),
.B2(n_1321),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1359),
.A2(n_1289),
.B(n_1353),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1353),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1353),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1289),
.A2(n_1445),
.B1(n_1419),
.B2(n_1301),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1419),
.B(n_1445),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1313),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1313),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1433),
.A2(n_1349),
.B1(n_1335),
.B2(n_1331),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1331),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1308),
.Y(n_1546)
);

BUFx12f_ASAP7_75t_L g1547 ( 
.A(n_1331),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1308),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1308),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1442),
.A2(n_1249),
.B1(n_773),
.B2(n_1409),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1288),
.B(n_1319),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1409),
.B(n_1431),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1367),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1296),
.Y(n_1555)
);

INVx6_ASAP7_75t_L g1556 ( 
.A(n_1443),
.Y(n_1556)
);

INVx6_ASAP7_75t_L g1557 ( 
.A(n_1443),
.Y(n_1557)
);

CKINVDCx16_ASAP7_75t_R g1558 ( 
.A(n_1414),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1377),
.A2(n_1127),
.B1(n_1217),
.B2(n_612),
.Y(n_1559)
);

CKINVDCx11_ASAP7_75t_R g1560 ( 
.A(n_1284),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1316),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1346),
.A2(n_1094),
.B1(n_1103),
.B2(n_1218),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1294),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1375),
.A2(n_1217),
.B1(n_1237),
.B2(n_1129),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1288),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1307),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1406),
.A2(n_669),
.B1(n_618),
.B2(n_773),
.Y(n_1568)
);

INVx6_ASAP7_75t_L g1569 ( 
.A(n_1443),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1316),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1392),
.A2(n_1217),
.B(n_1427),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1294),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1294),
.Y(n_1574)
);

BUFx2_ASAP7_75t_SL g1575 ( 
.A(n_1446),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1443),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1405),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1406),
.A2(n_669),
.B1(n_618),
.B2(n_773),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1427),
.A2(n_1249),
.B1(n_1392),
.B2(n_1346),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1405),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1342),
.Y(n_1582)
);

INVx6_ASAP7_75t_L g1583 ( 
.A(n_1443),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1346),
.A2(n_1094),
.B1(n_1103),
.B2(n_1218),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1442),
.A2(n_1249),
.B1(n_773),
.B2(n_1409),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1377),
.A2(n_1127),
.B1(n_1217),
.B2(n_612),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1427),
.A2(n_1249),
.B1(n_1392),
.B2(n_1346),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1392),
.A2(n_1217),
.B(n_1427),
.Y(n_1590)
);

INVx8_ASAP7_75t_L g1591 ( 
.A(n_1424),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1294),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1294),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1371),
.A2(n_1217),
.B1(n_943),
.B2(n_809),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1294),
.Y(n_1597)
);

BUFx12f_ASAP7_75t_L g1598 ( 
.A(n_1284),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1397),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1288),
.B(n_1319),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1296),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1294),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1554),
.B(n_1472),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1474),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1495),
.Y(n_1605)
);

CKINVDCx6p67_ASAP7_75t_R g1606 ( 
.A(n_1558),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1496),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1554),
.B(n_1455),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1455),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1565),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1472),
.B(n_1464),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1529),
.A2(n_1467),
.B(n_1531),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1503),
.Y(n_1613)
);

AO31x2_ASAP7_75t_L g1614 ( 
.A1(n_1534),
.A2(n_1518),
.A3(n_1538),
.B(n_1539),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1527),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1506),
.Y(n_1616)
);

AO21x1_ASAP7_75t_SL g1617 ( 
.A1(n_1507),
.A2(n_1511),
.B(n_1491),
.Y(n_1617)
);

AO21x2_ASAP7_75t_L g1618 ( 
.A1(n_1537),
.A2(n_1534),
.B(n_1518),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1541),
.B(n_1565),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1491),
.A2(n_1530),
.B(n_1546),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1504),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1568),
.B(n_1579),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1453),
.Y(n_1623)
);

AOI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1531),
.A2(n_1529),
.B(n_1511),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1454),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1454),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1461),
.A2(n_1505),
.B(n_1562),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1467),
.A2(n_1507),
.B(n_1544),
.Y(n_1628)
);

CKINVDCx11_ASAP7_75t_R g1629 ( 
.A(n_1560),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1452),
.B(n_1457),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1555),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1475),
.A2(n_1500),
.B(n_1587),
.C(n_1559),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1520),
.A2(n_1543),
.B(n_1536),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1462),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1551),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1553),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1520),
.A2(n_1505),
.B(n_1562),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1469),
.B(n_1563),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1600),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1573),
.B(n_1574),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1600),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1584),
.B(n_1501),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1543),
.A2(n_1527),
.B(n_1535),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1547),
.Y(n_1647)
);

AND2x6_ASAP7_75t_L g1648 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1649)
);

INVxp33_ASAP7_75t_L g1650 ( 
.A(n_1493),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1559),
.A2(n_1587),
.B1(n_1588),
.B2(n_1566),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1597),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1504),
.Y(n_1653)
);

AOI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1517),
.A2(n_1584),
.B(n_1528),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1545),
.A2(n_1589),
.B(n_1580),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1456),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1545),
.A2(n_1526),
.B(n_1517),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1572),
.A2(n_1590),
.B1(n_1466),
.B2(n_1589),
.Y(n_1658)
);

OAI322xp33_ASAP7_75t_L g1659 ( 
.A1(n_1580),
.A2(n_1499),
.A3(n_1564),
.B1(n_1489),
.B2(n_1485),
.C1(n_1478),
.C2(n_1550),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1473),
.B(n_1477),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1509),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1510),
.B(n_1540),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1591),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1542),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1515),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1494),
.A2(n_1512),
.B(n_1567),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1525),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1591),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1522),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1502),
.Y(n_1670)
);

CKINVDCx6p67_ASAP7_75t_R g1671 ( 
.A(n_1463),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1522),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1471),
.B(n_1516),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1591),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1510),
.B(n_1540),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1549),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1521),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1487),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1490),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1533),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1486),
.B(n_1548),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1459),
.A2(n_1599),
.B(n_1482),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1483),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1552),
.A2(n_1592),
.B(n_1585),
.Y(n_1684)
);

OAI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1571),
.A2(n_1576),
.B(n_1595),
.C(n_1596),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1599),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1479),
.A2(n_1519),
.B(n_1523),
.Y(n_1687)
);

AOI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1486),
.A2(n_1508),
.B(n_1581),
.Y(n_1688)
);

CKINVDCx8_ASAP7_75t_R g1689 ( 
.A(n_1575),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1519),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1519),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1524),
.Y(n_1692)
);

AND2x2_ASAP7_75t_SL g1693 ( 
.A(n_1480),
.B(n_1492),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1470),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1476),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1582),
.B(n_1481),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1498),
.B(n_1586),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1476),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1488),
.A2(n_1497),
.B1(n_1583),
.B2(n_1577),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1481),
.B(n_1556),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1557),
.A2(n_1569),
.B1(n_1583),
.B2(n_1577),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1557),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1569),
.A2(n_1577),
.B1(n_1598),
.B2(n_1484),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1569),
.Y(n_1704)
);

AND2x2_ASAP7_75t_SL g1705 ( 
.A(n_1578),
.B(n_1458),
.Y(n_1705)
);

AND2x4_ASAP7_75t_SL g1706 ( 
.A(n_1578),
.B(n_1465),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1468),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1460),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1561),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1570),
.B(n_1541),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1529),
.A2(n_1467),
.B(n_1531),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1635),
.B(n_1646),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1608),
.B(n_1637),
.Y(n_1713)
);

AOI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1658),
.A2(n_1633),
.B(n_1627),
.C(n_1659),
.Y(n_1714)
);

O2A1O1Ixp33_ASAP7_75t_L g1715 ( 
.A1(n_1627),
.A2(n_1611),
.B(n_1622),
.C(n_1638),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1612),
.A2(n_1711),
.B(n_1628),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1710),
.B(n_1656),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1612),
.A2(n_1711),
.B(n_1628),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_SL g1719 ( 
.A1(n_1688),
.A2(n_1653),
.B(n_1621),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1632),
.Y(n_1720)
);

O2A1O1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1603),
.A2(n_1660),
.B(n_1644),
.C(n_1684),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1634),
.A2(n_1657),
.B(n_1687),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1651),
.A2(n_1661),
.B(n_1675),
.C(n_1662),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1662),
.A2(n_1675),
.B1(n_1685),
.B2(n_1655),
.C(n_1669),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1629),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1647),
.B(n_1619),
.Y(n_1726)
);

AO32x2_ASAP7_75t_L g1727 ( 
.A1(n_1615),
.A2(n_1653),
.A3(n_1621),
.B1(n_1617),
.B2(n_1663),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1650),
.B(n_1632),
.Y(n_1728)
);

INVx4_ASAP7_75t_SL g1729 ( 
.A(n_1708),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1647),
.B(n_1619),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1631),
.B(n_1630),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1673),
.A2(n_1693),
.B(n_1672),
.C(n_1669),
.Y(n_1732)
);

AO32x2_ASAP7_75t_L g1733 ( 
.A1(n_1615),
.A2(n_1653),
.A3(n_1617),
.B1(n_1674),
.B2(n_1668),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1639),
.B(n_1642),
.Y(n_1735)
);

AO21x1_ASAP7_75t_L g1736 ( 
.A1(n_1677),
.A2(n_1692),
.B(n_1652),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1652),
.B(n_1639),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1654),
.A2(n_1624),
.B(n_1657),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1642),
.B(n_1649),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1604),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1640),
.B(n_1708),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1654),
.A2(n_1624),
.B(n_1682),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1709),
.B(n_1696),
.C(n_1697),
.D(n_1616),
.Y(n_1743)
);

AO32x2_ASAP7_75t_L g1744 ( 
.A1(n_1663),
.A2(n_1674),
.A3(n_1668),
.B1(n_1616),
.B2(n_1655),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1693),
.A2(n_1672),
.B1(n_1689),
.B2(n_1703),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1689),
.A2(n_1681),
.B1(n_1703),
.B2(n_1699),
.C(n_1692),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1628),
.A2(n_1681),
.B(n_1610),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1628),
.B(n_1704),
.C(n_1698),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1604),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1645),
.A2(n_1676),
.B(n_1664),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1616),
.A2(n_1670),
.B(n_1709),
.C(n_1667),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1686),
.B(n_1696),
.Y(n_1752)
);

AO32x2_ASAP7_75t_L g1753 ( 
.A1(n_1618),
.A2(n_1620),
.A3(n_1679),
.B1(n_1678),
.B2(n_1666),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1698),
.B(n_1704),
.C(n_1609),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1623),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1606),
.B(n_1700),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1671),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1707),
.B(n_1683),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1693),
.A2(n_1705),
.B1(n_1667),
.B2(n_1665),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1625),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1618),
.A2(n_1702),
.B(n_1694),
.C(n_1695),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1671),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1690),
.A2(n_1691),
.B(n_1680),
.C(n_1676),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1626),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1636),
.B(n_1643),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1706),
.B(n_1705),
.Y(n_1766)
);

CKINVDCx16_ASAP7_75t_R g1767 ( 
.A(n_1759),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1714),
.A2(n_1679),
.B1(n_1705),
.B2(n_1641),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1760),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1750),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1754),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1727),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1764),
.B(n_1643),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1712),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1740),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1735),
.B(n_1605),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1754),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1750),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1749),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1755),
.B(n_1641),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1607),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1752),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1713),
.B(n_1620),
.Y(n_1783)
);

INVxp67_ASAP7_75t_SL g1784 ( 
.A(n_1747),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1727),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1737),
.B(n_1613),
.Y(n_1786)
);

OA21x2_ASAP7_75t_L g1787 ( 
.A1(n_1738),
.A2(n_1664),
.B(n_1680),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1726),
.B(n_1607),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1753),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1753),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1727),
.Y(n_1791)
);

INVxp33_ASAP7_75t_L g1792 ( 
.A(n_1741),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1753),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1730),
.B(n_1717),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1731),
.B(n_1648),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1734),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1719),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1765),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1763),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1748),
.Y(n_1800)
);

INVxp67_ASAP7_75t_SL g1801 ( 
.A(n_1748),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1736),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1733),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1744),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1744),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1784),
.B(n_1744),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1784),
.B(n_1733),
.Y(n_1807)
);

OAI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1768),
.A2(n_1724),
.B1(n_1745),
.B2(n_1743),
.Y(n_1808)
);

AND2x2_ASAP7_75t_SL g1809 ( 
.A(n_1767),
.B(n_1724),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1797),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1803),
.B(n_1772),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1771),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1803),
.B(n_1733),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1775),
.Y(n_1814)
);

AOI322xp5_ASAP7_75t_L g1815 ( 
.A1(n_1767),
.A2(n_1723),
.A3(n_1714),
.B1(n_1732),
.B2(n_1715),
.C1(n_1721),
.C2(n_1728),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1775),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1770),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1797),
.Y(n_1818)
);

NAND4xp25_ASAP7_75t_L g1819 ( 
.A(n_1768),
.B(n_1751),
.C(n_1743),
.D(n_1766),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1785),
.B(n_1791),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1771),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1779),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1777),
.B(n_1761),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1770),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1770),
.Y(n_1825)
);

INVxp33_ASAP7_75t_L g1826 ( 
.A(n_1774),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1785),
.B(n_1738),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1802),
.A2(n_1745),
.B1(n_1678),
.B2(n_1746),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1778),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1799),
.B(n_1751),
.C(n_1746),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_SL g1831 ( 
.A(n_1802),
.B(n_1742),
.C(n_1762),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1776),
.B(n_1742),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1776),
.B(n_1716),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1800),
.A2(n_1759),
.B1(n_1722),
.B2(n_1718),
.C(n_1716),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1781),
.B(n_1718),
.Y(n_1835)
);

AO21x2_ASAP7_75t_L g1836 ( 
.A1(n_1801),
.A2(n_1790),
.B(n_1789),
.Y(n_1836)
);

INVx4_ASAP7_75t_L g1837 ( 
.A(n_1797),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1787),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1799),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1783),
.B(n_1614),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1787),
.Y(n_1841)
);

NOR2x1_ASAP7_75t_L g1842 ( 
.A(n_1796),
.B(n_1720),
.Y(n_1842)
);

BUFx3_ASAP7_75t_L g1843 ( 
.A(n_1787),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1804),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1843),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1810),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1823),
.Y(n_1847)
);

INVx4_ASAP7_75t_L g1848 ( 
.A(n_1818),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1814),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1807),
.B(n_1782),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1814),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1814),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1812),
.B(n_1783),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1813),
.B(n_1794),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1810),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1843),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1816),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1843),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1839),
.B(n_1725),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1812),
.B(n_1769),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1816),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1823),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1807),
.B(n_1782),
.Y(n_1863)
);

NAND2x1_ASAP7_75t_SL g1864 ( 
.A(n_1821),
.B(n_1807),
.Y(n_1864)
);

NOR2x1_ASAP7_75t_L g1865 ( 
.A(n_1818),
.B(n_1796),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1813),
.B(n_1788),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1813),
.B(n_1788),
.Y(n_1867)
);

NAND2x1_ASAP7_75t_L g1868 ( 
.A(n_1842),
.B(n_1796),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1821),
.B(n_1769),
.Y(n_1869)
);

AND2x2_ASAP7_75t_SL g1870 ( 
.A(n_1809),
.B(n_1795),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1810),
.B(n_1795),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1816),
.Y(n_1872)
);

INVx6_ASAP7_75t_L g1873 ( 
.A(n_1818),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1839),
.B(n_1773),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1822),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1810),
.B(n_1818),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1820),
.B(n_1794),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1822),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1811),
.B(n_1773),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1843),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1844),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1838),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1818),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1822),
.B(n_1780),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1811),
.B(n_1786),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1833),
.B(n_1798),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1838),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1844),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1838),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1877),
.B(n_1811),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1849),
.Y(n_1891)
);

NAND2x1p5_ASAP7_75t_L g1892 ( 
.A(n_1848),
.B(n_1809),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1849),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1873),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1859),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1845),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1851),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1864),
.A2(n_1806),
.B(n_1827),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1847),
.B(n_1832),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1874),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1877),
.B(n_1820),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1847),
.B(n_1832),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1851),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1852),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1845),
.Y(n_1905)
);

OAI21xp33_ASAP7_75t_L g1906 ( 
.A1(n_1864),
.A2(n_1806),
.B(n_1827),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1876),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1852),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1866),
.B(n_1820),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1862),
.B(n_1832),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1845),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1866),
.B(n_1827),
.Y(n_1912)
);

NAND2x1p5_ASAP7_75t_L g1913 ( 
.A(n_1848),
.B(n_1809),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1862),
.B(n_1806),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1857),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1857),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1874),
.B(n_1833),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1861),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_SL g1919 ( 
.A(n_1870),
.B(n_1809),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1886),
.B(n_1833),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1861),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1886),
.B(n_1835),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1866),
.B(n_1818),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1856),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1872),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.B(n_1837),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1886),
.B(n_1835),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1860),
.B(n_1835),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1860),
.B(n_1830),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1869),
.B(n_1830),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1871),
.B(n_1837),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1872),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1867),
.B(n_1837),
.Y(n_1933)
);

NAND2x1_ASAP7_75t_L g1934 ( 
.A(n_1873),
.B(n_1871),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1875),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1875),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1892),
.B(n_1871),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1892),
.B(n_1871),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1929),
.B(n_1850),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1892),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1913),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1930),
.B(n_1850),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1913),
.B(n_1876),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1900),
.B(n_1850),
.Y(n_1944)
);

AND2x2_ASAP7_75t_SL g1945 ( 
.A(n_1919),
.B(n_1870),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1899),
.B(n_1863),
.Y(n_1946)
);

NOR2x1p5_ASAP7_75t_L g1947 ( 
.A(n_1895),
.B(n_1831),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1891),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1913),
.B(n_1876),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1890),
.B(n_1876),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1895),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1891),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1893),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1902),
.B(n_1879),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1910),
.B(n_1881),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1914),
.B(n_1881),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1890),
.B(n_1846),
.Y(n_1957)
);

AOI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1898),
.A2(n_1906),
.B1(n_1808),
.B2(n_1880),
.C(n_1858),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1893),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1901),
.B(n_1846),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1907),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1896),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1901),
.B(n_1855),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1897),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1920),
.B(n_1863),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1922),
.B(n_1879),
.Y(n_1966)
);

AO22x1_ASAP7_75t_L g1967 ( 
.A1(n_1912),
.A2(n_1757),
.B1(n_1888),
.B2(n_1856),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1897),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1903),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1927),
.B(n_1917),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1903),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1928),
.B(n_1869),
.Y(n_1972)
);

INVx4_ASAP7_75t_L g1973 ( 
.A(n_1907),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1909),
.B(n_1855),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1904),
.B(n_1888),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1951),
.B(n_1934),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1951),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1958),
.A2(n_1939),
.B1(n_1942),
.B2(n_1815),
.C(n_1841),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1947),
.A2(n_1870),
.B1(n_1808),
.B2(n_1828),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1948),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1961),
.B(n_1912),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1947),
.A2(n_1828),
.B1(n_1834),
.B2(n_1873),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1948),
.Y(n_1983)
);

OAI32xp33_ASAP7_75t_L g1984 ( 
.A1(n_1944),
.A2(n_1856),
.A3(n_1858),
.B1(n_1880),
.B2(n_1853),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1945),
.B(n_1931),
.Y(n_1985)
);

OAI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1946),
.A2(n_1819),
.B1(n_1831),
.B2(n_1834),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1961),
.B(n_1909),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1945),
.A2(n_1836),
.B1(n_1880),
.B2(n_1858),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1957),
.B(n_1960),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1973),
.B(n_1970),
.Y(n_1990)
);

NOR3xp33_ASAP7_75t_L g1991 ( 
.A(n_1973),
.B(n_1819),
.C(n_1896),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1952),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1956),
.A2(n_1841),
.B1(n_1838),
.B2(n_1924),
.C(n_1911),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1940),
.A2(n_1841),
.B1(n_1804),
.B2(n_1805),
.Y(n_1994)
);

OAI21xp33_ASAP7_75t_L g1995 ( 
.A1(n_1957),
.A2(n_1926),
.B(n_1923),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1952),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1973),
.B(n_1967),
.C(n_1955),
.Y(n_1997)
);

OAI222xp33_ASAP7_75t_L g1998 ( 
.A1(n_1940),
.A2(n_1841),
.B1(n_1853),
.B2(n_1815),
.C1(n_1805),
.C2(n_1840),
.Y(n_1998)
);

OAI322xp33_ASAP7_75t_L g1999 ( 
.A1(n_1955),
.A2(n_1956),
.A3(n_1972),
.B1(n_1954),
.B2(n_1945),
.C1(n_1975),
.C2(n_1966),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1960),
.B(n_1931),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1953),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1963),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1953),
.Y(n_2003)
);

OAI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1940),
.A2(n_1815),
.B(n_1894),
.Y(n_2004)
);

INVxp33_ASAP7_75t_L g2005 ( 
.A(n_1989),
.Y(n_2005)
);

OAI211xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1991),
.A2(n_1997),
.B(n_1978),
.C(n_1976),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1977),
.B(n_1963),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1990),
.B(n_1973),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1981),
.B(n_1966),
.Y(n_2009)
);

O2A1O1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1979),
.A2(n_1998),
.B(n_1991),
.C(n_1999),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1987),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_1997),
.B(n_1941),
.C(n_1962),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1980),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1983),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_2000),
.Y(n_2015)
);

OAI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1988),
.A2(n_1982),
.B1(n_2004),
.B2(n_1993),
.C(n_1985),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_2002),
.B(n_1937),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1992),
.B(n_1954),
.Y(n_2018)
);

AOI21xp33_ASAP7_75t_SL g2019 ( 
.A1(n_1986),
.A2(n_1967),
.B(n_1894),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1996),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2001),
.B(n_1974),
.Y(n_2021)
);

AOI222xp33_ASAP7_75t_L g2022 ( 
.A1(n_1998),
.A2(n_1962),
.B1(n_1959),
.B2(n_1968),
.C1(n_1971),
.C2(n_1969),
.Y(n_2022)
);

NOR4xp25_ASAP7_75t_L g2023 ( 
.A(n_2003),
.B(n_1941),
.C(n_1962),
.D(n_1975),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1984),
.A2(n_1934),
.B(n_1943),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1995),
.Y(n_2025)
);

OAI31xp33_ASAP7_75t_L g2026 ( 
.A1(n_1994),
.A2(n_1941),
.A3(n_1938),
.B(n_1937),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1977),
.B(n_1974),
.Y(n_2027)
);

AOI221xp5_ASAP7_75t_L g2028 ( 
.A1(n_2010),
.A2(n_1959),
.B1(n_1971),
.B2(n_1969),
.C(n_1968),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_2022),
.B(n_1848),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2018),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_2022),
.A2(n_1964),
.B(n_1949),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2027),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_2023),
.A2(n_1964),
.B(n_1949),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_2027),
.B(n_1848),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_2005),
.B(n_1938),
.Y(n_2035)
);

XNOR2x2_ASAP7_75t_L g2036 ( 
.A(n_2012),
.B(n_1943),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2015),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2006),
.B(n_1883),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2007),
.Y(n_2039)
);

XOR2x2_ASAP7_75t_L g2040 ( 
.A(n_2016),
.B(n_1965),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2011),
.B(n_1972),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2009),
.Y(n_2042)
);

XNOR2x1_ASAP7_75t_L g2043 ( 
.A(n_2036),
.B(n_2011),
.Y(n_2043)
);

NAND4xp25_ASAP7_75t_L g2044 ( 
.A(n_2028),
.B(n_2008),
.C(n_2017),
.D(n_2025),
.Y(n_2044)
);

NOR3xp33_ASAP7_75t_L g2045 ( 
.A(n_2041),
.B(n_2019),
.C(n_2014),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2035),
.B(n_2021),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2032),
.Y(n_2047)
);

NAND4xp25_ASAP7_75t_L g2048 ( 
.A(n_2038),
.B(n_2024),
.C(n_2020),
.D(n_2013),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_2042),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_2041),
.B(n_1950),
.Y(n_2050)
);

NAND4xp25_ASAP7_75t_L g2051 ( 
.A(n_2031),
.B(n_2026),
.C(n_1950),
.D(n_1931),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2030),
.B(n_1923),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2037),
.B(n_1926),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_2039),
.B(n_1905),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2034),
.B(n_1873),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2040),
.B(n_1933),
.Y(n_2056)
);

OAI211xp5_ASAP7_75t_L g2057 ( 
.A1(n_2033),
.A2(n_1883),
.B(n_1837),
.C(n_1933),
.Y(n_2057)
);

OAI21xp33_ASAP7_75t_L g2058 ( 
.A1(n_2033),
.A2(n_1911),
.B(n_1905),
.Y(n_2058)
);

OAI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2043),
.A2(n_2029),
.B(n_1924),
.Y(n_2059)
);

OAI221xp5_ASAP7_75t_L g2060 ( 
.A1(n_2058),
.A2(n_1889),
.B1(n_1882),
.B2(n_1887),
.C(n_1873),
.Y(n_2060)
);

NAND4xp25_ASAP7_75t_L g2061 ( 
.A(n_2045),
.B(n_1665),
.C(n_1667),
.D(n_1837),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2050),
.B(n_1863),
.Y(n_2062)
);

AOI211xp5_ASAP7_75t_L g2063 ( 
.A1(n_2048),
.A2(n_1936),
.B(n_1935),
.C(n_1932),
.Y(n_2063)
);

AOI211xp5_ASAP7_75t_SL g2064 ( 
.A1(n_2047),
.A2(n_1908),
.B(n_1935),
.C(n_1932),
.Y(n_2064)
);

INVx1_ASAP7_75t_SL g2065 ( 
.A(n_2049),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2056),
.B(n_1854),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_2046),
.B(n_2044),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2065),
.Y(n_2068)
);

AOI322xp5_ASAP7_75t_L g2069 ( 
.A1(n_2067),
.A2(n_2053),
.A3(n_2052),
.B1(n_1887),
.B2(n_1889),
.C1(n_1882),
.C2(n_2055),
.Y(n_2069)
);

OAI21xp33_ASAP7_75t_L g2070 ( 
.A1(n_2061),
.A2(n_2051),
.B(n_2057),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2062),
.A2(n_2054),
.B1(n_1936),
.B2(n_1925),
.Y(n_2071)
);

AOI322xp5_ASAP7_75t_L g2072 ( 
.A1(n_2066),
.A2(n_1889),
.A3(n_1887),
.B1(n_1882),
.B2(n_1789),
.C1(n_1790),
.C2(n_1793),
.Y(n_2072)
);

AOI222xp33_ASAP7_75t_L g2073 ( 
.A1(n_2059),
.A2(n_1793),
.B1(n_1790),
.B2(n_1825),
.C1(n_1829),
.C2(n_1817),
.Y(n_2073)
);

OAI221xp5_ASAP7_75t_SL g2074 ( 
.A1(n_2063),
.A2(n_2060),
.B1(n_2064),
.B2(n_1885),
.C(n_1921),
.Y(n_2074)
);

AOI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2065),
.A2(n_1836),
.B1(n_1817),
.B2(n_1824),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2068),
.B(n_2070),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2069),
.B(n_1904),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_2074),
.B(n_2071),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2075),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_2073),
.B(n_1908),
.Y(n_2080)
);

XNOR2xp5_ASAP7_75t_L g2081 ( 
.A(n_2072),
.B(n_1706),
.Y(n_2081)
);

NAND3xp33_ASAP7_75t_SL g2082 ( 
.A(n_2076),
.B(n_1701),
.C(n_1885),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2077),
.Y(n_2083)
);

NOR2x1p5_ASAP7_75t_L g2084 ( 
.A(n_2079),
.B(n_1837),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2078),
.B(n_1915),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_2084),
.B(n_2085),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_2083),
.Y(n_2087)
);

OAI22x1_ASAP7_75t_L g2088 ( 
.A1(n_2087),
.A2(n_2081),
.B1(n_2080),
.B2(n_2082),
.Y(n_2088)
);

AOI221x1_ASAP7_75t_L g2089 ( 
.A1(n_2088),
.A2(n_2086),
.B1(n_1925),
.B2(n_1921),
.C(n_1918),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_2088),
.Y(n_2090)
);

AO22x1_ASAP7_75t_L g2091 ( 
.A1(n_2090),
.A2(n_2086),
.B1(n_1918),
.B2(n_1916),
.Y(n_2091)
);

AOI22x1_ASAP7_75t_L g2092 ( 
.A1(n_2089),
.A2(n_1916),
.B1(n_1915),
.B2(n_1758),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_2091),
.A2(n_1836),
.B(n_1884),
.Y(n_2093)
);

OAI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2092),
.A2(n_1829),
.B(n_1825),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2094),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_SL g2096 ( 
.A1(n_2095),
.A2(n_2093),
.B(n_1792),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2096),
.Y(n_2097)
);

OAI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_2097),
.A2(n_1729),
.B1(n_1865),
.B2(n_1868),
.C(n_1878),
.Y(n_2098)
);

AOI211xp5_ASAP7_75t_L g2099 ( 
.A1(n_2098),
.A2(n_1729),
.B(n_1756),
.C(n_1826),
.Y(n_2099)
);


endmodule