module fake_jpeg_7555_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_46),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_37),
.Y(n_62)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_15),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_32),
.Y(n_59)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_56),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_19),
.CON(n_54),
.SN(n_54)
);

OR2x2_ASAP7_75t_SL g112 ( 
.A(n_54),
.B(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_23),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_70),
.C(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_29),
.B1(n_18),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_76),
.B1(n_27),
.B2(n_49),
.Y(n_80)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_18),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_45),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_80),
.A2(n_81),
.B1(n_88),
.B2(n_90),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_93),
.Y(n_122)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_49),
.B1(n_25),
.B2(n_26),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_87),
.A2(n_98),
.B1(n_117),
.B2(n_93),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_42),
.B1(n_37),
.B2(n_17),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_37),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_99),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_42),
.B1(n_17),
.B2(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_107),
.B1(n_109),
.B2(n_63),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_13),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_102),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_44),
.B(n_33),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_78),
.C(n_1),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_26),
.B1(n_16),
.B2(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_10),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_43),
.B1(n_33),
.B2(n_39),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_0),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_115),
.B1(n_9),
.B2(n_2),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_44),
.B1(n_45),
.B2(n_39),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_116),
.B1(n_85),
.B2(n_82),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_55),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_64),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_58),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_116),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_15),
.B1(n_14),
.B2(n_11),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_121),
.B1(n_123),
.B2(n_127),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_74),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_66),
.B1(n_62),
.B2(n_40),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_62),
.B1(n_40),
.B2(n_72),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_135),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_131),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_2),
.B(n_4),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_146),
.B1(n_147),
.B2(n_116),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_127),
.B1(n_118),
.B2(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_143),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_1),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_94),
.B(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_149),
.A2(n_162),
.B(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_139),
.A2(n_81),
.B1(n_112),
.B2(n_80),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_156),
.B1(n_164),
.B2(n_168),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_158),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_147),
.B1(n_143),
.B2(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_89),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_99),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_161),
.B(n_178),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_99),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_109),
.B(n_89),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_102),
.B1(n_104),
.B2(n_101),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_95),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_107),
.B1(n_92),
.B2(n_101),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_172),
.B1(n_176),
.B2(n_182),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_113),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_173),
.B(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_82),
.B1(n_83),
.B2(n_95),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_108),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_114),
.C(n_96),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_130),
.C(n_138),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_91),
.B1(n_100),
.B2(n_86),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_119),
.A2(n_114),
.B(n_96),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_130),
.B1(n_128),
.B2(n_135),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_149),
.Y(n_232)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_194),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_208),
.B(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_141),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_197),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_206),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_133),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_161),
.C(n_175),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_161),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_133),
.A3(n_141),
.B1(n_138),
.B2(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_203),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_151),
.A2(n_138),
.B1(n_132),
.B2(n_91),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_204),
.B1(n_214),
.B2(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_150),
.A2(n_168),
.B1(n_151),
.B2(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_155),
.A2(n_4),
.B(n_5),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_162),
.A2(n_132),
.B1(n_100),
.B2(n_86),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_198),
.C(n_188),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_188),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_224),
.B1(n_238),
.B2(n_240),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_178),
.B1(n_158),
.B2(n_171),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_235),
.B(n_159),
.Y(n_253)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_228),
.B1(n_183),
.B2(n_204),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_191),
.B1(n_214),
.B2(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_241),
.C(n_149),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_161),
.B(n_159),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_265),
.C(n_266),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_249),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_211),
.B(n_208),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_252),
.B(n_253),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_233),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_205),
.B1(n_187),
.B2(n_189),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_258),
.B1(n_244),
.B2(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_262),
.B1(n_229),
.B2(n_238),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g258 ( 
.A1(n_223),
.A2(n_199),
.B1(n_211),
.B2(n_191),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_183),
.CI(n_213),
.CON(n_261),
.SN(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_225),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_237),
.A2(n_215),
.B1(n_203),
.B2(n_173),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_195),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_260),
.B1(n_226),
.B2(n_258),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_232),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_274),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_234),
.B1(n_217),
.B2(n_240),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_273),
.B1(n_278),
.B2(n_280),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_216),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_216),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_261),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_281),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_217),
.B1(n_242),
.B2(n_243),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_220),
.C(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_257),
.C(n_197),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_231),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_227),
.B1(n_225),
.B2(n_218),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_171),
.B1(n_153),
.B2(n_212),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_181),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_154),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_248),
.CI(n_261),
.CON(n_287),
.SN(n_287)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_287),
.B(n_271),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_262),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_289),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_296),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_294),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_251),
.B1(n_264),
.B2(n_248),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_300),
.B1(n_270),
.B2(n_284),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_218),
.C(n_224),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_153),
.B1(n_86),
.B2(n_154),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_4),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_5),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_283),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_310),
.B1(n_290),
.B2(n_296),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_269),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_311),
.C(n_292),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_278),
.B(n_268),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_4),
.C(n_5),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_320),
.B(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_293),
.C(n_286),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_289),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_309),
.CI(n_303),
.CON(n_322),
.SN(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_303),
.Y(n_324)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_320),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_286),
.B(n_7),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_6),
.B1(n_8),
.B2(n_315),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_324),
.C(n_326),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_332),
.C(n_334),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_336),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_333),
.B(n_6),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);


endmodule