module fake_jpeg_3526_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_57),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_35),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_59),
.B(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_40),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_67),
.Y(n_70)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_30),
.B(n_3),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_2),
.C(n_6),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_30),
.A3(n_26),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_3),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.C(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_9),
.C(n_10),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_65),
.B1(n_61),
.B2(n_11),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_12),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_76),
.C(n_75),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_80),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_73),
.A3(n_69),
.B1(n_16),
.B2(n_18),
.C1(n_19),
.C2(n_14),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_15),
.CI(n_21),
.CON(n_85),
.SN(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_22),
.Y(n_86)
);


endmodule