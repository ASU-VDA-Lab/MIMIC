module fake_aes_3108_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx1_ASAP7_75t_SL g4 ( .A(n_0), .Y(n_4) );
NAND3xp33_ASAP7_75t_L g5 ( .A(n_3), .B(n_4), .C(n_0), .Y(n_5) );
NOR2x1_ASAP7_75t_R g6 ( .A(n_3), .B(n_0), .Y(n_6) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx3_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
OAI221xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_6), .B1(n_1), .B2(n_2), .C(n_0), .Y(n_9) );
OA211x2_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_1), .B(n_2), .C(n_8), .Y(n_10) );
OAI22xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_2), .B1(n_8), .B2(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
endmodule