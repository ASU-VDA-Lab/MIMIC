module fake_netlist_6_924_n_5262 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5262);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5262;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_5229;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_695;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_4062;
wire n_3902;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_1077;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_4598;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3777;
wire n_4203;
wire n_3641;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4145;
wire n_3121;
wire n_4821;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_1266;
wire n_709;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3910;
wire n_3812;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_697;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1475;
wire n_716;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2969;
wire n_2787;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_641),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_89),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_68),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_642),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_483),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_160),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_541),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_427),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_123),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_171),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_161),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_181),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_443),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_544),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_600),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_424),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_524),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_293),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_305),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_145),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_667),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_497),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_496),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_417),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_197),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_484),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_520),
.Y(n_720)
);

CKINVDCx16_ASAP7_75t_R g721 ( 
.A(n_541),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_431),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_208),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_66),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_460),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_687),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_635),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_663),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_250),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_15),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_660),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_354),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_25),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_78),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_381),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_168),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_583),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_687),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_78),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_683),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_145),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_672),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_251),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_676),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_184),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_225),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_43),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_592),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_312),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_249),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_522),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_634),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_354),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_161),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_539),
.Y(n_755)
);

CKINVDCx16_ASAP7_75t_R g756 ( 
.A(n_545),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_239),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_33),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_615),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_325),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_60),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_351),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_562),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_270),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_336),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_204),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_538),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_575),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_33),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_92),
.Y(n_770)
);

CKINVDCx14_ASAP7_75t_R g771 ( 
.A(n_73),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_623),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_673),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_568),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_289),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_603),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_596),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_310),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_65),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_273),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_605),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_291),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_664),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_162),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_320),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_542),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_607),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_190),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_630),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_540),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_353),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_493),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_309),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_632),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_564),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_163),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_574),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_442),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_669),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_666),
.Y(n_800)
);

CKINVDCx14_ASAP7_75t_R g801 ( 
.A(n_238),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_55),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_85),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_114),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_236),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_543),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_329),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_488),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_604),
.Y(n_809)
);

BUFx5_ASAP7_75t_L g810 ( 
.A(n_257),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_86),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_666),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_583),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_399),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_97),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_120),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_473),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_101),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_21),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_602),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_12),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_314),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_76),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_191),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_430),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_383),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_134),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_18),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_110),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_123),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_692),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_562),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_20),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_515),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_68),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_548),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_309),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_665),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_614),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_68),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_514),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_415),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_123),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_597),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_13),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_61),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_206),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_311),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_405),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_501),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_185),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_50),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_333),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_691),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_84),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_481),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_203),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_97),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_501),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_175),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_250),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_504),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_508),
.Y(n_863)
);

CKINVDCx16_ASAP7_75t_R g864 ( 
.A(n_609),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_477),
.Y(n_865)
);

BUFx5_ASAP7_75t_L g866 ( 
.A(n_559),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_653),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_163),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_603),
.Y(n_869)
);

BUFx5_ASAP7_75t_L g870 ( 
.A(n_351),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_537),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_325),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_516),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_378),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_446),
.Y(n_875)
);

BUFx5_ASAP7_75t_L g876 ( 
.A(n_330),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_121),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_441),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_133),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_288),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_14),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_56),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_445),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_632),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_533),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_101),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_503),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_154),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_91),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_436),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_417),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_479),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_598),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_189),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_331),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_442),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_490),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_80),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_502),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_491),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_674),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_534),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_480),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_70),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_242),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_340),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_487),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_686),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_410),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_504),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_629),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_368),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_681),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_176),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_75),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_216),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_91),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_226),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_670),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_193),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_106),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_387),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_386),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_359),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_627),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_286),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_547),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_311),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_79),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_256),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_380),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_162),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_160),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_241),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_308),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_387),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_334),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_208),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_576),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_549),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_513),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_447),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_674),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_404),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_41),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_187),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_112),
.Y(n_947)
);

BUFx10_ASAP7_75t_L g948 ( 
.A(n_490),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_518),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_423),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_389),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_395),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_525),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_51),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_124),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_128),
.Y(n_956)
);

CKINVDCx16_ASAP7_75t_R g957 ( 
.A(n_86),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_668),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_58),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_670),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_688),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_491),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_308),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_130),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_129),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_287),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_408),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_193),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_564),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_427),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_559),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_197),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_594),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_397),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_317),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_378),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_435),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_148),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_622),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_2),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_594),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_642),
.Y(n_982)
);

BUFx10_ASAP7_75t_L g983 ( 
.A(n_67),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_36),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_337),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_407),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_384),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_327),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_404),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_396),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_131),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_129),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_234),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_269),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_113),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_576),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_675),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_32),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_676),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_597),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_261),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_187),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_225),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_246),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_191),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_650),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_28),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_390),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_407),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_395),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_167),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_485),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_350),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_671),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_143),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_455),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_248),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_358),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_11),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_152),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_103),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_437),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_41),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_10),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_369),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_645),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_422),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_20),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_5),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_771),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_810),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_957),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_801),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_810),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_802),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_721),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_756),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_838),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_810),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_864),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_930),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_810),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_700),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_694),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_759),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_810),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_810),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_763),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_702),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_765),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_810),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_772),
.Y(n_1052)
);

BUFx5_ASAP7_75t_L g1053 ( 
.A(n_697),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_810),
.Y(n_1054)
);

BUFx5_ASAP7_75t_L g1055 ( 
.A(n_698),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_866),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_866),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_774),
.Y(n_1058)
);

INVxp33_ASAP7_75t_L g1059 ( 
.A(n_846),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_776),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_866),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_777),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_866),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_866),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_866),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_778),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_998),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_866),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_784),
.Y(n_1069)
);

CKINVDCx16_ASAP7_75t_R g1070 ( 
.A(n_702),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_787),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_735),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_866),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_790),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_870),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_870),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_870),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_769),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_791),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_870),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_769),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_794),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_795),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_870),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_816),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_870),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_870),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_796),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_870),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_798),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_876),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_L g1092 ( 
.A(n_872),
.B(n_0),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_769),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_700),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_876),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_876),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_799),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_876),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_876),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_876),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_876),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_876),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_769),
.Y(n_1103)
);

INVxp33_ASAP7_75t_L g1104 ( 
.A(n_818),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_769),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_806),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_882),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_882),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_807),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_808),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_750),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_695),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_882),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_882),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_882),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_998),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_724),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_696),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_734),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_745),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_747),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_702),
.Y(n_1122)
);

BUFx5_ASAP7_75t_L g1123 ( 
.A(n_712),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_758),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_779),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_715),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_761),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_770),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_803),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_811),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_815),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_804),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_835),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_819),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_852),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_855),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_881),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_821),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_886),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_889),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_917),
.Y(n_1141)
);

INVxp33_ASAP7_75t_L g1142 ( 
.A(n_947),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_828),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_879),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_700),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_700),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_733),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_700),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_829),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_954),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_753),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_896),
.B(n_0),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_830),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_733),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_959),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_840),
.Y(n_1156)
);

CKINVDCx16_ASAP7_75t_R g1157 ( 
.A(n_983),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_715),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_984),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_843),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1007),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1024),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_845),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_722),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_722),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_730),
.B(n_1),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_766),
.Y(n_1167)
);

INVxp33_ASAP7_75t_L g1168 ( 
.A(n_1011),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_757),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_766),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_858),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_980),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_783),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_736),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_783),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_736),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_849),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_877),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_849),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_865),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_898),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_865),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_958),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_736),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_958),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_962),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_962),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_904),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1008),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1008),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_823),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_736),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_983),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_736),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_788),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_764),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_788),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_921),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_788),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_767),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_788),
.Y(n_1201)
);

BUFx5_ASAP7_75t_L g1202 ( 
.A(n_714),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_788),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_834),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_834),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_834),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_929),
.Y(n_1207)
);

CKINVDCx14_ASAP7_75t_R g1208 ( 
.A(n_983),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_834),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_834),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_994),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_994),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_994),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_994),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_980),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_703),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_994),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1026),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1026),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_792),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_945),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1029),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_995),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1026),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1026),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_854),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1026),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_812),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_820),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_824),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_825),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_826),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1023),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1023),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_827),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_719),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_726),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_841),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_727),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_842),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_729),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_738),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_737),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_742),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_844),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_738),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_847),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_850),
.Y(n_1248)
);

BUFx8_ASAP7_75t_SL g1249 ( 
.A(n_833),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_853),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_856),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_746),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_703),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_751),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_703),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_995),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_875),
.B(n_912),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_751),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_760),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_887),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_859),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_768),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_888),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_861),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_773),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_775),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_781),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_863),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_782),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_867),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_785),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_786),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_789),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_760),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_869),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_793),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_871),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_797),
.Y(n_1278)
);

BUFx10_ASAP7_75t_L g1279 ( 
.A(n_1019),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_800),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_874),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_813),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_814),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_832),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_837),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_857),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_878),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_860),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_875),
.B(n_0),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_805),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_880),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_868),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_884),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_805),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_890),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_873),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_831),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_883),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_915),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_831),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_891),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_894),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_885),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_892),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_893),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_895),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_899),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_903),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_926),
.Y(n_1309)
);

BUFx5_ASAP7_75t_L g1310 ( 
.A(n_916),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_920),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_836),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_897),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_836),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_900),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_901),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_924),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_925),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_713),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_902),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_713),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_905),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_906),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_931),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_908),
.Y(n_1325)
);

CKINVDCx16_ASAP7_75t_R g1326 ( 
.A(n_713),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_935),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_910),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_936),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_848),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_822),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_848),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_911),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_939),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_940),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_970),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_941),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_913),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_914),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_942),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1019),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1016),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_943),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_918),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_964),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1021),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_964),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_919),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_922),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_951),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_952),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_953),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_822),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_976),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_956),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_960),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_923),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_965),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_927),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_928),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_967),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_932),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_822),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_976),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_969),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_933),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_972),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_991),
.Y(n_1368)
);

INVxp33_ASAP7_75t_L g1369 ( 
.A(n_991),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_973),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_974),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1021),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_975),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_982),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_985),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_987),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_989),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1028),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_934),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1000),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_937),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1028),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_938),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_944),
.Y(n_1384)
);

CKINVDCx16_ASAP7_75t_R g1385 ( 
.A(n_851),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1004),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1005),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1014),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_946),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1018),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1020),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_912),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_949),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_739),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1033),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1078),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1030),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1072),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1081),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1072),
.Y(n_1400)
);

INVxp67_ASAP7_75t_SL g1401 ( 
.A(n_1093),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1111),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1103),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1111),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1107),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1228),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1151),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1108),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_1037),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1151),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1169),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1113),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1229),
.B(n_950),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1230),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1067),
.B(n_955),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1231),
.Y(n_1416)
);

CKINVDCx16_ASAP7_75t_R g1417 ( 
.A(n_1208),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1036),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1114),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1126),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1232),
.B(n_699),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1235),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1115),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1238),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1240),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1245),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1038),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1192),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1199),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_L g1430 ( 
.A(n_1247),
.B(n_1),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1169),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1196),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1302),
.Y(n_1433)
);

CKINVDCx14_ASAP7_75t_R g1434 ( 
.A(n_1032),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1248),
.B(n_699),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1126),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1201),
.Y(n_1437)
);

INVxp67_ASAP7_75t_SL g1438 ( 
.A(n_1158),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1203),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1383),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1204),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1196),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1384),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1205),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1389),
.B(n_851),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1209),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1394),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1211),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1213),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1214),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1217),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1393),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1346),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1158),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1040),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1174),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1200),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1218),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1206),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1112),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1118),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1105),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1224),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1225),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1125),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1132),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1134),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1227),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1041),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1067),
.B(n_701),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1105),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1138),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1143),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1149),
.B(n_1153),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1219),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1219),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1294),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1147),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1200),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1312),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1043),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1041),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1043),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1035),
.B(n_704),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1043),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1220),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1156),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1160),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1163),
.B(n_701),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1327),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1094),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1094),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1336),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1171),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1094),
.Y(n_1495)
);

NOR2xp67_ASAP7_75t_L g1496 ( 
.A(n_1178),
.B(n_1),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1195),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1181),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1174),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1195),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1195),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1145),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_L g1503 ( 
.A(n_1188),
.B(n_2),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1145),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1116),
.B(n_705),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1198),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1146),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1146),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1148),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1207),
.B(n_705),
.Y(n_1510)
);

CKINVDCx16_ASAP7_75t_R g1511 ( 
.A(n_1049),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1148),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1206),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1176),
.Y(n_1514)
);

CKINVDCx16_ASAP7_75t_R g1515 ( 
.A(n_1070),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1220),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1176),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1221),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1154),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1226),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1184),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1172),
.Y(n_1522)
);

XOR2xp5_ASAP7_75t_L g1523 ( 
.A(n_1226),
.B(n_706),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1184),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1206),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1222),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1194),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1044),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1044),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1194),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1045),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1260),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1197),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1197),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1045),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1116),
.B(n_706),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1048),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1210),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1048),
.Y(n_1539)
);

CKINVDCx16_ASAP7_75t_R g1540 ( 
.A(n_1122),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1210),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1370),
.B(n_1289),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1174),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1215),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1050),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1236),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1237),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1050),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1239),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1255),
.B(n_725),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1052),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1241),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1257),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1052),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1243),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1058),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1058),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_1249),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1191),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1253),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1223),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1244),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1260),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1263),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1252),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1262),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1265),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1060),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1266),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1164),
.B(n_707),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1256),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1267),
.Y(n_1572)
);

INVxp33_ASAP7_75t_SL g1573 ( 
.A(n_1152),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1269),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1165),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1263),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1060),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_L g1578 ( 
.A(n_1062),
.B(n_1066),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1271),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1062),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1066),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1069),
.Y(n_1582)
);

INVxp33_ASAP7_75t_L g1583 ( 
.A(n_1249),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1272),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1309),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1069),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1309),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1273),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1071),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1206),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1341),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1071),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1253),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1276),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1074),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1342),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1278),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1342),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1372),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1074),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1167),
.B(n_707),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1280),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1282),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1079),
.B(n_708),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1283),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1212),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1079),
.B(n_708),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1212),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1372),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1284),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1082),
.B(n_709),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1082),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1083),
.B(n_709),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1378),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1083),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1285),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1378),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1286),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1088),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1288),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1088),
.B(n_710),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1090),
.Y(n_1622)
);

CKINVDCx16_ASAP7_75t_R g1623 ( 
.A(n_1157),
.Y(n_1623)
);

CKINVDCx16_ASAP7_75t_R g1624 ( 
.A(n_1193),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1090),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1321),
.Y(n_1626)
);

INVxp33_ASAP7_75t_L g1627 ( 
.A(n_1104),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1097),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1382),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1097),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1292),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1382),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1296),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1298),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1104),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1106),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1321),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_1326),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1303),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1304),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1305),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1306),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1307),
.Y(n_1643)
);

CKINVDCx16_ASAP7_75t_R g1644 ( 
.A(n_1385),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1308),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1311),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1212),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1353),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1212),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1353),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1299),
.Y(n_1651)
);

CKINVDCx16_ASAP7_75t_R g1652 ( 
.A(n_1279),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1317),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1106),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1109),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1109),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1110),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_1110),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1318),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1324),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1250),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1329),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1334),
.Y(n_1663)
);

BUFx6f_ASAP7_75t_SL g1664 ( 
.A(n_1279),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1250),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1251),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1251),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1261),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1261),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1335),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1170),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1337),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1340),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1264),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1242),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1173),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1264),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1268),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_1268),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1085),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_1270),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1343),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1270),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1275),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1242),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1350),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1351),
.Y(n_1687)
);

CKINVDCx16_ASAP7_75t_R g1688 ( 
.A(n_1279),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1275),
.B(n_710),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1255),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1277),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1277),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1281),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1352),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1281),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1355),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1356),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1242),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1287),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1331),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1459),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1475),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1462),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1476),
.B(n_1246),
.Y(n_1704)
);

AND2x6_ASAP7_75t_L g1705 ( 
.A(n_1542),
.B(n_1031),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1420),
.B(n_1246),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1447),
.B(n_1369),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1459),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1459),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1481),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1559),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1459),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1456),
.B(n_1034),
.Y(n_1713)
);

INVx6_ASAP7_75t_L g1714 ( 
.A(n_1542),
.Y(n_1714)
);

BUFx8_ASAP7_75t_L g1715 ( 
.A(n_1664),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1647),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_L g1717 ( 
.A(n_1415),
.B(n_1053),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1647),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1462),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1553),
.B(n_1542),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1664),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1502),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1647),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1483),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1456),
.B(n_1039),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1399),
.B(n_1046),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1675),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1651),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1401),
.B(n_1047),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1504),
.Y(n_1730)
);

NOR2x1_ASAP7_75t_L g1731 ( 
.A(n_1499),
.B(n_1578),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1690),
.B(n_1287),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1396),
.B(n_1054),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1575),
.B(n_1369),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1513),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1507),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1546),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1513),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1436),
.B(n_1056),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1438),
.B(n_1254),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1573),
.B(n_1291),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1547),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1454),
.B(n_1057),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1485),
.A2(n_1063),
.B(n_1061),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1508),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1543),
.A2(n_1051),
.B(n_1042),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1575),
.B(n_1254),
.Y(n_1747)
);

BUFx12f_ASAP7_75t_L g1748 ( 
.A(n_1455),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1491),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1525),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1509),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1492),
.A2(n_1065),
.B(n_1064),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1499),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1477),
.B(n_1068),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1671),
.B(n_1258),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1573),
.B(n_1291),
.Y(n_1756)
);

OA21x2_ASAP7_75t_L g1757 ( 
.A1(n_1495),
.A2(n_1075),
.B(n_1073),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1484),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1671),
.Y(n_1759)
);

BUFx8_ASAP7_75t_SL g1760 ( 
.A(n_1398),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1525),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1512),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1514),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1590),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1676),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1676),
.B(n_1258),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1489),
.B(n_1293),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1433),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1474),
.B(n_1076),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1517),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1497),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1675),
.B(n_1274),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1521),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1500),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1480),
.B(n_1077),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1501),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1403),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1524),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1428),
.A2(n_1087),
.B(n_1080),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1429),
.A2(n_1091),
.B(n_1089),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1527),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1490),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1405),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1408),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1412),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1437),
.A2(n_1096),
.B(n_1095),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1510),
.B(n_1293),
.Y(n_1787)
);

OAI22x1_ASAP7_75t_SL g1788 ( 
.A1(n_1599),
.A2(n_716),
.B1(n_717),
.B2(n_711),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1549),
.A2(n_1142),
.B1(n_1168),
.B2(n_1144),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1530),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1590),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1685),
.B(n_1098),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1606),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1685),
.B(n_1099),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1606),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1533),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1608),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1523),
.A2(n_1651),
.B1(n_1657),
.B2(n_1655),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1698),
.B(n_1100),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1608),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1552),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1649),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1698),
.B(n_1274),
.Y(n_1803)
);

INVx4_ASAP7_75t_L g1804 ( 
.A(n_1649),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1555),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1562),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1421),
.B(n_1295),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1565),
.B(n_1297),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1423),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1604),
.A2(n_1301),
.B1(n_1313),
.B2(n_1295),
.Y(n_1811)
);

BUFx12f_ASAP7_75t_L g1812 ( 
.A(n_1455),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1439),
.B(n_1101),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1534),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1538),
.Y(n_1815)
);

INVx5_ASAP7_75t_L g1816 ( 
.A(n_1445),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1441),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1444),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1446),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1448),
.A2(n_1102),
.B(n_1449),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1550),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1566),
.B(n_1297),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1435),
.B(n_1301),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1450),
.Y(n_1824)
);

AND2x2_ASAP7_75t_SL g1825 ( 
.A(n_1607),
.B(n_1166),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1541),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1611),
.B(n_1313),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1451),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1458),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1471),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1463),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1464),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1468),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1567),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1569),
.B(n_1300),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1613),
.A2(n_1316),
.B1(n_1320),
.B2(n_1315),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1560),
.B(n_1053),
.Y(n_1837)
);

CKINVDCx16_ASAP7_75t_R g1838 ( 
.A(n_1417),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_L g1839 ( 
.A(n_1621),
.B(n_1175),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1493),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1572),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1574),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1579),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1689),
.A2(n_1316),
.B1(n_1320),
.B2(n_1315),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1584),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1398),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1588),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1594),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1597),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1602),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1680),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1603),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1605),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1610),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1478),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1616),
.Y(n_1856)
);

AND2x2_ASAP7_75t_SL g1857 ( 
.A(n_1539),
.B(n_1242),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1618),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1620),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1627),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1635),
.B(n_1300),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1631),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1655),
.A2(n_716),
.B1(n_717),
.B2(n_711),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1633),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1634),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1593),
.B(n_1053),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1639),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1640),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1664),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1641),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1642),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1643),
.Y(n_1872)
);

OAI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1570),
.A2(n_1051),
.B(n_1042),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1645),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1646),
.Y(n_1875)
);

AND2x6_ASAP7_75t_L g1876 ( 
.A(n_1653),
.B(n_1084),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1659),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1601),
.A2(n_1086),
.B(n_1084),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1700),
.B(n_1314),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1648),
.B(n_1053),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1660),
.Y(n_1881)
);

OA21x2_ASAP7_75t_L g1882 ( 
.A1(n_1662),
.A2(n_1086),
.B(n_1314),
.Y(n_1882)
);

CKINVDCx8_ASAP7_75t_R g1883 ( 
.A(n_1409),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1663),
.Y(n_1884)
);

INVx6_ASAP7_75t_L g1885 ( 
.A(n_1652),
.Y(n_1885)
);

OA21x2_ASAP7_75t_L g1886 ( 
.A1(n_1670),
.A2(n_1345),
.B(n_1332),
.Y(n_1886)
);

INVx6_ASAP7_75t_L g1887 ( 
.A(n_1688),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1672),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1650),
.B(n_1053),
.Y(n_1889)
);

OA21x2_ASAP7_75t_L g1890 ( 
.A1(n_1673),
.A2(n_1345),
.B(n_1332),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1682),
.B(n_1347),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1686),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1626),
.B(n_1053),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1687),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1694),
.B(n_1347),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1696),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1697),
.Y(n_1897)
);

OA21x2_ASAP7_75t_L g1898 ( 
.A1(n_1470),
.A2(n_1536),
.B(n_1505),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1496),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1453),
.B(n_1322),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1503),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1637),
.Y(n_1902)
);

BUFx12f_ASAP7_75t_L g1903 ( 
.A(n_1397),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1519),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1430),
.B(n_1358),
.Y(n_1905)
);

OA21x2_ASAP7_75t_L g1906 ( 
.A1(n_1522),
.A2(n_1179),
.B(n_1177),
.Y(n_1906)
);

OAI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1506),
.A2(n_1182),
.B(n_1180),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1518),
.A2(n_1185),
.B(n_1183),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1544),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1545),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1561),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1683),
.B(n_1053),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1571),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1434),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1591),
.B(n_1392),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1615),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1622),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1414),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1406),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1422),
.A2(n_1323),
.B1(n_1325),
.B2(n_1322),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_L g1921 ( 
.A1(n_1469),
.A2(n_1187),
.B(n_1186),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1482),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1418),
.B(n_1361),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1424),
.B(n_1323),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_SL g1925 ( 
.A1(n_1657),
.A2(n_720),
.B1(n_723),
.B2(n_718),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1425),
.A2(n_1328),
.B1(n_1333),
.B2(n_1325),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1460),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1426),
.A2(n_1333),
.B1(n_1338),
.B2(n_1328),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1414),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1461),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1465),
.B(n_1055),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1466),
.B(n_1338),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1467),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1472),
.B(n_1055),
.Y(n_1934)
);

BUFx8_ASAP7_75t_L g1935 ( 
.A(n_1511),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1473),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1487),
.B(n_1055),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1488),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1494),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1498),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1526),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1416),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1416),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1427),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1440),
.B(n_1055),
.Y(n_1945)
);

XNOR2x2_ASAP7_75t_L g1946 ( 
.A(n_1599),
.B(n_762),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1440),
.B(n_1392),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1443),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1443),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1452),
.A2(n_1190),
.B(n_1189),
.Y(n_1950)
);

INVx4_ASAP7_75t_L g1951 ( 
.A(n_1452),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1528),
.B(n_1055),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1529),
.B(n_1055),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1531),
.B(n_1055),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1535),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1537),
.B(n_1123),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1548),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1551),
.B(n_1365),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1554),
.Y(n_1959)
);

OA21x2_ASAP7_75t_L g1960 ( 
.A1(n_1600),
.A2(n_1234),
.B(n_1233),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1395),
.A2(n_1344),
.B1(n_1348),
.B2(n_1339),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1600),
.B(n_1339),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1556),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1557),
.B(n_1344),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1397),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1568),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1577),
.B(n_1348),
.Y(n_1967)
);

OA21x2_ASAP7_75t_L g1968 ( 
.A1(n_1612),
.A2(n_1371),
.B(n_1367),
.Y(n_1968)
);

OA21x2_ASAP7_75t_L g1969 ( 
.A1(n_1612),
.A2(n_1374),
.B(n_1373),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1580),
.B(n_1392),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1581),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1582),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1586),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1589),
.B(n_1375),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_SL g1975 ( 
.A1(n_1658),
.A2(n_720),
.B1(n_723),
.B2(n_718),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1592),
.B(n_1349),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1595),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1665),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1619),
.B(n_1349),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1666),
.A2(n_1377),
.B(n_1376),
.Y(n_1980)
);

OA21x2_ASAP7_75t_L g1981 ( 
.A1(n_1619),
.A2(n_1386),
.B(n_1380),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1674),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1677),
.B(n_1392),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1691),
.B(n_1123),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1692),
.B(n_1123),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1695),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1658),
.A2(n_1661),
.B1(n_1668),
.B2(n_1667),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1625),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1625),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1714),
.A2(n_1630),
.B1(n_1636),
.B2(n_1628),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1714),
.A2(n_1654),
.B1(n_1628),
.B2(n_1636),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1707),
.B(n_1142),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1707),
.B(n_1768),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1719),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1840),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1734),
.B(n_1331),
.Y(n_1996)
);

AO22x2_ASAP7_75t_L g1997 ( 
.A1(n_1989),
.A2(n_1363),
.B1(n_809),
.B2(n_817),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1886),
.Y(n_1998)
);

AO22x2_ASAP7_75t_L g1999 ( 
.A1(n_1989),
.A2(n_1363),
.B1(n_839),
.B2(n_907),
.Y(n_1999)
);

AO22x2_ASAP7_75t_L g2000 ( 
.A1(n_1821),
.A2(n_909),
.B1(n_992),
.B2(n_780),
.Y(n_2000)
);

OAI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1714),
.A2(n_1654),
.B1(n_1656),
.B2(n_1630),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1719),
.Y(n_2002)
);

AO22x2_ASAP7_75t_L g2003 ( 
.A1(n_1821),
.A2(n_1009),
.B1(n_1022),
.B2(n_1006),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1714),
.Y(n_2004)
);

OA22x2_ASAP7_75t_L g2005 ( 
.A1(n_1863),
.A2(n_1319),
.B1(n_1216),
.B2(n_1656),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1734),
.B(n_1357),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1912),
.A2(n_1168),
.B1(n_1359),
.B2(n_1357),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1886),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1720),
.B(n_1359),
.Y(n_2009)
);

OR2x6_ASAP7_75t_L g2010 ( 
.A(n_1840),
.B(n_1092),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1886),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1827),
.B(n_1395),
.Y(n_2012)
);

AO22x2_ASAP7_75t_L g2013 ( 
.A1(n_1988),
.A2(n_1388),
.B1(n_1390),
.B2(n_1387),
.Y(n_2013)
);

OAI22xp33_ASAP7_75t_SL g2014 ( 
.A1(n_1899),
.A2(n_1362),
.B1(n_1366),
.B2(n_1360),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1719),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1861),
.B(n_1360),
.Y(n_2016)
);

OAI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1758),
.A2(n_1362),
.B1(n_1379),
.B2(n_1366),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1825),
.A2(n_1381),
.B1(n_1379),
.B2(n_1661),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1703),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1825),
.A2(n_1381),
.B1(n_1668),
.B2(n_1667),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1703),
.Y(n_2021)
);

OAI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1808),
.A2(n_1059),
.B1(n_1644),
.B2(n_1540),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1720),
.A2(n_1678),
.B1(n_1679),
.B2(n_1669),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1890),
.Y(n_2024)
);

AO22x1_ASAP7_75t_SL g2025 ( 
.A1(n_1946),
.A2(n_1917),
.B1(n_1910),
.B2(n_1949),
.Y(n_2025)
);

OAI22xp33_ASAP7_75t_SL g2026 ( 
.A1(n_1901),
.A2(n_731),
.B1(n_732),
.B2(n_728),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1711),
.Y(n_2027)
);

OAI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1816),
.A2(n_1059),
.B1(n_1623),
.B2(n_1515),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1861),
.B(n_1624),
.Y(n_2029)
);

AO22x2_ASAP7_75t_L g2030 ( 
.A1(n_1988),
.A2(n_1391),
.B1(n_948),
.B2(n_851),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1772),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1860),
.B(n_1558),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1782),
.B(n_1120),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1772),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1772),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1857),
.B(n_1669),
.Y(n_2036)
);

OAI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1816),
.A2(n_731),
.B1(n_732),
.B2(n_728),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1767),
.B(n_1678),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1726),
.B(n_1123),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1857),
.A2(n_1681),
.B1(n_1684),
.B2(n_1679),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1960),
.A2(n_1684),
.B1(n_1693),
.B2(n_1681),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1890),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1787),
.B(n_1693),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1947),
.B(n_1120),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1947),
.B(n_1120),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1890),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1882),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1759),
.B(n_1117),
.Y(n_2048)
);

OAI22xp33_ASAP7_75t_SL g2049 ( 
.A1(n_1945),
.A2(n_741),
.B1(n_743),
.B2(n_740),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1918),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_SL g2051 ( 
.A1(n_1846),
.A2(n_1614),
.B1(n_1617),
.B2(n_1609),
.Y(n_2051)
);

OR2x6_ASAP7_75t_L g2052 ( 
.A(n_1938),
.B(n_1119),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1803),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1970),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1960),
.A2(n_1699),
.B1(n_1123),
.B2(n_1310),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1911),
.B(n_1583),
.Y(n_2056)
);

AO22x2_ASAP7_75t_L g2057 ( 
.A1(n_1949),
.A2(n_948),
.B1(n_1124),
.B2(n_1121),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1803),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1960),
.A2(n_1898),
.B1(n_1769),
.B2(n_1705),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1970),
.B(n_1699),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1803),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1722),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1816),
.A2(n_741),
.B1(n_743),
.B2(n_740),
.Y(n_2063)
);

OAI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1816),
.A2(n_748),
.B1(n_749),
.B2(n_744),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1898),
.A2(n_1705),
.B1(n_1823),
.B2(n_1807),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1898),
.A2(n_1202),
.B1(n_1310),
.B2(n_1123),
.Y(n_2066)
);

AO22x2_ASAP7_75t_L g2067 ( 
.A1(n_1961),
.A2(n_948),
.B1(n_1128),
.B2(n_1127),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1705),
.A2(n_1202),
.B1(n_1310),
.B2(n_1123),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1722),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_1983),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1705),
.A2(n_1310),
.B1(n_1202),
.B2(n_1638),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1705),
.A2(n_1310),
.B1(n_1202),
.B2(n_1638),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1704),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1705),
.A2(n_1310),
.B1(n_1202),
.B2(n_1130),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1983),
.B(n_1129),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1729),
.B(n_1202),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1730),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1730),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1882),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1968),
.A2(n_1310),
.B1(n_1202),
.B2(n_1133),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_SL g2081 ( 
.A1(n_1846),
.A2(n_1614),
.B1(n_1617),
.B2(n_1609),
.Y(n_2081)
);

OA22x2_ASAP7_75t_L g2082 ( 
.A1(n_1925),
.A2(n_977),
.B1(n_996),
.B2(n_754),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1736),
.Y(n_2083)
);

OAI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_1816),
.A2(n_1911),
.B1(n_1953),
.B2(n_1952),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1847),
.B(n_1259),
.Y(n_2085)
);

AO22x2_ASAP7_75t_L g2086 ( 
.A1(n_1910),
.A2(n_1135),
.B1(n_1136),
.B2(n_1131),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1954),
.A2(n_748),
.B1(n_749),
.B2(n_744),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_1968),
.A2(n_1139),
.B1(n_1140),
.B2(n_1137),
.Y(n_2088)
);

OAI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_1956),
.A2(n_754),
.B1(n_755),
.B2(n_752),
.Y(n_2089)
);

OAI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_1984),
.A2(n_755),
.B1(n_862),
.B2(n_752),
.Y(n_2090)
);

OR2x6_ASAP7_75t_L g2091 ( 
.A(n_1938),
.B(n_1141),
.Y(n_2091)
);

OA22x2_ASAP7_75t_L g2092 ( 
.A1(n_1975),
.A2(n_990),
.B1(n_1010),
.B2(n_968),
.Y(n_2092)
);

OAI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_1985),
.A2(n_961),
.B1(n_963),
.B2(n_862),
.Y(n_2093)
);

OR2x6_ASAP7_75t_L g2094 ( 
.A(n_1938),
.B(n_1150),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1736),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1704),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1745),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_1968),
.A2(n_1981),
.B1(n_1969),
.B2(n_1756),
.Y(n_2098)
);

AO22x2_ASAP7_75t_L g2099 ( 
.A1(n_1917),
.A2(n_1159),
.B1(n_1161),
.B2(n_1155),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_1851),
.B(n_1162),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1969),
.A2(n_1290),
.B1(n_1330),
.B2(n_1259),
.Y(n_2101)
);

AO22x2_ASAP7_75t_L g2102 ( 
.A1(n_1928),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1745),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1969),
.A2(n_1981),
.B1(n_1741),
.B2(n_1839),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_1981),
.A2(n_1290),
.B1(n_1330),
.B2(n_1259),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1751),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1879),
.B(n_1259),
.Y(n_2107)
);

OR2x6_ASAP7_75t_L g2108 ( 
.A(n_1938),
.B(n_1290),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1879),
.B(n_1290),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1751),
.Y(n_2110)
);

NAND3x1_ASAP7_75t_L g2111 ( 
.A(n_1920),
.B(n_1632),
.C(n_1629),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1762),
.Y(n_2112)
);

OR2x6_ASAP7_75t_L g2113 ( 
.A(n_1938),
.B(n_1330),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_SL g2114 ( 
.A1(n_1918),
.A2(n_1632),
.B1(n_1629),
.B2(n_1402),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1900),
.B(n_1400),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1762),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1958),
.A2(n_1354),
.B1(n_1364),
.B2(n_1330),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1882),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_1958),
.A2(n_1364),
.B1(n_1368),
.B2(n_1354),
.Y(n_2119)
);

AO22x2_ASAP7_75t_L g2120 ( 
.A1(n_1916),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2120)
);

OAI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1739),
.A2(n_963),
.B1(n_966),
.B2(n_961),
.Y(n_2121)
);

OAI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_1743),
.A2(n_968),
.B1(n_971),
.B2(n_966),
.Y(n_2122)
);

NAND2xp33_ASAP7_75t_SL g2123 ( 
.A(n_1943),
.B(n_971),
.Y(n_2123)
);

OAI22xp33_ASAP7_75t_SL g2124 ( 
.A1(n_1841),
.A2(n_978),
.B1(n_979),
.B2(n_977),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1763),
.Y(n_2125)
);

OAI22xp33_ASAP7_75t_SL g2126 ( 
.A1(n_1841),
.A2(n_979),
.B1(n_981),
.B2(n_978),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1915),
.B(n_1354),
.Y(n_2127)
);

AOI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_1958),
.A2(n_1364),
.B1(n_1368),
.B2(n_1354),
.Y(n_2128)
);

OAI22xp5_ASAP7_75t_SL g2129 ( 
.A1(n_1987),
.A2(n_1402),
.B1(n_1404),
.B2(n_1400),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1931),
.A2(n_986),
.B1(n_988),
.B2(n_981),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1763),
.Y(n_2131)
);

OR2x6_ASAP7_75t_L g2132 ( 
.A(n_1885),
.B(n_1364),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1915),
.B(n_1368),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1704),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1974),
.B(n_1368),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1770),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1746),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1902),
.A2(n_988),
.B1(n_990),
.B2(n_986),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1746),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1770),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1773),
.Y(n_2141)
);

AO22x2_ASAP7_75t_L g2142 ( 
.A1(n_1916),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2142)
);

OAI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1902),
.A2(n_996),
.B1(n_997),
.B2(n_993),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1974),
.A2(n_997),
.B1(n_999),
.B2(n_993),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1974),
.B(n_1855),
.Y(n_2145)
);

AO22x2_ASAP7_75t_L g2146 ( 
.A1(n_1946),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2146)
);

AO22x2_ASAP7_75t_L g2147 ( 
.A1(n_1957),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1923),
.A2(n_1001),
.B1(n_1002),
.B2(n_999),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1923),
.A2(n_1002),
.B1(n_1003),
.B2(n_1001),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1773),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1855),
.B(n_1003),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1923),
.A2(n_1012),
.B1(n_1013),
.B2(n_1010),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1904),
.B(n_1012),
.Y(n_2153)
);

INVx8_ASAP7_75t_L g2154 ( 
.A(n_1748),
.Y(n_2154)
);

OAI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1842),
.A2(n_1015),
.B1(n_1017),
.B2(n_1013),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1811),
.B(n_1404),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1778),
.Y(n_2157)
);

OR2x6_ASAP7_75t_L g2158 ( 
.A(n_1885),
.B(n_1407),
.Y(n_2158)
);

AO22x2_ASAP7_75t_L g2159 ( 
.A1(n_1957),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1706),
.A2(n_1017),
.B1(n_1025),
.B2(n_1015),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1706),
.A2(n_1027),
.B1(n_1025),
.B2(n_1407),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1904),
.B(n_1851),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_1789),
.B(n_1027),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1820),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1778),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1948),
.B(n_1432),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1820),
.Y(n_2167)
);

OAI22xp33_ASAP7_75t_L g2168 ( 
.A1(n_1842),
.A2(n_1411),
.B1(n_1431),
.B2(n_1410),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_1728),
.B(n_1909),
.Y(n_2169)
);

AO22x2_ASAP7_75t_L g2170 ( 
.A1(n_1959),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1781),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1781),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1948),
.B(n_1432),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1759),
.B(n_9),
.Y(n_2174)
);

AO22x2_ASAP7_75t_L g2175 ( 
.A1(n_1959),
.A2(n_1963),
.B1(n_1972),
.B2(n_1962),
.Y(n_2175)
);

OAI22xp33_ASAP7_75t_R g2176 ( 
.A1(n_1964),
.A2(n_1411),
.B1(n_1431),
.B2(n_1410),
.Y(n_2176)
);

BUFx2_ASAP7_75t_L g2177 ( 
.A(n_1728),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1849),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1706),
.A2(n_1457),
.B1(n_1479),
.B2(n_1442),
.Y(n_2179)
);

BUFx10_ASAP7_75t_L g2180 ( 
.A(n_1932),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1820),
.Y(n_2181)
);

NAND2xp33_ASAP7_75t_SL g2182 ( 
.A(n_1943),
.B(n_1955),
.Y(n_2182)
);

OR2x6_ASAP7_75t_L g2183 ( 
.A(n_1885),
.B(n_1442),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_1934),
.A2(n_1479),
.B1(n_1486),
.B2(n_1457),
.Y(n_2184)
);

AO22x2_ASAP7_75t_L g2185 ( 
.A1(n_1963),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_1727),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_SL g2187 ( 
.A1(n_1929),
.A2(n_1516),
.B1(n_1520),
.B2(n_1486),
.Y(n_2187)
);

OA22x2_ASAP7_75t_L g2188 ( 
.A1(n_1836),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_1913),
.B(n_12),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1755),
.B(n_1587),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_1755),
.B(n_1587),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_1740),
.A2(n_1520),
.B1(n_1532),
.B2(n_1516),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_1906),
.B(n_13),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1790),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1790),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1905),
.B(n_1532),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1766),
.B(n_1563),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1905),
.B(n_1563),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1796),
.Y(n_2199)
);

OAI22xp33_ASAP7_75t_SL g2200 ( 
.A1(n_1858),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_2200)
);

OAI22xp33_ASAP7_75t_L g2201 ( 
.A1(n_1858),
.A2(n_1576),
.B1(n_1585),
.B2(n_1564),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1929),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1766),
.B(n_1564),
.Y(n_2203)
);

AND2x2_ASAP7_75t_SL g2204 ( 
.A(n_1943),
.B(n_1576),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1951),
.B(n_1585),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1951),
.B(n_1596),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1796),
.Y(n_2207)
);

AO22x2_ASAP7_75t_L g2208 ( 
.A1(n_1979),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1844),
.B(n_1596),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1814),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1814),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_1951),
.B(n_1598),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1815),
.Y(n_2213)
);

OAI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_1859),
.A2(n_1598),
.B1(n_18),
.B2(n_16),
.Y(n_2214)
);

OAI22xp33_ASAP7_75t_SL g2215 ( 
.A1(n_1859),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_1906),
.B(n_1944),
.Y(n_2216)
);

OAI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_1867),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_1740),
.A2(n_125),
.B1(n_126),
.B2(n_124),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_1740),
.A2(n_1866),
.B1(n_1880),
.B2(n_1837),
.Y(n_2219)
);

OAI22xp5_ASAP7_75t_SL g2220 ( 
.A1(n_1942),
.A2(n_28),
.B1(n_36),
.B2(n_19),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_1926),
.B(n_21),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1815),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1826),
.Y(n_2223)
);

AOI22x1_ASAP7_75t_SL g2224 ( 
.A1(n_1942),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1889),
.A2(n_126),
.B1(n_127),
.B2(n_125),
.Y(n_2225)
);

AND2x2_ASAP7_75t_SL g2226 ( 
.A(n_1943),
.B(n_22),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1967),
.B(n_680),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1727),
.Y(n_2228)
);

BUFx10_ASAP7_75t_L g2229 ( 
.A(n_1976),
.Y(n_2229)
);

OAI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_1867),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_2230)
);

INVxp67_ASAP7_75t_L g2231 ( 
.A(n_1905),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1847),
.B(n_1853),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_SL g2233 ( 
.A1(n_1965),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1847),
.B(n_24),
.Y(n_2234)
);

OAI22xp33_ASAP7_75t_L g2235 ( 
.A1(n_1896),
.A2(n_1854),
.B1(n_1868),
.B2(n_1853),
.Y(n_2235)
);

OA22x2_ASAP7_75t_L g2236 ( 
.A1(n_1944),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2236)
);

OR2x6_ASAP7_75t_L g2237 ( 
.A(n_1885),
.B(n_26),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_1732),
.B(n_26),
.Y(n_2238)
);

OR2x6_ASAP7_75t_L g2239 ( 
.A(n_1887),
.B(n_27),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1853),
.B(n_27),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1971),
.B(n_1977),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1937),
.A2(n_128),
.B1(n_130),
.B2(n_127),
.Y(n_2242)
);

OAI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_1896),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2243)
);

OAI22xp33_ASAP7_75t_L g2244 ( 
.A1(n_1854),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1826),
.Y(n_2245)
);

AND2x2_ASAP7_75t_SL g2246 ( 
.A(n_1943),
.B(n_29),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1895),
.Y(n_2247)
);

OAI22xp33_ASAP7_75t_SL g2248 ( 
.A1(n_1737),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2248)
);

OA22x2_ASAP7_75t_L g2249 ( 
.A1(n_1922),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1830),
.Y(n_2250)
);

OAI22xp33_ASAP7_75t_SL g2251 ( 
.A1(n_1742),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2251)
);

OAI22xp33_ASAP7_75t_R g2252 ( 
.A1(n_1798),
.A2(n_43),
.B1(n_51),
.B2(n_34),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_1854),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1830),
.Y(n_2254)
);

OAI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_1868),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_2255)
);

OA22x2_ASAP7_75t_L g2256 ( 
.A1(n_1971),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2256)
);

OAI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_1868),
.A2(n_1877),
.B1(n_1884),
.B2(n_1872),
.Y(n_2257)
);

AOI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_1906),
.A2(n_132),
.B1(n_133),
.B2(n_131),
.Y(n_2258)
);

INVx8_ASAP7_75t_L g2259 ( 
.A(n_1748),
.Y(n_2259)
);

OAI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_1872),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_1801),
.A2(n_134),
.B1(n_135),
.B2(n_132),
.Y(n_2261)
);

AND2x2_ASAP7_75t_SL g2262 ( 
.A(n_1986),
.B(n_1955),
.Y(n_2262)
);

OAI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_1872),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1833),
.Y(n_2264)
);

AOI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_1805),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_1977),
.B(n_692),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1833),
.Y(n_2267)
);

NAND2x1p5_ASAP7_75t_L g2268 ( 
.A(n_1753),
.B(n_40),
.Y(n_2268)
);

OAI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_1877),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2269)
);

AO22x2_ASAP7_75t_L g2270 ( 
.A1(n_1982),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_2270)
);

INVx8_ASAP7_75t_L g2271 ( 
.A(n_1812),
.Y(n_2271)
);

OAI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_1877),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_2272)
);

AO22x2_ASAP7_75t_L g2273 ( 
.A1(n_1982),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1765),
.B(n_46),
.Y(n_2274)
);

AO22x2_ASAP7_75t_L g2275 ( 
.A1(n_1919),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1834),
.Y(n_2276)
);

OAI22xp33_ASAP7_75t_SL g2277 ( 
.A1(n_1806),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1710),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1834),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1927),
.B(n_682),
.Y(n_2280)
);

OR2x6_ASAP7_75t_L g2281 ( 
.A(n_1887),
.B(n_48),
.Y(n_2281)
);

OAI22xp33_ASAP7_75t_SL g2282 ( 
.A1(n_1870),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2282)
);

OAI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_1884),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_1765),
.B(n_52),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1710),
.Y(n_2285)
);

AO22x2_ASAP7_75t_L g2286 ( 
.A1(n_1919),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2286)
);

OR2x6_ASAP7_75t_L g2287 ( 
.A(n_1887),
.B(n_53),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1724),
.Y(n_2288)
);

OAI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_1884),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1724),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_1871),
.A2(n_137),
.B1(n_138),
.B2(n_136),
.Y(n_2291)
);

INVx3_ASAP7_75t_SL g2292 ( 
.A(n_1914),
.Y(n_2292)
);

OAI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_1848),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1927),
.B(n_138),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1749),
.Y(n_2295)
);

AOI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_1894),
.A2(n_140),
.B1(n_141),
.B2(n_139),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_SL g2297 ( 
.A1(n_1702),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_2297)
);

AOI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_1713),
.A2(n_140),
.B1(n_141),
.B2(n_139),
.Y(n_2298)
);

AO22x2_ASAP7_75t_L g2299 ( 
.A1(n_1933),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2299)
);

AO22x2_ASAP7_75t_L g2300 ( 
.A1(n_1933),
.A2(n_1936),
.B1(n_1940),
.B2(n_1939),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1749),
.Y(n_2301)
);

AO22x2_ASAP7_75t_L g2302 ( 
.A1(n_1936),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_1725),
.A2(n_143),
.B1(n_144),
.B2(n_142),
.Y(n_2303)
);

AO22x2_ASAP7_75t_L g2304 ( 
.A1(n_1939),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2304)
);

OAI22xp33_ASAP7_75t_SL g2305 ( 
.A1(n_1702),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1927),
.B(n_688),
.Y(n_2306)
);

OAI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_1848),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_1980),
.Y(n_2308)
);

OR2x6_ASAP7_75t_L g2309 ( 
.A(n_1887),
.B(n_1955),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_1849),
.A2(n_1875),
.B1(n_1881),
.B2(n_1921),
.Y(n_2310)
);

AND2x2_ASAP7_75t_SL g2311 ( 
.A(n_2226),
.B(n_1955),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2031),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2034),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_L g2314 ( 
.A1(n_2221),
.A2(n_1845),
.B1(n_1850),
.B2(n_1843),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2065),
.B(n_1955),
.Y(n_2315)
);

INVx3_ASAP7_75t_L g2316 ( 
.A(n_2004),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_2054),
.B(n_2070),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1998),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2053),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_2262),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1998),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2008),
.Y(n_2322)
);

INVx11_ASAP7_75t_L g2323 ( 
.A(n_2154),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2127),
.B(n_1754),
.Y(n_2324)
);

INVxp33_ASAP7_75t_L g2325 ( 
.A(n_1995),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2075),
.B(n_1966),
.Y(n_2326)
);

AOI22xp33_ASAP7_75t_L g2327 ( 
.A1(n_2238),
.A2(n_1845),
.B1(n_1850),
.B2(n_1843),
.Y(n_2327)
);

NOR2x1p5_ASAP7_75t_L g2328 ( 
.A(n_2009),
.B(n_1721),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2058),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2008),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2011),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_2012),
.B(n_1993),
.Y(n_2332)
);

INVx1_ASAP7_75t_SL g2333 ( 
.A(n_2162),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2104),
.B(n_1966),
.Y(n_2334)
);

NOR3xp33_ASAP7_75t_L g2335 ( 
.A(n_2184),
.B(n_1924),
.C(n_1838),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2098),
.B(n_1966),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2011),
.Y(n_2337)
);

XNOR2xp5_ASAP7_75t_L g2338 ( 
.A(n_2114),
.B(n_1788),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2024),
.Y(n_2339)
);

AND2x6_ASAP7_75t_L g2340 ( 
.A(n_2164),
.B(n_1966),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2024),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2042),
.Y(n_2342)
);

INVx3_ASAP7_75t_L g2343 ( 
.A(n_2004),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2059),
.A2(n_1940),
.B1(n_1731),
.B2(n_1966),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_R g2345 ( 
.A(n_2177),
.B(n_1965),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2042),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2046),
.Y(n_2347)
);

NAND2xp33_ASAP7_75t_SL g2348 ( 
.A(n_2227),
.B(n_1986),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2046),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2047),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2061),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2073),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2073),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_1992),
.B(n_1973),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_2035),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2309),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2047),
.Y(n_2357)
);

BUFx3_ASAP7_75t_L g2358 ( 
.A(n_2309),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2178),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2038),
.B(n_1973),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2241),
.B(n_1986),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2079),
.Y(n_2362)
);

INVx8_ASAP7_75t_L g2363 ( 
.A(n_2108),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2178),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2096),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2079),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2133),
.B(n_1775),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2055),
.B(n_2186),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2190),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2118),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2096),
.Y(n_2371)
);

INVx2_ASAP7_75t_SL g2372 ( 
.A(n_2191),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2107),
.B(n_1733),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2118),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_2178),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_2029),
.Y(n_2376)
);

BUFx6f_ASAP7_75t_L g2377 ( 
.A(n_2035),
.Y(n_2377)
);

NAND2xp33_ASAP7_75t_SL g2378 ( 
.A(n_2280),
.B(n_1973),
.Y(n_2378)
);

AOI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_2246),
.A2(n_1845),
.B1(n_1850),
.B2(n_1843),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_2027),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_2043),
.B(n_1973),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2137),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2137),
.Y(n_2383)
);

AOI22xp5_ASAP7_75t_L g2384 ( 
.A1(n_2231),
.A2(n_1893),
.B1(n_1717),
.B2(n_1921),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2016),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_2308),
.A2(n_1845),
.B1(n_1850),
.B2(n_1843),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_2197),
.Y(n_2387)
);

CKINVDCx11_ASAP7_75t_R g2388 ( 
.A(n_2292),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2134),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2139),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2134),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2109),
.B(n_1843),
.Y(n_2392)
);

INVx4_ASAP7_75t_L g2393 ( 
.A(n_2186),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_SL g2394 ( 
.A(n_2050),
.B(n_1812),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2139),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2194),
.Y(n_2396)
);

INVx1_ASAP7_75t_SL g2397 ( 
.A(n_2169),
.Y(n_2397)
);

AOI22xp33_ASAP7_75t_L g2398 ( 
.A1(n_2193),
.A2(n_1850),
.B1(n_1864),
.B2(n_1845),
.Y(n_2398)
);

NAND3xp33_ASAP7_75t_L g2399 ( 
.A(n_2115),
.B(n_1978),
.C(n_1973),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_2228),
.Y(n_2400)
);

INVx4_ASAP7_75t_L g2401 ( 
.A(n_2228),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2194),
.Y(n_2402)
);

AOI22xp33_ASAP7_75t_L g2403 ( 
.A1(n_2247),
.A2(n_1874),
.B1(n_1864),
.B2(n_1771),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_2154),
.Y(n_2404)
);

AND2x6_ASAP7_75t_L g2405 ( 
.A(n_2164),
.B(n_1986),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2207),
.Y(n_2406)
);

NAND2xp33_ASAP7_75t_SL g2407 ( 
.A(n_2294),
.B(n_1986),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2207),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_2019),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2222),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2222),
.Y(n_2411)
);

OAI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2216),
.A2(n_1941),
.B1(n_1930),
.B2(n_1881),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2223),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2278),
.B(n_1864),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2108),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_2021),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2278),
.B(n_1950),
.Y(n_2417)
);

BUFx8_ASAP7_75t_SL g2418 ( 
.A(n_2158),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2285),
.B(n_1864),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2223),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2145),
.B(n_1864),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_1996),
.B(n_1980),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2100),
.B(n_1930),
.Y(n_2423)
);

INVx5_ASAP7_75t_L g2424 ( 
.A(n_2113),
.Y(n_2424)
);

INVx3_ASAP7_75t_L g2425 ( 
.A(n_2167),
.Y(n_2425)
);

INVx4_ASAP7_75t_L g2426 ( 
.A(n_2113),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2245),
.Y(n_2427)
);

NOR2x1p5_ASAP7_75t_L g2428 ( 
.A(n_2056),
.B(n_1721),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2017),
.B(n_1941),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2245),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_2259),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2254),
.Y(n_2432)
);

NAND3xp33_ASAP7_75t_SL g2433 ( 
.A(n_2018),
.B(n_2020),
.C(n_2040),
.Y(n_2433)
);

INVx1_ASAP7_75t_SL g2434 ( 
.A(n_2203),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_2259),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2254),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2285),
.Y(n_2437)
);

INVx4_ASAP7_75t_L g2438 ( 
.A(n_2300),
.Y(n_2438)
);

AND2x6_ASAP7_75t_L g2439 ( 
.A(n_2167),
.B(n_1753),
.Y(n_2439)
);

BUFx4f_ASAP7_75t_L g2440 ( 
.A(n_2306),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2288),
.Y(n_2441)
);

INVx6_ASAP7_75t_L g2442 ( 
.A(n_2132),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_2158),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2007),
.B(n_1883),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2181),
.Y(n_2445)
);

BUFx4f_ASAP7_75t_L g2446 ( 
.A(n_2204),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2288),
.Y(n_2447)
);

OR2x6_ASAP7_75t_L g2448 ( 
.A(n_2271),
.B(n_1903),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2181),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2290),
.Y(n_2450)
);

BUFx3_ASAP7_75t_L g2451 ( 
.A(n_2271),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2290),
.Y(n_2452)
);

OR2x6_ASAP7_75t_L g2453 ( 
.A(n_2052),
.B(n_1903),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2183),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2044),
.B(n_1883),
.Y(n_2455)
);

AOI22xp33_ASAP7_75t_L g2456 ( 
.A1(n_2295),
.A2(n_1874),
.B1(n_1771),
.B2(n_1776),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2219),
.A2(n_1875),
.B1(n_1878),
.B2(n_1869),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2295),
.Y(n_2458)
);

AND2x2_ASAP7_75t_SL g2459 ( 
.A(n_2258),
.B(n_1878),
.Y(n_2459)
);

INVx8_ASAP7_75t_L g2460 ( 
.A(n_2052),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2301),
.A2(n_1874),
.B1(n_1774),
.B2(n_1776),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2084),
.B(n_1874),
.Y(n_2462)
);

INVxp33_ASAP7_75t_L g2463 ( 
.A(n_2033),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2301),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2025),
.B(n_1914),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2045),
.B(n_1869),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2264),
.B(n_1874),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_L g2468 ( 
.A1(n_2267),
.A2(n_1774),
.B1(n_1783),
.B2(n_1777),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2062),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2069),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2077),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2276),
.B(n_1777),
.Y(n_2472)
);

AOI22xp33_ASAP7_75t_L g2473 ( 
.A1(n_2279),
.A2(n_1783),
.B1(n_1785),
.B2(n_1784),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2078),
.Y(n_2474)
);

CKINVDCx20_ASAP7_75t_R g2475 ( 
.A(n_2051),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_2300),
.Y(n_2476)
);

BUFx10_ASAP7_75t_L g2477 ( 
.A(n_2202),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2310),
.B(n_1818),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_2083),
.A2(n_1784),
.B1(n_1810),
.B2(n_1785),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2095),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2232),
.B(n_1810),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2071),
.B(n_1818),
.Y(n_2482)
);

OAI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2039),
.A2(n_1873),
.B(n_1878),
.Y(n_2483)
);

BUFx3_ASAP7_75t_L g2484 ( 
.A(n_2183),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2097),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2174),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2006),
.B(n_1950),
.Y(n_2487)
);

CKINVDCx14_ASAP7_75t_R g2488 ( 
.A(n_2081),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2103),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2106),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2110),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2112),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_2072),
.B(n_1818),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2235),
.B(n_1817),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2257),
.B(n_1818),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_1994),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2116),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2125),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2131),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2136),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2140),
.Y(n_2501)
);

AND2x6_ASAP7_75t_L g2502 ( 
.A(n_2066),
.B(n_1852),
.Y(n_2502)
);

AND2x2_ASAP7_75t_SL g2503 ( 
.A(n_2218),
.B(n_1717),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2141),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_1990),
.B(n_1760),
.Y(n_2505)
);

INVxp67_ASAP7_75t_SL g2506 ( 
.A(n_2002),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2088),
.B(n_1817),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2001),
.B(n_1818),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2266),
.B(n_2151),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2174),
.B(n_1852),
.Y(n_2510)
);

INVx1_ASAP7_75t_SL g2511 ( 
.A(n_2166),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2150),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2157),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2165),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2153),
.B(n_1907),
.Y(n_2515)
);

OAI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2091),
.A2(n_2094),
.B1(n_2010),
.B2(n_2041),
.Y(n_2516)
);

INVx4_ASAP7_75t_L g2517 ( 
.A(n_2015),
.Y(n_2517)
);

HB1xp67_ASAP7_75t_L g2518 ( 
.A(n_2274),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2171),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2172),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2195),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2274),
.Y(n_2522)
);

BUFx3_ASAP7_75t_L g2523 ( 
.A(n_2048),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2199),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_2036),
.B(n_1760),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2210),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2211),
.B(n_1819),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2213),
.B(n_1819),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2250),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2085),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2234),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2048),
.Y(n_2532)
);

INVx3_ASAP7_75t_L g2533 ( 
.A(n_2284),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2240),
.Y(n_2534)
);

XNOR2xp5_ASAP7_75t_L g2535 ( 
.A(n_2129),
.B(n_1907),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2284),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2076),
.B(n_1824),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2180),
.B(n_1856),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2080),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2013),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2013),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2091),
.B(n_1908),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2094),
.B(n_1908),
.Y(n_2543)
);

INVx6_ASAP7_75t_L g2544 ( 
.A(n_2132),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2135),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_1991),
.B(n_1831),
.Y(n_2546)
);

BUFx2_ASAP7_75t_L g2547 ( 
.A(n_2173),
.Y(n_2547)
);

INVx5_ASAP7_75t_L g2548 ( 
.A(n_2237),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2086),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2256),
.Y(n_2550)
);

INVx3_ASAP7_75t_L g2551 ( 
.A(n_2175),
.Y(n_2551)
);

AOI22xp33_ASAP7_75t_L g2552 ( 
.A1(n_2188),
.A2(n_1824),
.B1(n_1829),
.B2(n_1828),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2086),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2275),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2163),
.A2(n_1828),
.B1(n_1832),
.B2(n_1829),
.Y(n_2555)
);

INVx6_ASAP7_75t_L g2556 ( 
.A(n_2180),
.Y(n_2556)
);

INVx2_ASAP7_75t_SL g2557 ( 
.A(n_2060),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2099),
.Y(n_2558)
);

BUFx2_ASAP7_75t_L g2559 ( 
.A(n_2237),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2275),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2229),
.B(n_2022),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2286),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2286),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2099),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2101),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2105),
.Y(n_2566)
);

INVxp67_ASAP7_75t_SL g2567 ( 
.A(n_2117),
.Y(n_2567)
);

OAI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_2175),
.A2(n_1832),
.B1(n_1862),
.B2(n_1856),
.Y(n_2568)
);

INVx4_ASAP7_75t_SL g2569 ( 
.A(n_2239),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2119),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2089),
.B(n_1862),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2229),
.B(n_1865),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2090),
.B(n_1865),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2168),
.B(n_1888),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2128),
.Y(n_2575)
);

AND2x6_ASAP7_75t_L g2576 ( 
.A(n_2068),
.B(n_1888),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2236),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2182),
.B(n_1831),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2010),
.B(n_1895),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2299),
.Y(n_2580)
);

INVx2_ASAP7_75t_SL g2581 ( 
.A(n_2189),
.Y(n_2581)
);

AOI22xp33_ASAP7_75t_L g2582 ( 
.A1(n_2121),
.A2(n_1892),
.B1(n_1897),
.B2(n_1876),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2201),
.B(n_1892),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2299),
.Y(n_2584)
);

INVx4_ASAP7_75t_L g2585 ( 
.A(n_2302),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2302),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2304),
.Y(n_2587)
);

INVx5_ASAP7_75t_L g2588 ( 
.A(n_2239),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2304),
.Y(n_2589)
);

INVx2_ASAP7_75t_SL g2590 ( 
.A(n_2281),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2270),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2270),
.Y(n_2592)
);

INVx4_ASAP7_75t_L g2593 ( 
.A(n_2273),
.Y(n_2593)
);

NAND3xp33_ASAP7_75t_L g2594 ( 
.A(n_2156),
.B(n_1897),
.C(n_1715),
.Y(n_2594)
);

OAI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2242),
.A2(n_1723),
.B1(n_1813),
.B2(n_1727),
.Y(n_2595)
);

INVx2_ASAP7_75t_SL g2596 ( 
.A(n_2281),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2273),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2120),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2120),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2142),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2122),
.A2(n_1876),
.B1(n_1831),
.B2(n_1780),
.Y(n_2601)
);

BUFx10_ASAP7_75t_L g2602 ( 
.A(n_2209),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2142),
.Y(n_2603)
);

OAI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2225),
.A2(n_1831),
.B1(n_1804),
.B2(n_1792),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2249),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2074),
.B(n_2049),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2208),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2208),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2268),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2093),
.A2(n_1876),
.B1(n_1831),
.B2(n_1780),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2147),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2147),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2159),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2160),
.B(n_1747),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2272),
.Y(n_2615)
);

INVxp67_ASAP7_75t_L g2616 ( 
.A(n_2032),
.Y(n_2616)
);

INVxp67_ASAP7_75t_SL g2617 ( 
.A(n_2179),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2159),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2082),
.A2(n_1876),
.B1(n_1780),
.B2(n_1786),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2287),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2187),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2192),
.B(n_1747),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2170),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_2205),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2092),
.A2(n_1876),
.B1(n_1786),
.B2(n_1779),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2170),
.Y(n_2626)
);

INVx2_ASAP7_75t_SL g2627 ( 
.A(n_2287),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2298),
.Y(n_2628)
);

BUFx2_ASAP7_75t_L g2629 ( 
.A(n_2206),
.Y(n_2629)
);

INVx3_ASAP7_75t_L g2630 ( 
.A(n_2185),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2220),
.B(n_1738),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2028),
.B(n_1738),
.Y(n_2632)
);

INVx4_ASAP7_75t_L g2633 ( 
.A(n_2185),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2130),
.B(n_1747),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2196),
.B(n_1935),
.Y(n_2635)
);

INVxp67_ASAP7_75t_L g2636 ( 
.A(n_2198),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2102),
.Y(n_2637)
);

AND2x6_ASAP7_75t_L g2638 ( 
.A(n_2303),
.B(n_1738),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2000),
.B(n_1809),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2014),
.B(n_1738),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2000),
.B(n_1809),
.Y(n_2641)
);

INVx1_ASAP7_75t_SL g2642 ( 
.A(n_2212),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2102),
.Y(n_2643)
);

BUFx3_ASAP7_75t_L g2644 ( 
.A(n_2005),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2146),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2003),
.B(n_1809),
.Y(n_2646)
);

OAI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2087),
.A2(n_1873),
.B(n_1786),
.Y(n_2647)
);

AND2x6_ASAP7_75t_L g2648 ( 
.A(n_2261),
.B(n_1738),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2037),
.B(n_1804),
.Y(n_2649)
);

CKINVDCx20_ASAP7_75t_R g2650 ( 
.A(n_2023),
.Y(n_2650)
);

AOI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2123),
.A2(n_1876),
.B1(n_1723),
.B2(n_1804),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2146),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2067),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2063),
.B(n_1723),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2067),
.A2(n_1779),
.B1(n_1752),
.B2(n_1757),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2057),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2057),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_SL g2658 ( 
.A(n_2064),
.B(n_1750),
.Y(n_2658)
);

BUFx10_ASAP7_75t_L g2659 ( 
.A(n_2111),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2244),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2253),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2255),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2161),
.A2(n_1835),
.B1(n_1891),
.B2(n_1822),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2265),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2260),
.Y(n_2665)
);

AO22x2_ASAP7_75t_L g2666 ( 
.A1(n_2633),
.A2(n_2224),
.B1(n_2176),
.B2(n_2252),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2332),
.B(n_2509),
.Y(n_2667)
);

BUFx3_ASAP7_75t_L g2668 ( 
.A(n_2404),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2360),
.B(n_2144),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2359),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2464),
.Y(n_2671)
);

INVxp67_ASAP7_75t_L g2672 ( 
.A(n_2509),
.Y(n_2672)
);

OAI22xp5_ASAP7_75t_SL g2673 ( 
.A1(n_2650),
.A2(n_2252),
.B1(n_2176),
.B2(n_2148),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2311),
.A2(n_2296),
.B1(n_2291),
.B2(n_2269),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2464),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2534),
.B(n_1779),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2377),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2406),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2406),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2427),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2427),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_2359),
.Y(n_2682)
);

INVx4_ASAP7_75t_L g2683 ( 
.A(n_2359),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2531),
.B(n_1744),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2437),
.Y(n_2685)
);

INVx3_ASAP7_75t_L g2686 ( 
.A(n_2377),
.Y(n_2686)
);

AND2x6_ASAP7_75t_L g2687 ( 
.A(n_2320),
.B(n_2149),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2333),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2471),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2441),
.Y(n_2690)
);

BUFx4f_ASAP7_75t_L g2691 ( 
.A(n_2448),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2447),
.Y(n_2692)
);

INVxp67_ASAP7_75t_L g2693 ( 
.A(n_2547),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2311),
.A2(n_2283),
.B1(n_2289),
.B2(n_2263),
.Y(n_2694)
);

NAND3xp33_ASAP7_75t_L g2695 ( 
.A(n_2381),
.B(n_2583),
.C(n_2574),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2450),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2380),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2471),
.Y(n_2698)
);

BUFx2_ASAP7_75t_L g2699 ( 
.A(n_2376),
.Y(n_2699)
);

INVx3_ASAP7_75t_L g2700 ( 
.A(n_2377),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2490),
.Y(n_2701)
);

INVx4_ASAP7_75t_L g2702 ( 
.A(n_2359),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2511),
.B(n_2152),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2388),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2397),
.B(n_2138),
.Y(n_2705)
);

AO22x2_ASAP7_75t_L g2706 ( 
.A1(n_2633),
.A2(n_2224),
.B1(n_2233),
.B2(n_2214),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2354),
.B(n_1822),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2531),
.B(n_2373),
.Y(n_2708)
);

AOI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_2503),
.A2(n_2433),
.B1(n_2628),
.B2(n_2515),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2490),
.Y(n_2710)
);

AND2x6_ASAP7_75t_L g2711 ( 
.A(n_2320),
.B(n_1750),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2326),
.B(n_2354),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2492),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2492),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2452),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2364),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2324),
.B(n_1744),
.Y(n_2717)
);

AND2x6_ASAP7_75t_L g2718 ( 
.A(n_2320),
.B(n_2445),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2458),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2396),
.Y(n_2720)
);

INVx4_ASAP7_75t_L g2721 ( 
.A(n_2364),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2518),
.Y(n_2722)
);

OAI22x1_ASAP7_75t_R g2723 ( 
.A1(n_2475),
.A2(n_1935),
.B1(n_1715),
.B2(n_2026),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_2364),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2326),
.B(n_2003),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2364),
.Y(n_2726)
);

AO22x2_ASAP7_75t_L g2727 ( 
.A1(n_2633),
.A2(n_1999),
.B1(n_1997),
.B2(n_2030),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2498),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_L g2729 ( 
.A(n_2616),
.B(n_2143),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2402),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2408),
.Y(n_2731)
);

AND2x6_ASAP7_75t_L g2732 ( 
.A(n_2320),
.B(n_1750),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2410),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_2375),
.Y(n_2734)
);

INVx4_ASAP7_75t_SL g2735 ( 
.A(n_2340),
.Y(n_2735)
);

HB1xp67_ASAP7_75t_L g2736 ( 
.A(n_2369),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2325),
.B(n_2155),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2411),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2375),
.Y(n_2739)
);

BUFx6f_ASAP7_75t_L g2740 ( 
.A(n_2375),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2413),
.Y(n_2741)
);

AO22x2_ASAP7_75t_L g2742 ( 
.A1(n_2585),
.A2(n_2593),
.B1(n_2608),
.B2(n_2607),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2498),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2504),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2504),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2519),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2420),
.Y(n_2747)
);

AOI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2503),
.A2(n_2307),
.B1(n_2293),
.B2(n_2230),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_L g2749 ( 
.A(n_2325),
.B(n_2124),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_L g2750 ( 
.A1(n_2607),
.A2(n_2243),
.B1(n_2217),
.B2(n_2215),
.Y(n_2750)
);

INVxp67_ASAP7_75t_SL g2751 ( 
.A(n_2318),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2519),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2486),
.B(n_1822),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2430),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2432),
.Y(n_2755)
);

OR2x6_ASAP7_75t_L g2756 ( 
.A(n_2460),
.B(n_2448),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2367),
.B(n_1744),
.Y(n_2757)
);

AND2x2_ASAP7_75t_SL g2758 ( 
.A(n_2446),
.B(n_1715),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2486),
.B(n_1835),
.Y(n_2759)
);

BUFx6f_ASAP7_75t_L g2760 ( 
.A(n_2375),
.Y(n_2760)
);

NAND3x1_ASAP7_75t_L g2761 ( 
.A(n_2505),
.B(n_1935),
.C(n_2126),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2385),
.B(n_2434),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2520),
.Y(n_2763)
);

AND2x6_ASAP7_75t_L g2764 ( 
.A(n_2445),
.B(n_1750),
.Y(n_2764)
);

BUFx3_ASAP7_75t_L g2765 ( 
.A(n_2404),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2423),
.B(n_2557),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2481),
.B(n_1752),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2557),
.B(n_1997),
.Y(n_2768)
);

BUFx3_ASAP7_75t_L g2769 ( 
.A(n_2431),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_SL g2770 ( 
.A1(n_2650),
.A2(n_1999),
.B1(n_2251),
.B2(n_2248),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2388),
.Y(n_2771)
);

BUFx2_ASAP7_75t_L g2772 ( 
.A(n_2629),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2436),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2520),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2526),
.Y(n_2775)
);

AND2x4_ASAP7_75t_L g2776 ( 
.A(n_2486),
.B(n_1835),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2312),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2313),
.Y(n_2778)
);

BUFx6f_ASAP7_75t_L g2779 ( 
.A(n_2415),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2319),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2329),
.Y(n_2781)
);

INVx2_ASAP7_75t_SL g2782 ( 
.A(n_2423),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2415),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2351),
.Y(n_2784)
);

BUFx4f_ASAP7_75t_L g2785 ( 
.A(n_2448),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2463),
.B(n_2277),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_2415),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2463),
.B(n_2282),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2449),
.Y(n_2789)
);

AOI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2515),
.A2(n_2030),
.B1(n_1891),
.B2(n_2200),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2526),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2369),
.B(n_2372),
.Y(n_2792)
);

INVx2_ASAP7_75t_SL g2793 ( 
.A(n_2579),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2372),
.B(n_1891),
.Y(n_2794)
);

NAND2xp33_ASAP7_75t_L g2795 ( 
.A(n_2340),
.B(n_1750),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2449),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2318),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2422),
.A2(n_2305),
.B1(n_2297),
.B2(n_1799),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2409),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2321),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2321),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2322),
.Y(n_2802)
);

NAND2x1p5_ASAP7_75t_L g2803 ( 
.A(n_2393),
.B(n_2400),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2409),
.Y(n_2804)
);

INVx4_ASAP7_75t_L g2805 ( 
.A(n_2424),
.Y(n_2805)
);

BUFx2_ASAP7_75t_L g2806 ( 
.A(n_2629),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2322),
.Y(n_2807)
);

AND2x4_ASAP7_75t_L g2808 ( 
.A(n_2486),
.B(n_1701),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2636),
.B(n_1761),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2330),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2446),
.B(n_1761),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_2642),
.B(n_1761),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2330),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2331),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2331),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2387),
.B(n_1752),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2337),
.Y(n_2817)
);

HB1xp67_ASAP7_75t_L g2818 ( 
.A(n_2387),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2337),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2415),
.Y(n_2820)
);

INVx3_ASAP7_75t_L g2821 ( 
.A(n_2377),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2409),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2339),
.Y(n_2823)
);

AO22x2_ASAP7_75t_L g2824 ( 
.A1(n_2585),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2422),
.A2(n_1757),
.B1(n_1764),
.B2(n_1761),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2339),
.B(n_2341),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2341),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2342),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2342),
.B(n_2346),
.Y(n_2829)
);

OR2x2_ASAP7_75t_L g2830 ( 
.A(n_2617),
.B(n_1794),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2346),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2347),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2347),
.B(n_1757),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2349),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2349),
.B(n_1735),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2522),
.B(n_1701),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2416),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2455),
.B(n_1735),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2416),
.Y(n_2839)
);

AOI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2664),
.A2(n_1791),
.B1(n_1793),
.B2(n_1735),
.Y(n_2840)
);

INVx5_ASAP7_75t_L g2841 ( 
.A(n_2340),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2466),
.B(n_1791),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2350),
.B(n_1791),
.Y(n_2843)
);

INVx8_ASAP7_75t_L g2844 ( 
.A(n_2363),
.Y(n_2844)
);

HB1xp67_ASAP7_75t_L g2845 ( 
.A(n_2438),
.Y(n_2845)
);

OR2x6_ASAP7_75t_L g2846 ( 
.A(n_2460),
.B(n_1761),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_SL g2847 ( 
.A(n_2446),
.B(n_1764),
.Y(n_2847)
);

BUFx6f_ASAP7_75t_L g2848 ( 
.A(n_2442),
.Y(n_2848)
);

BUFx2_ASAP7_75t_L g2849 ( 
.A(n_2559),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2416),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2412),
.B(n_1764),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2355),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2522),
.B(n_1701),
.Y(n_2853)
);

BUFx10_ASAP7_75t_L g2854 ( 
.A(n_2444),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2382),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2350),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2357),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2622),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2357),
.Y(n_2859)
);

HB1xp67_ASAP7_75t_L g2860 ( 
.A(n_2438),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2362),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2362),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2382),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2366),
.B(n_2370),
.Y(n_2864)
);

INVx3_ASAP7_75t_L g2865 ( 
.A(n_2355),
.Y(n_2865)
);

OAI221xp5_ASAP7_75t_L g2866 ( 
.A1(n_2552),
.A2(n_1802),
.B1(n_1793),
.B2(n_1764),
.C(n_1797),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2366),
.B(n_1793),
.Y(n_2867)
);

BUFx10_ASAP7_75t_L g2868 ( 
.A(n_2635),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2370),
.Y(n_2869)
);

INVx4_ASAP7_75t_L g2870 ( 
.A(n_2424),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2429),
.B(n_1764),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2383),
.Y(n_2872)
);

AOI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2487),
.A2(n_1797),
.B1(n_1800),
.B2(n_1795),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2383),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2374),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2374),
.B(n_1802),
.Y(n_2876)
);

AOI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2664),
.A2(n_1802),
.B1(n_1718),
.B2(n_1716),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2472),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2390),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2527),
.Y(n_2880)
);

AO22x2_ASAP7_75t_L g2881 ( 
.A1(n_2585),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_2487),
.A2(n_1797),
.B1(n_1800),
.B2(n_1795),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2537),
.B(n_1795),
.Y(n_2883)
);

OAI22xp33_ASAP7_75t_L g2884 ( 
.A1(n_2593),
.A2(n_1797),
.B1(n_1800),
.B2(n_1795),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2528),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2579),
.B(n_693),
.Y(n_2886)
);

BUFx6f_ASAP7_75t_L g2887 ( 
.A(n_2442),
.Y(n_2887)
);

INVx4_ASAP7_75t_L g2888 ( 
.A(n_2424),
.Y(n_2888)
);

BUFx2_ASAP7_75t_L g2889 ( 
.A(n_2559),
.Y(n_2889)
);

BUFx4f_ASAP7_75t_L g2890 ( 
.A(n_2448),
.Y(n_2890)
);

AO22x2_ASAP7_75t_L g2891 ( 
.A1(n_2593),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2522),
.B(n_1716),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2469),
.Y(n_2893)
);

BUFx3_ASAP7_75t_L g2894 ( 
.A(n_2431),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2442),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2435),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2602),
.B(n_142),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2470),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2602),
.B(n_1795),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_2522),
.B(n_1716),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2474),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2494),
.B(n_1797),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2480),
.Y(n_2903)
);

OR2x2_ASAP7_75t_L g2904 ( 
.A(n_2622),
.B(n_1800),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2602),
.B(n_1800),
.Y(n_2905)
);

INVx4_ASAP7_75t_L g2906 ( 
.A(n_2424),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2581),
.B(n_144),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_2355),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2438),
.A2(n_1718),
.B1(n_1716),
.B2(n_1709),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2485),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2489),
.Y(n_2911)
);

AND2x4_ASAP7_75t_L g2912 ( 
.A(n_2523),
.B(n_1716),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2491),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2497),
.Y(n_2914)
);

BUFx4f_ASAP7_75t_L g2915 ( 
.A(n_2460),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2499),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2390),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2500),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2395),
.Y(n_2919)
);

BUFx3_ASAP7_75t_L g2920 ( 
.A(n_2435),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2501),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2425),
.B(n_1718),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2581),
.Y(n_2923)
);

INVx2_ASAP7_75t_SL g2924 ( 
.A(n_2454),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2624),
.B(n_146),
.Y(n_2925)
);

NAND3xp33_ASAP7_75t_L g2926 ( 
.A(n_2399),
.B(n_1718),
.C(n_1709),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2512),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2513),
.Y(n_2928)
);

NAND2xp33_ASAP7_75t_L g2929 ( 
.A(n_2340),
.B(n_1718),
.Y(n_2929)
);

AND2x4_ASAP7_75t_L g2930 ( 
.A(n_2523),
.B(n_1708),
.Y(n_2930)
);

INVxp67_ASAP7_75t_L g2931 ( 
.A(n_2605),
.Y(n_2931)
);

NAND3xp33_ASAP7_75t_SL g2932 ( 
.A(n_2561),
.B(n_67),
.C(n_69),
.Y(n_2932)
);

NAND2x1p5_ASAP7_75t_L g2933 ( 
.A(n_2393),
.B(n_1708),
.Y(n_2933)
);

OA22x2_ASAP7_75t_L g2934 ( 
.A1(n_2645),
.A2(n_2652),
.B1(n_2630),
.B2(n_2611),
.Y(n_2934)
);

BUFx2_ASAP7_75t_L g2935 ( 
.A(n_2624),
.Y(n_2935)
);

AND2x4_ASAP7_75t_L g2936 ( 
.A(n_2536),
.B(n_2533),
.Y(n_2936)
);

AOI22x1_ASAP7_75t_L g2937 ( 
.A1(n_2539),
.A2(n_1709),
.B1(n_1712),
.B2(n_1708),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2514),
.Y(n_2938)
);

INVxp67_ASAP7_75t_L g2939 ( 
.A(n_2361),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2521),
.Y(n_2940)
);

AO22x2_ASAP7_75t_L g2941 ( 
.A1(n_2608),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2533),
.B(n_1708),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2316),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_L g2944 ( 
.A(n_2442),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2614),
.B(n_679),
.Y(n_2945)
);

AND2x4_ASAP7_75t_L g2946 ( 
.A(n_2533),
.B(n_2317),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2538),
.B(n_1708),
.Y(n_2947)
);

INVxp67_ASAP7_75t_L g2948 ( 
.A(n_2361),
.Y(n_2948)
);

OAI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2554),
.A2(n_1712),
.B1(n_1709),
.B2(n_71),
.Y(n_2949)
);

AOI22xp5_ASAP7_75t_L g2950 ( 
.A1(n_2551),
.A2(n_1712),
.B1(n_1709),
.B2(n_147),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2614),
.B(n_679),
.Y(n_2951)
);

BUFx6f_ASAP7_75t_L g2952 ( 
.A(n_2544),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2524),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2316),
.Y(n_2954)
);

CKINVDCx16_ASAP7_75t_R g2955 ( 
.A(n_2345),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2572),
.B(n_1712),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2317),
.B(n_680),
.Y(n_2957)
);

NAND2x1p5_ASAP7_75t_L g2958 ( 
.A(n_2393),
.B(n_1712),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2934),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2955),
.B(n_2548),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2667),
.B(n_2550),
.Y(n_2961)
);

A2O1A1Ixp33_ASAP7_75t_L g2962 ( 
.A1(n_2669),
.A2(n_2440),
.B(n_2348),
.C(n_2407),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2708),
.B(n_2550),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2858),
.B(n_2645),
.Y(n_2964)
);

AND2x6_ASAP7_75t_L g2965 ( 
.A(n_2950),
.B(n_2554),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2858),
.B(n_2652),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2672),
.B(n_2465),
.Y(n_2967)
);

A2O1A1Ixp33_ASAP7_75t_L g2968 ( 
.A1(n_2695),
.A2(n_2440),
.B(n_2348),
.C(n_2407),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2934),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2708),
.B(n_2550),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2678),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2680),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2712),
.B(n_2577),
.Y(n_2973)
);

INVx2_ASAP7_75t_SL g2974 ( 
.A(n_2697),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2685),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2668),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2681),
.Y(n_2977)
);

NAND2x1p5_ASAP7_75t_L g2978 ( 
.A(n_2805),
.B(n_2424),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2703),
.B(n_2639),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_L g2980 ( 
.A(n_2672),
.B(n_2465),
.Y(n_2980)
);

AOI22xp33_ASAP7_75t_L g2981 ( 
.A1(n_2932),
.A2(n_2615),
.B1(n_2661),
.B2(n_2660),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_2782),
.B(n_2548),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2690),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2692),
.Y(n_2984)
);

INVx2_ASAP7_75t_SL g2985 ( 
.A(n_2765),
.Y(n_2985)
);

NAND2xp33_ASAP7_75t_L g2986 ( 
.A(n_2695),
.B(n_2340),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2762),
.B(n_2548),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2878),
.B(n_2880),
.Y(n_2988)
);

BUFx6f_ASAP7_75t_L g2989 ( 
.A(n_2670),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2766),
.B(n_2548),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2885),
.B(n_2577),
.Y(n_2991)
);

INVx3_ASAP7_75t_L g2992 ( 
.A(n_2805),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2931),
.B(n_2577),
.Y(n_2993)
);

A2O1A1Ixp33_ASAP7_75t_L g2994 ( 
.A1(n_2709),
.A2(n_2440),
.B(n_2378),
.C(n_2315),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2931),
.B(n_2662),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2673),
.A2(n_2335),
.B1(n_2525),
.B2(n_2516),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2709),
.A2(n_2400),
.B1(n_2401),
.B2(n_2314),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2792),
.B(n_2665),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2671),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2693),
.B(n_2643),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2751),
.A2(n_2401),
.B1(n_2400),
.B2(n_2403),
.Y(n_3001)
);

O2A1O1Ixp5_ASAP7_75t_L g3002 ( 
.A1(n_2851),
.A2(n_2334),
.B(n_2315),
.C(n_2336),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2675),
.Y(n_3003)
);

NAND2x1_ASAP7_75t_L g3004 ( 
.A(n_2718),
.B(n_2401),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2932),
.A2(n_2630),
.B1(n_2535),
.B2(n_2553),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2699),
.B(n_2548),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2696),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_SL g3008 ( 
.A(n_2854),
.B(n_2588),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_SL g3009 ( 
.A1(n_2673),
.A2(n_2475),
.B1(n_2338),
.B2(n_2621),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2679),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2751),
.B(n_2317),
.Y(n_3011)
);

CKINVDCx5p33_ASAP7_75t_R g3012 ( 
.A(n_2704),
.Y(n_3012)
);

INVx2_ASAP7_75t_SL g3013 ( 
.A(n_2769),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2830),
.B(n_2600),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2715),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2693),
.B(n_2637),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2674),
.A2(n_2630),
.B1(n_2535),
.B2(n_2558),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2707),
.B(n_2603),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2854),
.B(n_2588),
.Y(n_3019)
);

OAI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2748),
.A2(n_2611),
.B1(n_2613),
.B2(n_2612),
.Y(n_3020)
);

INVxp67_ASAP7_75t_SL g3021 ( 
.A(n_2884),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2707),
.B(n_2555),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2719),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2855),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2863),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_2705),
.B(n_2637),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2688),
.B(n_2588),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2838),
.B(n_2589),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2725),
.B(n_2580),
.Y(n_3029)
);

AND2x4_ASAP7_75t_L g3030 ( 
.A(n_2793),
.B(n_2356),
.Y(n_3030)
);

HB1xp67_ASAP7_75t_L g3031 ( 
.A(n_2688),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2946),
.B(n_2588),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2720),
.Y(n_3033)
);

NAND3xp33_ASAP7_75t_L g3034 ( 
.A(n_2729),
.B(n_2594),
.C(n_2394),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2872),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2945),
.B(n_2592),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2874),
.Y(n_3037)
);

AOI22xp33_ASAP7_75t_L g3038 ( 
.A1(n_2674),
.A2(n_2549),
.B1(n_2564),
.B2(n_2562),
.Y(n_3038)
);

BUFx2_ASAP7_75t_L g3039 ( 
.A(n_2849),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2730),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2731),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2795),
.A2(n_2368),
.B(n_2334),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2737),
.B(n_2637),
.Y(n_3043)
);

NAND2xp33_ASAP7_75t_L g3044 ( 
.A(n_2718),
.B(n_2340),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2951),
.B(n_2587),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2733),
.Y(n_3046)
);

AOI22xp5_ASAP7_75t_L g3047 ( 
.A1(n_2687),
.A2(n_2609),
.B1(n_2344),
.B2(n_2443),
.Y(n_3047)
);

AND2x6_ASAP7_75t_SL g3048 ( 
.A(n_2749),
.B(n_2453),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2772),
.B(n_2643),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2886),
.B(n_2639),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2748),
.B(n_2584),
.Y(n_3051)
);

AOI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2687),
.A2(n_2788),
.B1(n_2786),
.B2(n_2935),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2806),
.B(n_2643),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2738),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2946),
.B(n_2588),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2794),
.B(n_2586),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2736),
.B(n_2597),
.Y(n_3057)
);

INVx2_ASAP7_75t_SL g3058 ( 
.A(n_2894),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_2824),
.A2(n_2562),
.B1(n_2563),
.B2(n_2560),
.Y(n_3059)
);

AND2x4_ASAP7_75t_L g3060 ( 
.A(n_2848),
.B(n_2356),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2879),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_L g3062 ( 
.A1(n_2824),
.A2(n_2563),
.B1(n_2591),
.B2(n_2560),
.Y(n_3062)
);

BUFx3_ASAP7_75t_L g3063 ( 
.A(n_2896),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2736),
.B(n_2510),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_2845),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2818),
.B(n_2510),
.Y(n_3066)
);

OAI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_2871),
.A2(n_2386),
.B1(n_2379),
.B2(n_2476),
.Y(n_3067)
);

CKINVDCx14_ASAP7_75t_R g3068 ( 
.A(n_2771),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2741),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2917),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2919),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2818),
.B(n_2510),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2957),
.B(n_2641),
.Y(n_3073)
);

OAI221xp5_ASAP7_75t_L g3074 ( 
.A1(n_2694),
.A2(n_2644),
.B1(n_2532),
.B2(n_2631),
.C(n_2656),
.Y(n_3074)
);

AOI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_2929),
.A2(n_2368),
.B(n_2478),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2881),
.A2(n_2591),
.B1(n_2613),
.B2(n_2612),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_2923),
.B(n_2620),
.Y(n_3077)
);

OR2x6_ASAP7_75t_L g3078 ( 
.A(n_2844),
.B(n_2460),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2687),
.B(n_2598),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2689),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_SL g3081 ( 
.A(n_2758),
.B(n_2477),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2848),
.B(n_2620),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2747),
.Y(n_3083)
);

AOI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2687),
.A2(n_2443),
.B1(n_2631),
.B2(n_2328),
.Y(n_3084)
);

BUFx6f_ASAP7_75t_L g3085 ( 
.A(n_2670),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2845),
.B(n_2598),
.Y(n_3086)
);

NAND2xp33_ASAP7_75t_L g3087 ( 
.A(n_2718),
.B(n_2405),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2860),
.B(n_2599),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2860),
.B(n_2599),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2698),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2842),
.B(n_2540),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2694),
.B(n_2541),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2754),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2755),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_SL g3095 ( 
.A(n_2848),
.B(n_2620),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2773),
.Y(n_3096)
);

A2O1A1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2939),
.A2(n_2378),
.B(n_2573),
.C(n_2571),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2887),
.B(n_2620),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2701),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2710),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2713),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2722),
.B(n_2476),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2750),
.B(n_2541),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2722),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2750),
.B(n_2618),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2742),
.B(n_2618),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_2768),
.B(n_2641),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2742),
.B(n_2623),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2881),
.A2(n_2623),
.B1(n_2626),
.B2(n_2656),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2777),
.B(n_2626),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_2939),
.B(n_2476),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2887),
.B(n_2477),
.Y(n_3112)
);

INVx4_ASAP7_75t_L g3113 ( 
.A(n_2844),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2887),
.B(n_2477),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2895),
.B(n_2569),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2714),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_2925),
.B(n_2646),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_SL g3118 ( 
.A(n_2895),
.B(n_2569),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2728),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2778),
.B(n_2646),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2897),
.B(n_2644),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2948),
.B(n_2551),
.Y(n_3122)
);

NOR2x2_ASAP7_75t_L g3123 ( 
.A(n_2756),
.B(n_2653),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2948),
.B(n_2551),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2780),
.B(n_2421),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2889),
.B(n_2653),
.Y(n_3126)
);

NOR2xp67_ASAP7_75t_L g3127 ( 
.A(n_2924),
.B(n_2451),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2844),
.Y(n_3128)
);

NAND2xp33_ASAP7_75t_L g3129 ( 
.A(n_2718),
.B(n_2405),
.Y(n_3129)
);

NAND2x1p5_ASAP7_75t_L g3130 ( 
.A(n_2870),
.B(n_2426),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2781),
.B(n_2421),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2904),
.Y(n_3132)
);

OR2x2_ASAP7_75t_L g3133 ( 
.A(n_2784),
.B(n_2454),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2812),
.B(n_2953),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_SL g3135 ( 
.A(n_2915),
.B(n_2451),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2789),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2796),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2743),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2893),
.B(n_2657),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2797),
.Y(n_3140)
);

NAND2xp33_ASAP7_75t_L g3141 ( 
.A(n_2841),
.B(n_2405),
.Y(n_3141)
);

NAND2x1_ASAP7_75t_L g3142 ( 
.A(n_2870),
.B(n_2888),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2898),
.B(n_2657),
.Y(n_3143)
);

INVx3_ASAP7_75t_L g3144 ( 
.A(n_2888),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2744),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2901),
.B(n_2545),
.Y(n_3146)
);

OR2x2_ASAP7_75t_L g3147 ( 
.A(n_2903),
.B(n_2484),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2884),
.A2(n_2478),
.B(n_2462),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2910),
.B(n_2473),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2745),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2911),
.B(n_2479),
.Y(n_3151)
);

OAI22xp5_ASAP7_75t_SL g3152 ( 
.A1(n_2770),
.A2(n_2338),
.B1(n_2621),
.B2(n_2488),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2913),
.B(n_2914),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2916),
.B(n_2663),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2918),
.B(n_2507),
.Y(n_3155)
);

INVx2_ASAP7_75t_SL g3156 ( 
.A(n_2920),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2746),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2800),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_SL g3159 ( 
.A(n_2915),
.B(n_2691),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2801),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_SL g3161 ( 
.A(n_2895),
.B(n_2569),
.Y(n_3161)
);

BUFx5_ASAP7_75t_L g3162 ( 
.A(n_2764),
.Y(n_3162)
);

AND2x4_ASAP7_75t_SL g3163 ( 
.A(n_2906),
.B(n_2952),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2802),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_2868),
.B(n_2488),
.Y(n_3165)
);

A2O1A1Ixp33_ASAP7_75t_L g3166 ( 
.A1(n_2809),
.A2(n_2336),
.B(n_2508),
.C(n_2606),
.Y(n_3166)
);

AND2x4_ASAP7_75t_SL g3167 ( 
.A(n_2906),
.B(n_2426),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2752),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2770),
.A2(n_2428),
.B1(n_2596),
.B2(n_2590),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2763),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_L g3171 ( 
.A(n_2921),
.B(n_2590),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2774),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2775),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2927),
.B(n_2468),
.Y(n_3174)
);

CKINVDCx5p33_ASAP7_75t_R g3175 ( 
.A(n_2868),
.Y(n_3175)
);

BUFx3_ASAP7_75t_L g3176 ( 
.A(n_2779),
.Y(n_3176)
);

INVx2_ASAP7_75t_SL g3177 ( 
.A(n_2779),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2791),
.Y(n_3178)
);

O2A1O1Ixp5_ASAP7_75t_L g3179 ( 
.A1(n_2811),
.A2(n_2462),
.B(n_2546),
.C(n_2640),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2928),
.B(n_2596),
.Y(n_3180)
);

OR2x2_ASAP7_75t_L g3181 ( 
.A(n_2938),
.B(n_2484),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2940),
.B(n_2567),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_3012),
.Y(n_3183)
);

NAND3xp33_ASAP7_75t_SL g3184 ( 
.A(n_2996),
.B(n_2950),
.C(n_2790),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3153),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2971),
.Y(n_3186)
);

CKINVDCx5p33_ASAP7_75t_R g3187 ( 
.A(n_3175),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_2965),
.A2(n_2666),
.B1(n_2706),
.B2(n_2891),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2972),
.Y(n_3189)
);

BUFx4f_ASAP7_75t_L g3190 ( 
.A(n_3078),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2975),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3092),
.B(n_2902),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_3113),
.Y(n_3193)
);

HB1xp67_ASAP7_75t_L g3194 ( 
.A(n_3065),
.Y(n_3194)
);

AOI22xp5_ASAP7_75t_L g3195 ( 
.A1(n_2967),
.A2(n_2706),
.B1(n_2666),
.B2(n_2891),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2983),
.Y(n_3196)
);

BUFx2_ASAP7_75t_L g3197 ( 
.A(n_3039),
.Y(n_3197)
);

INVx5_ASAP7_75t_L g3198 ( 
.A(n_2989),
.Y(n_3198)
);

BUFx6f_ASAP7_75t_L g3199 ( 
.A(n_2989),
.Y(n_3199)
);

OR2x2_ASAP7_75t_L g3200 ( 
.A(n_2979),
.B(n_2634),
.Y(n_3200)
);

OR2x2_ASAP7_75t_SL g3201 ( 
.A(n_3034),
.B(n_2556),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_3107),
.B(n_2907),
.Y(n_3202)
);

AND2x4_ASAP7_75t_L g3203 ( 
.A(n_3060),
.B(n_3078),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2977),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_3024),
.Y(n_3205)
);

INVx1_ASAP7_75t_SL g3206 ( 
.A(n_3031),
.Y(n_3206)
);

BUFx6f_ASAP7_75t_L g3207 ( 
.A(n_2989),
.Y(n_3207)
);

BUFx2_ASAP7_75t_L g3208 ( 
.A(n_3031),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2984),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3007),
.Y(n_3210)
);

INVxp67_ASAP7_75t_L g3211 ( 
.A(n_3104),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3025),
.Y(n_3212)
);

CKINVDCx5p33_ASAP7_75t_R g3213 ( 
.A(n_3068),
.Y(n_3213)
);

CKINVDCx8_ASAP7_75t_R g3214 ( 
.A(n_3048),
.Y(n_3214)
);

OR2x6_ASAP7_75t_SL g3215 ( 
.A(n_2995),
.B(n_3079),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_3052),
.B(n_2627),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3015),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2988),
.B(n_2627),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3023),
.Y(n_3219)
);

BUFx6f_ASAP7_75t_L g3220 ( 
.A(n_2989),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_3060),
.B(n_2756),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_3035),
.Y(n_3222)
);

INVx3_ASAP7_75t_L g3223 ( 
.A(n_3113),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3051),
.B(n_2902),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3037),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_3061),
.Y(n_3226)
);

AO22x1_ASAP7_75t_L g3227 ( 
.A1(n_3165),
.A2(n_3026),
.B1(n_2967),
.B2(n_2980),
.Y(n_3227)
);

INVx2_ASAP7_75t_SL g3228 ( 
.A(n_3063),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3070),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2965),
.B(n_2826),
.Y(n_3230)
);

AND2x6_ASAP7_75t_L g3231 ( 
.A(n_2959),
.B(n_2542),
.Y(n_3231)
);

INVx4_ASAP7_75t_L g3232 ( 
.A(n_3078),
.Y(n_3232)
);

INVx6_ASAP7_75t_L g3233 ( 
.A(n_3030),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3033),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_2976),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_3071),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_3182),
.B(n_2691),
.Y(n_3237)
);

BUFx6f_ASAP7_75t_L g3238 ( 
.A(n_3085),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_2980),
.B(n_2785),
.Y(n_3239)
);

BUFx2_ASAP7_75t_L g3240 ( 
.A(n_3104),
.Y(n_3240)
);

BUFx3_ASAP7_75t_L g3241 ( 
.A(n_2985),
.Y(n_3241)
);

INVx2_ASAP7_75t_SL g3242 ( 
.A(n_3013),
.Y(n_3242)
);

AND2x4_ASAP7_75t_L g3243 ( 
.A(n_3128),
.B(n_2756),
.Y(n_3243)
);

INVx1_ASAP7_75t_SL g3244 ( 
.A(n_3133),
.Y(n_3244)
);

OR2x2_ASAP7_75t_L g3245 ( 
.A(n_2961),
.B(n_2790),
.Y(n_3245)
);

NOR2xp33_ASAP7_75t_R g3246 ( 
.A(n_3159),
.B(n_2556),
.Y(n_3246)
);

O2A1O1Ixp33_ASAP7_75t_L g3247 ( 
.A1(n_3074),
.A2(n_2949),
.B(n_2606),
.C(n_2568),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2965),
.B(n_2826),
.Y(n_3248)
);

BUFx3_ASAP7_75t_L g3249 ( 
.A(n_3058),
.Y(n_3249)
);

NOR2xp33_ASAP7_75t_L g3250 ( 
.A(n_3043),
.B(n_3026),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3040),
.Y(n_3251)
);

INVx2_ASAP7_75t_SL g3252 ( 
.A(n_3156),
.Y(n_3252)
);

INVx2_ASAP7_75t_SL g3253 ( 
.A(n_2974),
.Y(n_3253)
);

NOR2xp33_ASAP7_75t_SL g3254 ( 
.A(n_3081),
.B(n_2841),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_3043),
.B(n_3117),
.Y(n_3255)
);

INVxp67_ASAP7_75t_L g3256 ( 
.A(n_3049),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_3176),
.Y(n_3257)
);

AOI22xp5_ASAP7_75t_L g3258 ( 
.A1(n_3005),
.A2(n_2727),
.B1(n_2949),
.B2(n_2761),
.Y(n_3258)
);

INVx2_ASAP7_75t_SL g3259 ( 
.A(n_3030),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3041),
.Y(n_3260)
);

HB1xp67_ASAP7_75t_L g3261 ( 
.A(n_3065),
.Y(n_3261)
);

OR2x2_ASAP7_75t_L g3262 ( 
.A(n_2998),
.B(n_2640),
.Y(n_3262)
);

BUFx2_ASAP7_75t_L g3263 ( 
.A(n_3121),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2965),
.B(n_2829),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2999),
.Y(n_3265)
);

AND2x4_ASAP7_75t_L g3266 ( 
.A(n_3128),
.B(n_2944),
.Y(n_3266)
);

HB1xp67_ASAP7_75t_L g3267 ( 
.A(n_3102),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3046),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2965),
.B(n_2829),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3020),
.B(n_2864),
.Y(n_3270)
);

INVxp67_ASAP7_75t_SL g3271 ( 
.A(n_3011),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3073),
.B(n_2727),
.Y(n_3272)
);

A2O1A1Ixp33_ASAP7_75t_L g3273 ( 
.A1(n_3148),
.A2(n_2947),
.B(n_2956),
.C(n_2866),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3054),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3003),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3069),
.Y(n_3276)
);

AOI22x1_ASAP7_75t_L g3277 ( 
.A1(n_3148),
.A2(n_2941),
.B1(n_2426),
.B2(n_2543),
.Y(n_3277)
);

INVx3_ASAP7_75t_SL g3278 ( 
.A(n_3123),
.Y(n_3278)
);

AND2x4_ASAP7_75t_L g3279 ( 
.A(n_3115),
.B(n_2944),
.Y(n_3279)
);

AOI22xp5_ASAP7_75t_L g3280 ( 
.A1(n_3005),
.A2(n_2941),
.B1(n_2798),
.B2(n_2417),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_3085),
.Y(n_3281)
);

BUFx2_ASAP7_75t_L g3282 ( 
.A(n_3147),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3083),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3020),
.B(n_2864),
.Y(n_3284)
);

BUFx4f_ASAP7_75t_L g3285 ( 
.A(n_3085),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_3010),
.Y(n_3286)
);

AOI211xp5_ASAP7_75t_L g3287 ( 
.A1(n_3152),
.A2(n_2508),
.B(n_2546),
.C(n_2457),
.Y(n_3287)
);

INVx5_ASAP7_75t_L g3288 ( 
.A(n_3085),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3080),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3093),
.Y(n_3290)
);

INVx5_ASAP7_75t_L g3291 ( 
.A(n_2992),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3094),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3096),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3090),
.Y(n_3294)
);

INVx3_ASAP7_75t_L g3295 ( 
.A(n_2978),
.Y(n_3295)
);

AND2x4_ASAP7_75t_L g3296 ( 
.A(n_3118),
.B(n_2944),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3103),
.B(n_2807),
.Y(n_3297)
);

NOR2xp67_ASAP7_75t_L g3298 ( 
.A(n_3155),
.B(n_2926),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3099),
.Y(n_3299)
);

INVx3_ASAP7_75t_SL g3300 ( 
.A(n_3181),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_3100),
.Y(n_3301)
);

INVx2_ASAP7_75t_SL g3302 ( 
.A(n_3177),
.Y(n_3302)
);

CKINVDCx5p33_ASAP7_75t_R g3303 ( 
.A(n_3009),
.Y(n_3303)
);

INVxp67_ASAP7_75t_L g3304 ( 
.A(n_3049),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3110),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_3050),
.B(n_2659),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3139),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3105),
.B(n_2810),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_3084),
.B(n_2659),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_3101),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3116),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3119),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3143),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3138),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_2978),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3038),
.B(n_2813),
.Y(n_3316)
);

CKINVDCx20_ASAP7_75t_R g3317 ( 
.A(n_2960),
.Y(n_3317)
);

INVx2_ASAP7_75t_SL g3318 ( 
.A(n_3163),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3145),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_3161),
.B(n_2952),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_3112),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3038),
.B(n_2814),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3150),
.Y(n_3323)
);

BUFx6f_ASAP7_75t_L g3324 ( 
.A(n_3114),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3136),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_3169),
.Y(n_3326)
);

AOI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_2981),
.A2(n_2798),
.B1(n_2417),
.B2(n_2648),
.Y(n_3327)
);

BUFx6f_ASAP7_75t_L g3328 ( 
.A(n_3082),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3137),
.Y(n_3329)
);

BUFx3_ASAP7_75t_L g3330 ( 
.A(n_3053),
.Y(n_3330)
);

NOR2xp67_ASAP7_75t_L g3331 ( 
.A(n_2992),
.B(n_2926),
.Y(n_3331)
);

AND2x4_ASAP7_75t_L g3332 ( 
.A(n_3032),
.B(n_2952),
.Y(n_3332)
);

CKINVDCx5p33_ASAP7_75t_R g3333 ( 
.A(n_3132),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3122),
.B(n_2815),
.Y(n_3334)
);

BUFx4f_ASAP7_75t_L g3335 ( 
.A(n_3130),
.Y(n_3335)
);

BUFx3_ASAP7_75t_L g3336 ( 
.A(n_3053),
.Y(n_3336)
);

INVx2_ASAP7_75t_SL g3337 ( 
.A(n_3077),
.Y(n_3337)
);

BUFx6f_ASAP7_75t_L g3338 ( 
.A(n_3095),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_3098),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3122),
.B(n_2817),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3140),
.Y(n_3341)
);

AOI22xp33_ASAP7_75t_L g3342 ( 
.A1(n_3017),
.A2(n_2659),
.B1(n_2417),
.B2(n_2543),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3157),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3158),
.Y(n_3344)
);

AND2x4_ASAP7_75t_L g3345 ( 
.A(n_3055),
.B(n_2358),
.Y(n_3345)
);

NAND3xp33_ASAP7_75t_L g3346 ( 
.A(n_2981),
.B(n_2632),
.C(n_2582),
.Y(n_3346)
);

HB1xp67_ASAP7_75t_L g3347 ( 
.A(n_3102),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3168),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3170),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3172),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3160),
.Y(n_3351)
);

HB1xp67_ASAP7_75t_L g3352 ( 
.A(n_3132),
.Y(n_3352)
);

AND2x6_ASAP7_75t_SL g3353 ( 
.A(n_3126),
.B(n_2453),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_3029),
.B(n_2936),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_3047),
.B(n_2785),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3057),
.Y(n_3356)
);

BUFx2_ASAP7_75t_L g3357 ( 
.A(n_2993),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3164),
.Y(n_3358)
);

INVx5_ASAP7_75t_L g3359 ( 
.A(n_3144),
.Y(n_3359)
);

AND2x4_ASAP7_75t_L g3360 ( 
.A(n_3127),
.B(n_2358),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_2963),
.B(n_2556),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_3017),
.A2(n_2542),
.B1(n_2648),
.B2(n_2576),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3173),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3124),
.B(n_2819),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2969),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_3134),
.B(n_2890),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3022),
.A2(n_3067),
.B1(n_3111),
.B2(n_2964),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_2970),
.B(n_2556),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3178),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_2973),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2991),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2987),
.B(n_2418),
.Y(n_3372)
);

HB1xp67_ASAP7_75t_L g3373 ( 
.A(n_3106),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3018),
.Y(n_3374)
);

INVx5_ASAP7_75t_L g3375 ( 
.A(n_3144),
.Y(n_3375)
);

BUFx6f_ASAP7_75t_L g3376 ( 
.A(n_3006),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_3146),
.Y(n_3377)
);

BUFx2_ASAP7_75t_L g3378 ( 
.A(n_3126),
.Y(n_3378)
);

AND2x2_ASAP7_75t_SL g3379 ( 
.A(n_3044),
.B(n_2890),
.Y(n_3379)
);

BUFx8_ASAP7_75t_L g3380 ( 
.A(n_3162),
.Y(n_3380)
);

HB1xp67_ASAP7_75t_L g3381 ( 
.A(n_3000),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_2964),
.B(n_2936),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3124),
.B(n_2823),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3086),
.Y(n_3384)
);

INVxp67_ASAP7_75t_SL g3385 ( 
.A(n_3021),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3088),
.Y(n_3386)
);

INVx2_ASAP7_75t_SL g3387 ( 
.A(n_3167),
.Y(n_3387)
);

BUFx6f_ASAP7_75t_L g3388 ( 
.A(n_3130),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3111),
.B(n_3097),
.Y(n_3389)
);

NOR2x1_ASAP7_75t_SL g3390 ( 
.A(n_3001),
.B(n_2841),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3021),
.B(n_2827),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_2966),
.B(n_2828),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3377),
.B(n_2966),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_3255),
.B(n_2418),
.Y(n_3394)
);

OA22x2_ASAP7_75t_L g3395 ( 
.A1(n_3195),
.A2(n_3045),
.B1(n_3036),
.B2(n_3108),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_3373),
.B(n_3120),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_3273),
.A2(n_3141),
.B(n_3129),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3250),
.B(n_3014),
.Y(n_3398)
);

AOI33xp33_ASAP7_75t_L g3399 ( 
.A1(n_3188),
.A2(n_3109),
.A3(n_3076),
.B1(n_3059),
.B2(n_3062),
.B3(n_2723),
.Y(n_3399)
);

O2A1O1Ixp33_ASAP7_75t_L g3400 ( 
.A1(n_3184),
.A2(n_2962),
.B(n_2994),
.C(n_2968),
.Y(n_3400)
);

NAND3xp33_ASAP7_75t_L g3401 ( 
.A(n_3287),
.B(n_3166),
.C(n_3154),
.Y(n_3401)
);

O2A1O1Ixp33_ASAP7_75t_L g3402 ( 
.A1(n_3184),
.A2(n_3027),
.B(n_2986),
.C(n_2990),
.Y(n_3402)
);

O2A1O1Ixp5_ASAP7_75t_L g3403 ( 
.A1(n_3237),
.A2(n_3179),
.B(n_3002),
.C(n_3075),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_SL g3404 ( 
.A(n_3321),
.B(n_3324),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3202),
.B(n_3000),
.Y(n_3405)
);

OAI22xp5_ASAP7_75t_L g3406 ( 
.A1(n_3258),
.A2(n_3109),
.B1(n_3076),
.B2(n_3059),
.Y(n_3406)
);

AND2x4_ASAP7_75t_SL g3407 ( 
.A(n_3360),
.B(n_2779),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_3321),
.B(n_3008),
.Y(n_3408)
);

INVxp67_ASAP7_75t_L g3409 ( 
.A(n_3282),
.Y(n_3409)
);

AND2x6_ASAP7_75t_L g3410 ( 
.A(n_3327),
.B(n_3280),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3194),
.Y(n_3411)
);

AOI33xp33_ASAP7_75t_L g3412 ( 
.A1(n_3195),
.A2(n_3062),
.A3(n_2529),
.B1(n_2625),
.B2(n_2619),
.B3(n_93),
.Y(n_3412)
);

A2O1A1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_3247),
.A2(n_3075),
.B(n_3042),
.C(n_3179),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_SL g3414 ( 
.A(n_3321),
.B(n_3019),
.Y(n_3414)
);

OAI22xp5_ASAP7_75t_L g3415 ( 
.A1(n_3258),
.A2(n_2453),
.B1(n_3028),
.B2(n_3091),
.Y(n_3415)
);

A2O1A1Ixp33_ASAP7_75t_L g3416 ( 
.A1(n_3247),
.A2(n_3042),
.B(n_3002),
.C(n_3171),
.Y(n_3416)
);

NOR3xp33_ASAP7_75t_L g3417 ( 
.A(n_3227),
.B(n_2982),
.C(n_3149),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3263),
.B(n_3016),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3374),
.B(n_3016),
.Y(n_3419)
);

OAI22xp5_ASAP7_75t_SL g3420 ( 
.A1(n_3326),
.A2(n_2453),
.B1(n_3180),
.B2(n_3171),
.Y(n_3420)
);

OAI21xp33_ASAP7_75t_L g3421 ( 
.A1(n_3367),
.A2(n_3135),
.B(n_3180),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3324),
.B(n_2899),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_3324),
.B(n_2905),
.Y(n_3423)
);

AOI22xp33_ASAP7_75t_L g3424 ( 
.A1(n_3355),
.A2(n_2576),
.B1(n_2759),
.B2(n_2753),
.Y(n_3424)
);

A2O1A1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_3287),
.A2(n_3087),
.B(n_2997),
.C(n_2866),
.Y(n_3425)
);

NOR3xp33_ASAP7_75t_L g3426 ( 
.A(n_3366),
.B(n_3174),
.C(n_3151),
.Y(n_3426)
);

NAND2xp33_ASAP7_75t_SL g3427 ( 
.A(n_3246),
.B(n_2783),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_3367),
.B(n_3064),
.Y(n_3428)
);

AOI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_3346),
.A2(n_3004),
.B(n_2578),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3265),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3300),
.B(n_3066),
.Y(n_3431)
);

OAI21xp33_ASAP7_75t_L g3432 ( 
.A1(n_3280),
.A2(n_3056),
.B(n_3072),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3370),
.B(n_3089),
.Y(n_3433)
);

INVxp67_ASAP7_75t_L g3434 ( 
.A(n_3197),
.Y(n_3434)
);

NOR2xp67_ASAP7_75t_L g3435 ( 
.A(n_3187),
.B(n_3253),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3239),
.B(n_2783),
.Y(n_3436)
);

OAI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3309),
.A2(n_2544),
.B1(n_3131),
.B2(n_3125),
.Y(n_3437)
);

BUFx6f_ASAP7_75t_L g3438 ( 
.A(n_3285),
.Y(n_3438)
);

INVx4_ASAP7_75t_L g3439 ( 
.A(n_3198),
.Y(n_3439)
);

NAND3xp33_ASAP7_75t_SL g3440 ( 
.A(n_3214),
.B(n_2327),
.C(n_2632),
.Y(n_3440)
);

BUFx4f_ASAP7_75t_L g3441 ( 
.A(n_3243),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3194),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3346),
.A2(n_3271),
.B(n_3254),
.Y(n_3443)
);

INVx3_ASAP7_75t_L g3444 ( 
.A(n_3388),
.Y(n_3444)
);

O2A1O1Ixp33_ASAP7_75t_L g3445 ( 
.A1(n_3216),
.A2(n_2847),
.B(n_2658),
.C(n_2654),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3357),
.B(n_2831),
.Y(n_3446)
);

OAI22x1_ASAP7_75t_L g3447 ( 
.A1(n_3277),
.A2(n_2937),
.B1(n_2834),
.B2(n_2856),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3275),
.Y(n_3448)
);

OR2x6_ASAP7_75t_SL g3449 ( 
.A(n_3213),
.B(n_2649),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3261),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3306),
.B(n_3317),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3185),
.B(n_2832),
.Y(n_3452)
);

O2A1O1Ixp33_ASAP7_75t_L g3453 ( 
.A1(n_3278),
.A2(n_2658),
.B(n_2578),
.C(n_2570),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3384),
.B(n_2857),
.Y(n_3454)
);

BUFx2_ASAP7_75t_L g3455 ( 
.A(n_3333),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3386),
.B(n_3356),
.Y(n_3456)
);

INVx3_ASAP7_75t_L g3457 ( 
.A(n_3388),
.Y(n_3457)
);

NOR2x1_ASAP7_75t_L g3458 ( 
.A(n_3330),
.B(n_3142),
.Y(n_3458)
);

CKINVDCx14_ASAP7_75t_R g3459 ( 
.A(n_3183),
.Y(n_3459)
);

BUFx6f_ASAP7_75t_L g3460 ( 
.A(n_3285),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3271),
.A2(n_2803),
.B(n_2493),
.Y(n_3461)
);

NOR3xp33_ASAP7_75t_L g3462 ( 
.A(n_3361),
.B(n_2759),
.C(n_2753),
.Y(n_3462)
);

INVx3_ASAP7_75t_L g3463 ( 
.A(n_3388),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_L g3464 ( 
.A(n_3303),
.B(n_2783),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3286),
.Y(n_3465)
);

BUFx3_ASAP7_75t_L g3466 ( 
.A(n_3257),
.Y(n_3466)
);

A2O1A1Ixp33_ASAP7_75t_L g3467 ( 
.A1(n_3327),
.A2(n_2363),
.B(n_2776),
.C(n_2493),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3186),
.Y(n_3468)
);

OAI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_3362),
.A2(n_2544),
.B1(n_2909),
.B2(n_2820),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3261),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3254),
.A2(n_2803),
.B(n_2482),
.Y(n_3471)
);

INVxp67_ASAP7_75t_L g3472 ( 
.A(n_3208),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3371),
.B(n_3244),
.Y(n_3473)
);

OR2x6_ASAP7_75t_L g3474 ( 
.A(n_3232),
.B(n_2846),
.Y(n_3474)
);

A2O1A1Ixp33_ASAP7_75t_L g3475 ( 
.A1(n_3218),
.A2(n_2363),
.B(n_2776),
.C(n_2482),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_3390),
.A2(n_2495),
.B(n_2883),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_3224),
.A2(n_2495),
.B(n_2883),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3244),
.B(n_2859),
.Y(n_3478)
);

O2A1O1Ixp33_ASAP7_75t_L g3479 ( 
.A1(n_3389),
.A2(n_2575),
.B(n_2595),
.C(n_2566),
.Y(n_3479)
);

NAND2x1p5_ASAP7_75t_L g3480 ( 
.A(n_3190),
.B(n_2683),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3342),
.A2(n_2576),
.B1(n_2648),
.B2(n_2502),
.Y(n_3481)
);

INVxp67_ASAP7_75t_L g3482 ( 
.A(n_3378),
.Y(n_3482)
);

BUFx2_ASAP7_75t_L g3483 ( 
.A(n_3336),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3305),
.B(n_2861),
.Y(n_3484)
);

A2O1A1Ixp33_ASAP7_75t_L g3485 ( 
.A1(n_3368),
.A2(n_2363),
.B(n_2384),
.C(n_2565),
.Y(n_3485)
);

OR2x6_ASAP7_75t_SL g3486 ( 
.A(n_3389),
.B(n_2676),
.Y(n_3486)
);

OR2x6_ASAP7_75t_SL g3487 ( 
.A(n_3245),
.B(n_2676),
.Y(n_3487)
);

NOR2xp33_ASAP7_75t_L g3488 ( 
.A(n_3201),
.B(n_2787),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3272),
.B(n_2816),
.Y(n_3489)
);

O2A1O1Ixp33_ASAP7_75t_L g3490 ( 
.A1(n_3256),
.A2(n_2604),
.B(n_2419),
.C(n_2414),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3307),
.B(n_2862),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3382),
.B(n_3259),
.Y(n_3492)
);

O2A1O1Ixp5_ASAP7_75t_L g3493 ( 
.A1(n_3224),
.A2(n_2647),
.B(n_2757),
.C(n_2717),
.Y(n_3493)
);

OAI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3298),
.A2(n_2502),
.B(n_2717),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_3376),
.B(n_2569),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3189),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3313),
.B(n_3354),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3192),
.A2(n_2825),
.B(n_2459),
.Y(n_3498)
);

A2O1A1Ixp33_ASAP7_75t_L g3499 ( 
.A1(n_3190),
.A2(n_3372),
.B(n_3298),
.C(n_3262),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3381),
.B(n_2869),
.Y(n_3500)
);

OAI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3256),
.A2(n_2544),
.B1(n_2820),
.B2(n_2787),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3204),
.Y(n_3502)
);

AOI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3345),
.A2(n_2648),
.B1(n_2638),
.B2(n_2912),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3376),
.B(n_2787),
.Y(n_3504)
);

AO21x1_ASAP7_75t_L g3505 ( 
.A1(n_3385),
.A2(n_2875),
.B(n_2702),
.Y(n_3505)
);

O2A1O1Ixp5_ASAP7_75t_L g3506 ( 
.A1(n_3192),
.A2(n_2757),
.B(n_2767),
.C(n_2392),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3205),
.Y(n_3507)
);

AOI21x1_ASAP7_75t_L g3508 ( 
.A1(n_3331),
.A2(n_2767),
.B(n_2395),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3335),
.A2(n_2459),
.B(n_2483),
.Y(n_3509)
);

OAI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3304),
.A2(n_2820),
.B1(n_2846),
.B2(n_2456),
.Y(n_3510)
);

NOR2x1_ASAP7_75t_L g3511 ( 
.A(n_3193),
.B(n_2846),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_SL g3512 ( 
.A(n_3376),
.B(n_2912),
.Y(n_3512)
);

O2A1O1Ixp33_ASAP7_75t_L g3513 ( 
.A1(n_3304),
.A2(n_2353),
.B(n_2365),
.C(n_2352),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3352),
.B(n_2799),
.Y(n_3514)
);

BUFx6f_ASAP7_75t_L g3515 ( 
.A(n_3241),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3373),
.B(n_2804),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3335),
.A2(n_2398),
.B(n_2873),
.Y(n_3517)
);

OA22x2_ASAP7_75t_L g3518 ( 
.A1(n_3267),
.A2(n_2930),
.B1(n_2686),
.B2(n_2700),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3206),
.B(n_2822),
.Y(n_3519)
);

O2A1O1Ixp33_ASAP7_75t_L g3520 ( 
.A1(n_3337),
.A2(n_2389),
.B(n_2391),
.C(n_2371),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3206),
.B(n_2837),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3233),
.B(n_2323),
.Y(n_3522)
);

NOR3xp33_ASAP7_75t_L g3523 ( 
.A(n_3200),
.B(n_2686),
.C(n_2677),
.Y(n_3523)
);

INVxp67_ASAP7_75t_L g3524 ( 
.A(n_3240),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3347),
.B(n_2839),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3392),
.B(n_2850),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_3379),
.B(n_3162),
.Y(n_3527)
);

O2A1O1Ixp33_ASAP7_75t_L g3528 ( 
.A1(n_3392),
.A2(n_2865),
.B(n_2908),
.C(n_2852),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_L g3529 ( 
.A(n_3233),
.B(n_2323),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_3228),
.B(n_2677),
.Y(n_3530)
);

BUFx2_ASAP7_75t_L g3531 ( 
.A(n_3221),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3211),
.B(n_2684),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3385),
.A2(n_2882),
.B1(n_2877),
.B2(n_2425),
.Y(n_3533)
);

OAI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_3270),
.A2(n_2877),
.B1(n_2425),
.B2(n_2655),
.Y(n_3534)
);

OAI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3215),
.A2(n_2461),
.B1(n_2930),
.B2(n_2601),
.Y(n_3535)
);

OR2x6_ASAP7_75t_SL g3536 ( 
.A(n_3230),
.B(n_2467),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3221),
.B(n_2808),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3212),
.Y(n_3538)
);

OAI22xp5_ASAP7_75t_L g3539 ( 
.A1(n_3230),
.A2(n_2610),
.B1(n_2821),
.B2(n_2700),
.Y(n_3539)
);

INVxp67_ASAP7_75t_L g3540 ( 
.A(n_3235),
.Y(n_3540)
);

O2A1O1Ixp33_ASAP7_75t_L g3541 ( 
.A1(n_3211),
.A2(n_2852),
.B(n_2908),
.C(n_2865),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3248),
.A2(n_2958),
.B(n_2933),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3191),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3196),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3328),
.B(n_3162),
.Y(n_3545)
);

NOR2xp33_ASAP7_75t_R g3546 ( 
.A(n_3318),
.B(n_2670),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3248),
.A2(n_2958),
.B(n_2933),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3369),
.B(n_2684),
.Y(n_3548)
);

O2A1O1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_3270),
.A2(n_2821),
.B(n_2836),
.C(n_2808),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_3209),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3210),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3334),
.B(n_2502),
.Y(n_3552)
);

INVxp33_ASAP7_75t_SL g3553 ( 
.A(n_3249),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3334),
.B(n_2502),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3345),
.B(n_2836),
.Y(n_3555)
);

O2A1O1Ixp5_ASAP7_75t_L g3556 ( 
.A1(n_3264),
.A2(n_2530),
.B(n_2922),
.C(n_2833),
.Y(n_3556)
);

O2A1O1Ixp5_ASAP7_75t_L g3557 ( 
.A1(n_3264),
.A2(n_2530),
.B(n_2922),
.C(n_2833),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3231),
.A2(n_2576),
.B1(n_2648),
.B2(n_2502),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3203),
.B(n_2853),
.Y(n_3559)
);

OAI21x1_ASAP7_75t_L g3560 ( 
.A1(n_3269),
.A2(n_2843),
.B(n_2835),
.Y(n_3560)
);

AND2x4_ASAP7_75t_L g3561 ( 
.A(n_3203),
.B(n_2682),
.Y(n_3561)
);

BUFx6f_ASAP7_75t_L g3562 ( 
.A(n_3199),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_3217),
.Y(n_3563)
);

AOI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3231),
.A2(n_2576),
.B1(n_2648),
.B2(n_2502),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_3269),
.A2(n_2843),
.B(n_2835),
.Y(n_3565)
);

AOI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3284),
.A2(n_2876),
.B(n_2867),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3340),
.B(n_2943),
.Y(n_3567)
);

AOI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3231),
.A2(n_2638),
.B1(n_2576),
.B2(n_2853),
.Y(n_3568)
);

AOI22xp33_ASAP7_75t_L g3569 ( 
.A1(n_3231),
.A2(n_2638),
.B1(n_2405),
.B2(n_2892),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_3199),
.Y(n_3570)
);

INVx8_ASAP7_75t_L g3571 ( 
.A(n_3198),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_SL g3572 ( 
.A1(n_3360),
.A2(n_2702),
.B1(n_2721),
.B2(n_2683),
.Y(n_3572)
);

AO221x1_ASAP7_75t_L g3573 ( 
.A1(n_3328),
.A2(n_2724),
.B1(n_2726),
.B2(n_2716),
.C(n_2682),
.Y(n_3573)
);

O2A1O1Ixp33_ASAP7_75t_L g3574 ( 
.A1(n_3284),
.A2(n_2954),
.B(n_2943),
.C(n_2343),
.Y(n_3574)
);

AOI221xp5_ASAP7_75t_L g3575 ( 
.A1(n_3365),
.A2(n_2506),
.B1(n_2942),
.B2(n_2496),
.C(n_2900),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3219),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3234),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3340),
.B(n_2954),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3297),
.A2(n_2876),
.B(n_2867),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_3297),
.A2(n_2735),
.B(n_2405),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3308),
.A2(n_2735),
.B(n_2405),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3308),
.A2(n_2735),
.B(n_3162),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_3331),
.A2(n_3162),
.B(n_2942),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_3242),
.B(n_2682),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3391),
.A2(n_3162),
.B(n_2840),
.Y(n_3585)
);

BUFx2_ASAP7_75t_L g3586 ( 
.A(n_3199),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3391),
.A2(n_2840),
.B(n_2892),
.Y(n_3587)
);

A2O1A1Ixp33_ASAP7_75t_L g3588 ( 
.A1(n_3316),
.A2(n_3322),
.B(n_3383),
.C(n_3364),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3364),
.A2(n_2900),
.B(n_2651),
.Y(n_3589)
);

OA22x2_ASAP7_75t_L g3590 ( 
.A1(n_3383),
.A2(n_2721),
.B1(n_2517),
.B2(n_2496),
.Y(n_3590)
);

NOR2xp33_ASAP7_75t_L g3591 ( 
.A(n_3252),
.B(n_2716),
.Y(n_3591)
);

BUFx3_ASAP7_75t_L g3592 ( 
.A(n_3207),
.Y(n_3592)
);

BUFx2_ASAP7_75t_L g3593 ( 
.A(n_3207),
.Y(n_3593)
);

NOR2xp67_ASAP7_75t_L g3594 ( 
.A(n_3387),
.B(n_3222),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3328),
.B(n_2716),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3225),
.B(n_2724),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_3338),
.B(n_2724),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_SL g3598 ( 
.A(n_3338),
.B(n_2726),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3316),
.A2(n_2517),
.B(n_2726),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3322),
.A2(n_2517),
.B(n_2734),
.Y(n_3600)
);

BUFx3_ASAP7_75t_L g3601 ( 
.A(n_3207),
.Y(n_3601)
);

OAI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_3251),
.A2(n_2734),
.B1(n_2740),
.B2(n_2739),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3226),
.B(n_2734),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_3332),
.B(n_2739),
.Y(n_3604)
);

BUFx3_ASAP7_75t_L g3605 ( 
.A(n_3220),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3229),
.B(n_2739),
.Y(n_3606)
);

OA21x2_ASAP7_75t_L g3607 ( 
.A1(n_3403),
.A2(n_3329),
.B(n_3325),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3405),
.B(n_3260),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3497),
.B(n_3268),
.Y(n_3609)
);

NAND3xp33_ASAP7_75t_L g3610 ( 
.A(n_3401),
.B(n_3276),
.C(n_3274),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3456),
.B(n_3283),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3413),
.A2(n_3359),
.B(n_3291),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3426),
.B(n_3243),
.Y(n_3613)
);

NOR2xp33_ASAP7_75t_L g3614 ( 
.A(n_3553),
.B(n_3353),
.Y(n_3614)
);

AOI221xp5_ASAP7_75t_SL g3615 ( 
.A1(n_3421),
.A2(n_3339),
.B1(n_3338),
.B2(n_3344),
.C(n_3341),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3508),
.A2(n_3358),
.B(n_3351),
.Y(n_3616)
);

BUFx12f_ASAP7_75t_L g3617 ( 
.A(n_3515),
.Y(n_3617)
);

INVx3_ASAP7_75t_SL g3618 ( 
.A(n_3515),
.Y(n_3618)
);

OAI21x1_ASAP7_75t_L g3619 ( 
.A1(n_3580),
.A2(n_3315),
.B(n_3295),
.Y(n_3619)
);

OAI21x1_ASAP7_75t_L g3620 ( 
.A1(n_3581),
.A2(n_3582),
.B(n_3476),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3473),
.B(n_3290),
.Y(n_3621)
);

AO31x2_ASAP7_75t_L g3622 ( 
.A1(n_3505),
.A2(n_3232),
.A3(n_3293),
.B(n_3292),
.Y(n_3622)
);

AO31x2_ASAP7_75t_L g3623 ( 
.A1(n_3447),
.A2(n_3236),
.A3(n_3294),
.B(n_3289),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3397),
.A2(n_3359),
.B(n_3291),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_3443),
.A2(n_3359),
.B(n_3291),
.Y(n_3625)
);

NAND2x1p5_ASAP7_75t_L g3626 ( 
.A(n_3458),
.B(n_3511),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3416),
.A2(n_3375),
.B(n_3288),
.Y(n_3627)
);

OAI21x1_ASAP7_75t_SL g3628 ( 
.A1(n_3402),
.A2(n_3301),
.B(n_3299),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3398),
.B(n_3310),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3588),
.B(n_3311),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3543),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3425),
.A2(n_3375),
.B(n_3288),
.Y(n_3632)
);

AOI21x1_ASAP7_75t_L g3633 ( 
.A1(n_3422),
.A2(n_3332),
.B(n_3296),
.Y(n_3633)
);

AOI221xp5_ASAP7_75t_SL g3634 ( 
.A1(n_3406),
.A2(n_3339),
.B1(n_3319),
.B2(n_3323),
.C(n_3314),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_SL g3635 ( 
.A(n_3499),
.B(n_3339),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3409),
.B(n_3312),
.Y(n_3636)
);

NAND2xp33_ASAP7_75t_L g3637 ( 
.A(n_3417),
.B(n_3193),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_SL g3638 ( 
.A(n_3441),
.B(n_3375),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3550),
.Y(n_3639)
);

AO31x2_ASAP7_75t_L g3640 ( 
.A1(n_3534),
.A2(n_3343),
.A3(n_3349),
.B(n_3348),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_SL g3641 ( 
.A1(n_3400),
.A2(n_3363),
.B(n_3350),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3418),
.B(n_3353),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3396),
.B(n_3279),
.Y(n_3643)
);

OAI21x1_ASAP7_75t_L g3644 ( 
.A1(n_3429),
.A2(n_3315),
.B(n_3295),
.Y(n_3644)
);

AOI211x1_ASAP7_75t_L g3645 ( 
.A1(n_3415),
.A2(n_156),
.B(n_168),
.C(n_148),
.Y(n_3645)
);

A2O1A1Ixp33_ASAP7_75t_L g3646 ( 
.A1(n_3399),
.A2(n_3279),
.B(n_3320),
.C(n_3296),
.Y(n_3646)
);

INVx3_ASAP7_75t_L g3647 ( 
.A(n_3444),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3544),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3461),
.A2(n_3223),
.B(n_2496),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3471),
.A2(n_3223),
.B(n_2343),
.Y(n_3650)
);

INVxp67_ASAP7_75t_SL g3651 ( 
.A(n_3563),
.Y(n_3651)
);

OAI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_3401),
.A2(n_2638),
.B(n_3320),
.Y(n_3652)
);

AOI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3509),
.A2(n_3288),
.B(n_3198),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3482),
.B(n_3220),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_L g3655 ( 
.A1(n_3542),
.A2(n_2343),
.B(n_2316),
.Y(n_3655)
);

AO32x2_ASAP7_75t_L g3656 ( 
.A1(n_3420),
.A2(n_3302),
.A3(n_3380),
.B1(n_71),
.B2(n_69),
.Y(n_3656)
);

AOI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_3498),
.A2(n_3266),
.B(n_3380),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3531),
.B(n_3220),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3477),
.A2(n_3266),
.B(n_2760),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3472),
.B(n_3238),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_SL g3661 ( 
.A(n_3441),
.B(n_3238),
.Y(n_3661)
);

OAI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3445),
.A2(n_2638),
.B(n_2439),
.Y(n_3662)
);

A2O1A1Ixp33_ASAP7_75t_L g3663 ( 
.A1(n_3412),
.A2(n_3281),
.B(n_3238),
.C(n_2740),
.Y(n_3663)
);

AO22x2_ASAP7_75t_L g3664 ( 
.A1(n_3411),
.A2(n_3281),
.B1(n_73),
.B2(n_70),
.Y(n_3664)
);

O2A1O1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_3440),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3594),
.B(n_3281),
.Y(n_3666)
);

OAI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3485),
.A2(n_2638),
.B(n_2439),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3524),
.B(n_146),
.Y(n_3668)
);

O2A1O1Ixp5_ASAP7_75t_L g3669 ( 
.A1(n_3494),
.A2(n_2439),
.B(n_2732),
.C(n_2711),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3419),
.B(n_147),
.Y(n_3670)
);

OAI21x1_ASAP7_75t_L g3671 ( 
.A1(n_3547),
.A2(n_2764),
.B(n_2732),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3442),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3393),
.B(n_149),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3558),
.A2(n_2760),
.B(n_2740),
.Y(n_3674)
);

INVx3_ASAP7_75t_L g3675 ( 
.A(n_3444),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3492),
.B(n_2760),
.Y(n_3676)
);

NAND2x1p5_ASAP7_75t_L g3677 ( 
.A(n_3483),
.B(n_2711),
.Y(n_3677)
);

INVx3_ASAP7_75t_L g3678 ( 
.A(n_3457),
.Y(n_3678)
);

INVx3_ASAP7_75t_L g3679 ( 
.A(n_3457),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3450),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3564),
.A2(n_2439),
.B(n_2764),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3517),
.A2(n_2439),
.B(n_2764),
.Y(n_3682)
);

OAI21x1_ASAP7_75t_L g3683 ( 
.A1(n_3556),
.A2(n_2732),
.B(n_2711),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3470),
.Y(n_3684)
);

OAI21x1_ASAP7_75t_L g3685 ( 
.A1(n_3557),
.A2(n_2732),
.B(n_2711),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_3437),
.B(n_2439),
.Y(n_3686)
);

OAI22x1_ASAP7_75t_L g3687 ( 
.A1(n_3551),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_3687)
);

OAI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3453),
.A2(n_3475),
.B(n_3574),
.Y(n_3688)
);

OAI21x1_ASAP7_75t_L g3689 ( 
.A1(n_3560),
.A2(n_72),
.B(n_74),
.Y(n_3689)
);

OAI21x1_ASAP7_75t_L g3690 ( 
.A1(n_3583),
.A2(n_75),
.B(n_76),
.Y(n_3690)
);

OAI21x1_ASAP7_75t_L g3691 ( 
.A1(n_3565),
.A2(n_76),
.B(n_77),
.Y(n_3691)
);

NAND2x1p5_ASAP7_75t_L g3692 ( 
.A(n_3423),
.B(n_675),
.Y(n_3692)
);

AOI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3602),
.A2(n_77),
.B(n_78),
.Y(n_3693)
);

HB1xp67_ASAP7_75t_L g3694 ( 
.A(n_3518),
.Y(n_3694)
);

OAI21x1_ASAP7_75t_L g3695 ( 
.A1(n_3585),
.A2(n_77),
.B(n_79),
.Y(n_3695)
);

AO31x2_ASAP7_75t_L g3696 ( 
.A1(n_3534),
.A2(n_81),
.A3(n_79),
.B(n_80),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3576),
.Y(n_3697)
);

OAI21x1_ASAP7_75t_L g3698 ( 
.A1(n_3587),
.A2(n_80),
.B(n_81),
.Y(n_3698)
);

OAI21x1_ASAP7_75t_L g3699 ( 
.A1(n_3506),
.A2(n_81),
.B(n_82),
.Y(n_3699)
);

OAI21x1_ASAP7_75t_L g3700 ( 
.A1(n_3566),
.A2(n_82),
.B(n_83),
.Y(n_3700)
);

OAI21x1_ASAP7_75t_L g3701 ( 
.A1(n_3579),
.A2(n_82),
.B(n_83),
.Y(n_3701)
);

OAI22x1_ASAP7_75t_L g3702 ( 
.A1(n_3577),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_3702)
);

HB1xp67_ASAP7_75t_L g3703 ( 
.A(n_3518),
.Y(n_3703)
);

BUFx2_ASAP7_75t_L g3704 ( 
.A(n_3434),
.Y(n_3704)
);

OAI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3479),
.A2(n_92),
.B(n_84),
.Y(n_3705)
);

NAND3x1_ASAP7_75t_L g3706 ( 
.A(n_3488),
.B(n_3451),
.C(n_3436),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3428),
.B(n_149),
.Y(n_3707)
);

A2O1A1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3467),
.A2(n_151),
.B(n_152),
.C(n_150),
.Y(n_3708)
);

A2O1A1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3568),
.A2(n_151),
.B(n_153),
.C(n_150),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3533),
.A2(n_85),
.B(n_86),
.Y(n_3710)
);

AOI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_3533),
.A2(n_87),
.B(n_88),
.Y(n_3711)
);

INVx5_ASAP7_75t_L g3712 ( 
.A(n_3571),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3433),
.B(n_153),
.Y(n_3713)
);

O2A1O1Ixp5_ASAP7_75t_SL g3714 ( 
.A1(n_3408),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_3714)
);

AOI21xp5_ASAP7_75t_L g3715 ( 
.A1(n_3494),
.A2(n_87),
.B(n_88),
.Y(n_3715)
);

OR2x2_ASAP7_75t_L g3716 ( 
.A(n_3552),
.B(n_154),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3430),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_SL g3718 ( 
.A1(n_3490),
.A2(n_156),
.B(n_155),
.Y(n_3718)
);

OAI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3589),
.A2(n_89),
.B(n_90),
.Y(n_3719)
);

OAI21x1_ASAP7_75t_L g3720 ( 
.A1(n_3599),
.A2(n_90),
.B(n_91),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3569),
.A2(n_90),
.B(n_92),
.Y(n_3721)
);

OAI21x1_ASAP7_75t_L g3722 ( 
.A1(n_3600),
.A2(n_93),
.B(n_94),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3448),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3446),
.B(n_155),
.Y(n_3724)
);

OAI21x1_ASAP7_75t_L g3725 ( 
.A1(n_3528),
.A2(n_93),
.B(n_94),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3535),
.A2(n_94),
.B(n_95),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3567),
.B(n_157),
.Y(n_3727)
);

CKINVDCx20_ASAP7_75t_R g3728 ( 
.A(n_3459),
.Y(n_3728)
);

AOI211x1_ASAP7_75t_L g3729 ( 
.A1(n_3414),
.A2(n_3432),
.B(n_3404),
.C(n_3495),
.Y(n_3729)
);

OAI21x1_ASAP7_75t_L g3730 ( 
.A1(n_3590),
.A2(n_95),
.B(n_96),
.Y(n_3730)
);

A2O1A1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3503),
.A2(n_158),
.B(n_159),
.C(n_157),
.Y(n_3731)
);

INVx1_ASAP7_75t_SL g3732 ( 
.A(n_3536),
.Y(n_3732)
);

AOI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3602),
.A2(n_95),
.B(n_96),
.Y(n_3733)
);

INVx2_ASAP7_75t_SL g3734 ( 
.A(n_3515),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3590),
.A2(n_96),
.B(n_97),
.Y(n_3735)
);

OAI21x1_ASAP7_75t_L g3736 ( 
.A1(n_3539),
.A2(n_98),
.B(n_99),
.Y(n_3736)
);

NAND3xp33_ASAP7_75t_L g3737 ( 
.A(n_3431),
.B(n_98),
.C(n_99),
.Y(n_3737)
);

BUFx3_ASAP7_75t_L g3738 ( 
.A(n_3466),
.Y(n_3738)
);

AO221x1_ASAP7_75t_L g3739 ( 
.A1(n_3463),
.A2(n_114),
.B1(n_122),
.B2(n_106),
.C(n_98),
.Y(n_3739)
);

OAI21x1_ASAP7_75t_L g3740 ( 
.A1(n_3493),
.A2(n_99),
.B(n_100),
.Y(n_3740)
);

AO31x2_ASAP7_75t_L g3741 ( 
.A1(n_3554),
.A2(n_102),
.A3(n_100),
.B(n_101),
.Y(n_3741)
);

AND2x4_ASAP7_75t_L g3742 ( 
.A(n_3463),
.B(n_100),
.Y(n_3742)
);

AND2x4_ASAP7_75t_L g3743 ( 
.A(n_3545),
.B(n_102),
.Y(n_3743)
);

INVx6_ASAP7_75t_L g3744 ( 
.A(n_3438),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3541),
.A2(n_102),
.B(n_103),
.Y(n_3745)
);

NAND3x1_ASAP7_75t_L g3746 ( 
.A(n_3464),
.B(n_103),
.C(n_104),
.Y(n_3746)
);

INVx4_ASAP7_75t_L g3747 ( 
.A(n_3571),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3465),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3578),
.B(n_158),
.Y(n_3749)
);

AOI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3427),
.A2(n_104),
.B(n_105),
.Y(n_3750)
);

A2O1A1Ixp33_ASAP7_75t_L g3751 ( 
.A1(n_3394),
.A2(n_3481),
.B(n_3549),
.C(n_3462),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3573),
.A2(n_104),
.B(n_105),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_SL g3753 ( 
.A(n_3439),
.B(n_3571),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3468),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3527),
.A2(n_105),
.B(n_106),
.Y(n_3755)
);

INVx2_ASAP7_75t_SL g3756 ( 
.A(n_3455),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3489),
.B(n_686),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_SL g3758 ( 
.A(n_3523),
.B(n_3435),
.Y(n_3758)
);

OAI22xp5_ASAP7_75t_L g3759 ( 
.A1(n_3449),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3759)
);

OAI21x1_ASAP7_75t_L g3760 ( 
.A1(n_3548),
.A2(n_107),
.B(n_108),
.Y(n_3760)
);

BUFx3_ASAP7_75t_L g3761 ( 
.A(n_3592),
.Y(n_3761)
);

AO31x2_ASAP7_75t_L g3762 ( 
.A1(n_3439),
.A2(n_109),
.A3(n_107),
.B(n_108),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3474),
.A2(n_109),
.B(n_110),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3478),
.B(n_3516),
.Y(n_3764)
);

OAI21x1_ASAP7_75t_L g3765 ( 
.A1(n_3526),
.A2(n_110),
.B(n_111),
.Y(n_3765)
);

OAI21x1_ASAP7_75t_SL g3766 ( 
.A1(n_3513),
.A2(n_111),
.B(n_112),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3474),
.A2(n_111),
.B(n_112),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3474),
.A2(n_113),
.B(n_114),
.Y(n_3768)
);

OAI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3484),
.A2(n_113),
.B(n_115),
.Y(n_3769)
);

BUFx6f_ASAP7_75t_L g3770 ( 
.A(n_3562),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3452),
.A2(n_3454),
.B(n_3491),
.Y(n_3771)
);

AOI21x1_ASAP7_75t_SL g3772 ( 
.A1(n_3500),
.A2(n_164),
.B(n_159),
.Y(n_3772)
);

OAI21x1_ASAP7_75t_L g3773 ( 
.A1(n_3532),
.A2(n_115),
.B(n_116),
.Y(n_3773)
);

OAI21x1_ASAP7_75t_SL g3774 ( 
.A1(n_3520),
.A2(n_115),
.B(n_116),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3512),
.A2(n_116),
.B(n_117),
.Y(n_3775)
);

CKINVDCx5p33_ASAP7_75t_R g3776 ( 
.A(n_3546),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3496),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3502),
.B(n_164),
.Y(n_3778)
);

INVxp67_ASAP7_75t_L g3779 ( 
.A(n_3584),
.Y(n_3779)
);

NOR2x1_ASAP7_75t_SL g3780 ( 
.A(n_3438),
.B(n_165),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3507),
.B(n_165),
.Y(n_3781)
);

OAI21x1_ASAP7_75t_L g3782 ( 
.A1(n_3395),
.A2(n_3538),
.B(n_3424),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3514),
.Y(n_3783)
);

BUFx6f_ASAP7_75t_L g3784 ( 
.A(n_3562),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3555),
.B(n_693),
.Y(n_3785)
);

OAI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3395),
.A2(n_117),
.B(n_118),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3525),
.B(n_166),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3486),
.B(n_166),
.Y(n_3788)
);

OAI21x1_ASAP7_75t_L g3789 ( 
.A1(n_3510),
.A2(n_117),
.B(n_118),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3540),
.B(n_167),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3519),
.B(n_169),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3596),
.A2(n_118),
.B(n_119),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3469),
.A2(n_119),
.B(n_120),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3521),
.B(n_169),
.Y(n_3794)
);

OAI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3410),
.A2(n_119),
.B(n_120),
.Y(n_3795)
);

OAI21x1_ASAP7_75t_L g3796 ( 
.A1(n_3603),
.A2(n_121),
.B(n_122),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3606),
.A2(n_121),
.B(n_122),
.Y(n_3797)
);

AO22x2_ASAP7_75t_L g3798 ( 
.A1(n_3501),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3487),
.B(n_170),
.Y(n_3799)
);

NAND2xp33_ASAP7_75t_L g3800 ( 
.A(n_3410),
.B(n_172),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3586),
.B(n_173),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_SL g3802 ( 
.A1(n_3575),
.A2(n_173),
.B(n_174),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3537),
.B(n_174),
.Y(n_3803)
);

OAI21x1_ASAP7_75t_L g3804 ( 
.A1(n_3480),
.A2(n_175),
.B(n_176),
.Y(n_3804)
);

NAND2x1p5_ASAP7_75t_L g3805 ( 
.A(n_3504),
.B(n_177),
.Y(n_3805)
);

OAI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_3480),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3595),
.A2(n_178),
.B(n_179),
.Y(n_3807)
);

NAND3xp33_ASAP7_75t_SL g3808 ( 
.A(n_3530),
.B(n_180),
.C(n_181),
.Y(n_3808)
);

AOI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3410),
.A2(n_183),
.B1(n_180),
.B2(n_182),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3593),
.Y(n_3810)
);

OAI21x1_ASAP7_75t_L g3811 ( 
.A1(n_3597),
.A2(n_182),
.B(n_183),
.Y(n_3811)
);

OAI21x1_ASAP7_75t_L g3812 ( 
.A1(n_3598),
.A2(n_184),
.B(n_185),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3570),
.A2(n_186),
.B(n_188),
.Y(n_3813)
);

BUFx4_ASAP7_75t_SL g3814 ( 
.A(n_3601),
.Y(n_3814)
);

INVx1_ASAP7_75t_SL g3815 ( 
.A(n_3605),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3410),
.B(n_186),
.Y(n_3816)
);

NAND3xp33_ASAP7_75t_L g3817 ( 
.A(n_3591),
.B(n_188),
.C(n_189),
.Y(n_3817)
);

AOI211x1_ASAP7_75t_L g3818 ( 
.A1(n_3559),
.A2(n_194),
.B(n_190),
.C(n_192),
.Y(n_3818)
);

OAI21x1_ASAP7_75t_L g3819 ( 
.A1(n_3570),
.A2(n_192),
.B(n_194),
.Y(n_3819)
);

CKINVDCx20_ASAP7_75t_R g3820 ( 
.A(n_3407),
.Y(n_3820)
);

AOI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_3522),
.A2(n_198),
.B1(n_195),
.B2(n_196),
.Y(n_3821)
);

AND2x4_ASAP7_75t_L g3822 ( 
.A(n_3561),
.B(n_195),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3572),
.A2(n_196),
.B(n_198),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3562),
.Y(n_3824)
);

BUFx2_ASAP7_75t_L g3825 ( 
.A(n_3561),
.Y(n_3825)
);

OAI21xp33_ASAP7_75t_L g3826 ( 
.A1(n_3529),
.A2(n_199),
.B(n_200),
.Y(n_3826)
);

NOR2xp67_ASAP7_75t_L g3827 ( 
.A(n_3604),
.B(n_199),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3438),
.B(n_691),
.Y(n_3828)
);

OAI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3460),
.A2(n_200),
.B(n_201),
.Y(n_3829)
);

BUFx2_ASAP7_75t_SL g3830 ( 
.A(n_3460),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3460),
.A2(n_201),
.B(n_202),
.Y(n_3831)
);

AND2x6_ASAP7_75t_SL g3832 ( 
.A(n_3394),
.B(n_202),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3497),
.B(n_203),
.Y(n_3833)
);

OAI21x1_ASAP7_75t_L g3834 ( 
.A1(n_3508),
.A2(n_204),
.B(n_205),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3543),
.Y(n_3835)
);

BUFx2_ASAP7_75t_L g3836 ( 
.A(n_3651),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3697),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3783),
.B(n_205),
.Y(n_3838)
);

AOI21xp5_ASAP7_75t_L g3839 ( 
.A1(n_3800),
.A2(n_206),
.B(n_207),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3732),
.B(n_207),
.Y(n_3840)
);

INVx4_ASAP7_75t_L g3841 ( 
.A(n_3776),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3662),
.A2(n_209),
.B(n_210),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3631),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3648),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3835),
.Y(n_3845)
);

AO31x2_ASAP7_75t_L g3846 ( 
.A1(n_3657),
.A2(n_211),
.A3(n_209),
.B(n_210),
.Y(n_3846)
);

OAI21xp33_ASAP7_75t_L g3847 ( 
.A1(n_3718),
.A2(n_211),
.B(n_212),
.Y(n_3847)
);

OR2x2_ASAP7_75t_L g3848 ( 
.A(n_3639),
.B(n_212),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3672),
.Y(n_3849)
);

AOI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3662),
.A2(n_213),
.B(n_214),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3680),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3684),
.Y(n_3852)
);

OAI21xp5_ASAP7_75t_L g3853 ( 
.A1(n_3715),
.A2(n_3705),
.B(n_3726),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3612),
.A2(n_213),
.B(n_214),
.Y(n_3854)
);

INVx2_ASAP7_75t_SL g3855 ( 
.A(n_3738),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3694),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3717),
.Y(n_3857)
);

CKINVDCx11_ASAP7_75t_R g3858 ( 
.A(n_3728),
.Y(n_3858)
);

OR2x6_ASAP7_75t_L g3859 ( 
.A(n_3627),
.B(n_215),
.Y(n_3859)
);

AOI22xp5_ASAP7_75t_L g3860 ( 
.A1(n_3809),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_3860)
);

A2O1A1Ixp33_ASAP7_75t_L g3861 ( 
.A1(n_3826),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_3861)
);

OAI21x1_ASAP7_75t_L g3862 ( 
.A1(n_3620),
.A2(n_218),
.B(n_219),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3610),
.A2(n_3667),
.B(n_3624),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3764),
.B(n_220),
.Y(n_3864)
);

AO31x2_ASAP7_75t_L g3865 ( 
.A1(n_3708),
.A2(n_222),
.A3(n_220),
.B(n_221),
.Y(n_3865)
);

NAND2x1p5_ASAP7_75t_L g3866 ( 
.A(n_3712),
.B(n_221),
.Y(n_3866)
);

OAI21x1_ASAP7_75t_L g3867 ( 
.A1(n_3671),
.A2(n_222),
.B(n_223),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3610),
.A2(n_223),
.B(n_224),
.Y(n_3868)
);

AOI21xp5_ASAP7_75t_L g3869 ( 
.A1(n_3667),
.A2(n_224),
.B(n_226),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3688),
.A2(n_227),
.B(n_228),
.Y(n_3870)
);

OAI21x1_ASAP7_75t_L g3871 ( 
.A1(n_3682),
.A2(n_227),
.B(n_228),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3771),
.B(n_229),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3688),
.A2(n_3632),
.B(n_3705),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3732),
.B(n_229),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3611),
.B(n_3609),
.Y(n_3875)
);

INVx4_ASAP7_75t_L g3876 ( 
.A(n_3618),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3653),
.A2(n_230),
.B(n_231),
.Y(n_3877)
);

OAI21x1_ASAP7_75t_L g3878 ( 
.A1(n_3655),
.A2(n_230),
.B(n_231),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3810),
.Y(n_3879)
);

INVx5_ASAP7_75t_L g3880 ( 
.A(n_3617),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3625),
.A2(n_232),
.B(n_233),
.Y(n_3881)
);

BUFx6f_ASAP7_75t_L g3882 ( 
.A(n_3770),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3723),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3643),
.B(n_232),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3613),
.A2(n_233),
.B(n_234),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3637),
.A2(n_235),
.B(n_236),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3681),
.A2(n_3795),
.B(n_3686),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3748),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3795),
.A2(n_235),
.B(n_237),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_3814),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3630),
.A2(n_237),
.B(n_238),
.Y(n_3891)
);

A2O1A1Ixp33_ASAP7_75t_L g3892 ( 
.A1(n_3826),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3751),
.A2(n_240),
.B(n_242),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3652),
.A2(n_243),
.B(n_244),
.Y(n_3894)
);

AO31x2_ASAP7_75t_L g3895 ( 
.A1(n_3710),
.A2(n_245),
.A3(n_243),
.B(n_244),
.Y(n_3895)
);

AO31x2_ASAP7_75t_L g3896 ( 
.A1(n_3711),
.A2(n_247),
.A3(n_245),
.B(n_246),
.Y(n_3896)
);

OAI21x1_ASAP7_75t_L g3897 ( 
.A1(n_3649),
.A2(n_247),
.B(n_248),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3621),
.B(n_249),
.Y(n_3898)
);

AO31x2_ASAP7_75t_L g3899 ( 
.A1(n_3709),
.A2(n_253),
.A3(n_251),
.B(n_252),
.Y(n_3899)
);

AO31x2_ASAP7_75t_L g3900 ( 
.A1(n_3731),
.A2(n_254),
.A3(n_252),
.B(n_253),
.Y(n_3900)
);

BUFx2_ASAP7_75t_SL g3901 ( 
.A(n_3820),
.Y(n_3901)
);

O2A1O1Ixp33_ASAP7_75t_SL g3902 ( 
.A1(n_3758),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_3902)
);

OAI21x1_ASAP7_75t_L g3903 ( 
.A1(n_3644),
.A2(n_255),
.B(n_257),
.Y(n_3903)
);

AOI21x1_ASAP7_75t_L g3904 ( 
.A1(n_3799),
.A2(n_258),
.B(n_259),
.Y(n_3904)
);

AO31x2_ASAP7_75t_L g3905 ( 
.A1(n_3687),
.A2(n_260),
.A3(n_258),
.B(n_259),
.Y(n_3905)
);

NOR2xp67_ASAP7_75t_SL g3906 ( 
.A(n_3737),
.B(n_260),
.Y(n_3906)
);

O2A1O1Ixp33_ASAP7_75t_SL g3907 ( 
.A1(n_3829),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_3907)
);

OAI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3809),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3642),
.B(n_264),
.Y(n_3909)
);

AND2x4_ASAP7_75t_L g3910 ( 
.A(n_3658),
.B(n_3825),
.Y(n_3910)
);

OAI21x1_ASAP7_75t_L g3911 ( 
.A1(n_3699),
.A2(n_265),
.B(n_266),
.Y(n_3911)
);

BUFx10_ASAP7_75t_L g3912 ( 
.A(n_3742),
.Y(n_3912)
);

OAI21x1_ASAP7_75t_L g3913 ( 
.A1(n_3683),
.A2(n_265),
.B(n_266),
.Y(n_3913)
);

BUFx6f_ASAP7_75t_L g3914 ( 
.A(n_3770),
.Y(n_3914)
);

OA22x2_ASAP7_75t_L g3915 ( 
.A1(n_3739),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_3915)
);

O2A1O1Ixp33_ASAP7_75t_SL g3916 ( 
.A1(n_3829),
.A2(n_3759),
.B(n_3816),
.C(n_3737),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3652),
.A2(n_3638),
.B(n_3669),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3659),
.A2(n_267),
.B(n_268),
.Y(n_3918)
);

AO31x2_ASAP7_75t_L g3919 ( 
.A1(n_3702),
.A2(n_272),
.A3(n_270),
.B(n_271),
.Y(n_3919)
);

OAI21x1_ASAP7_75t_L g3920 ( 
.A1(n_3685),
.A2(n_271),
.B(n_272),
.Y(n_3920)
);

OAI22x1_ASAP7_75t_L g3921 ( 
.A1(n_3704),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3754),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_L g3923 ( 
.A(n_3614),
.B(n_274),
.Y(n_3923)
);

O2A1O1Ixp5_ASAP7_75t_SL g3924 ( 
.A1(n_3635),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_3924)
);

AND2x4_ASAP7_75t_L g3925 ( 
.A(n_3747),
.B(n_276),
.Y(n_3925)
);

OAI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3665),
.A2(n_277),
.B(n_278),
.Y(n_3926)
);

INVx4_ASAP7_75t_L g3927 ( 
.A(n_3770),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3817),
.A2(n_278),
.B(n_279),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3817),
.A2(n_279),
.B(n_280),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3777),
.B(n_280),
.Y(n_3930)
);

BUFx6f_ASAP7_75t_L g3931 ( 
.A(n_3784),
.Y(n_3931)
);

OAI21xp5_ASAP7_75t_L g3932 ( 
.A1(n_3746),
.A2(n_281),
.B(n_282),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3608),
.B(n_281),
.Y(n_3933)
);

CKINVDCx20_ASAP7_75t_R g3934 ( 
.A(n_3761),
.Y(n_3934)
);

NOR2xp33_ASAP7_75t_L g3935 ( 
.A(n_3779),
.B(n_282),
.Y(n_3935)
);

O2A1O1Ixp33_ASAP7_75t_SL g3936 ( 
.A1(n_3788),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_3936)
);

AO31x2_ASAP7_75t_L g3937 ( 
.A1(n_3752),
.A2(n_3674),
.A3(n_3793),
.B(n_3663),
.Y(n_3937)
);

AO31x2_ASAP7_75t_L g3938 ( 
.A1(n_3747),
.A2(n_285),
.A3(n_283),
.B(n_284),
.Y(n_3938)
);

AO22x1_ASAP7_75t_L g3939 ( 
.A1(n_3712),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3753),
.A2(n_289),
.B(n_290),
.Y(n_3940)
);

BUFx2_ASAP7_75t_L g3941 ( 
.A(n_3703),
.Y(n_3941)
);

AOI31xp67_ASAP7_75t_L g3942 ( 
.A1(n_3821),
.A2(n_292),
.A3(n_290),
.B(n_291),
.Y(n_3942)
);

OAI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_3750),
.A2(n_292),
.B(n_293),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3616),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3607),
.Y(n_3945)
);

XNOR2xp5_ASAP7_75t_L g3946 ( 
.A(n_3706),
.B(n_294),
.Y(n_3946)
);

O2A1O1Ixp5_ASAP7_75t_L g3947 ( 
.A1(n_3763),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_3947)
);

AOI221x1_ASAP7_75t_L g3948 ( 
.A1(n_3664),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_298),
.Y(n_3948)
);

AO32x2_ASAP7_75t_L g3949 ( 
.A1(n_3756),
.A2(n_299),
.A3(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_3949)
);

OAI21x1_ASAP7_75t_L g3950 ( 
.A1(n_3740),
.A2(n_299),
.B(n_300),
.Y(n_3950)
);

OAI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3698),
.A2(n_301),
.B(n_302),
.Y(n_3951)
);

CKINVDCx5p33_ASAP7_75t_R g3952 ( 
.A(n_3734),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_SL g3953 ( 
.A(n_3729),
.B(n_3615),
.Y(n_3953)
);

A2O1A1Ixp33_ASAP7_75t_L g3954 ( 
.A1(n_3823),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_3954)
);

OAI22x1_ASAP7_75t_L g3955 ( 
.A1(n_3821),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3753),
.A2(n_304),
.B(n_306),
.Y(n_3956)
);

AOI221xp5_ASAP7_75t_SL g3957 ( 
.A1(n_3831),
.A2(n_3755),
.B1(n_3767),
.B2(n_3768),
.C(n_3775),
.Y(n_3957)
);

OAI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3645),
.A2(n_310),
.B1(n_306),
.B2(n_307),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3707),
.A2(n_307),
.B(n_312),
.Y(n_3959)
);

INVxp67_ASAP7_75t_SL g3960 ( 
.A(n_3607),
.Y(n_3960)
);

AOI221xp5_ASAP7_75t_SL g3961 ( 
.A1(n_3806),
.A2(n_3721),
.B1(n_3646),
.B2(n_3749),
.C(n_3727),
.Y(n_3961)
);

A2O1A1Ixp33_ASAP7_75t_L g3962 ( 
.A1(n_3736),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_3962)
);

BUFx10_ASAP7_75t_L g3963 ( 
.A(n_3742),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3629),
.B(n_313),
.Y(n_3964)
);

OAI21xp33_ASAP7_75t_L g3965 ( 
.A1(n_3664),
.A2(n_315),
.B(n_316),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3622),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3636),
.B(n_316),
.Y(n_3967)
);

BUFx10_ASAP7_75t_L g3968 ( 
.A(n_3803),
.Y(n_3968)
);

AO32x2_ASAP7_75t_L g3969 ( 
.A1(n_3656),
.A2(n_319),
.A3(n_317),
.B1(n_318),
.B2(n_320),
.Y(n_3969)
);

OAI21x1_ASAP7_75t_L g3970 ( 
.A1(n_3650),
.A2(n_318),
.B(n_319),
.Y(n_3970)
);

OAI21x1_ASAP7_75t_L g3971 ( 
.A1(n_3695),
.A2(n_321),
.B(n_322),
.Y(n_3971)
);

INVx2_ASAP7_75t_SL g3972 ( 
.A(n_3784),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_L g3973 ( 
.A(n_3832),
.B(n_321),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3622),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3622),
.Y(n_3975)
);

A2O1A1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3808),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3824),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3640),
.Y(n_3978)
);

OAI21x1_ASAP7_75t_L g3979 ( 
.A1(n_3834),
.A2(n_323),
.B(n_324),
.Y(n_3979)
);

AOI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3666),
.A2(n_3661),
.B(n_3628),
.Y(n_3980)
);

OAI21x1_ASAP7_75t_L g3981 ( 
.A1(n_3619),
.A2(n_326),
.B(n_327),
.Y(n_3981)
);

AO31x2_ASAP7_75t_L g3982 ( 
.A1(n_3696),
.A2(n_329),
.A3(n_326),
.B(n_328),
.Y(n_3982)
);

NOR2xp33_ASAP7_75t_L g3983 ( 
.A(n_3832),
.B(n_328),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3647),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3641),
.A2(n_330),
.B(n_331),
.Y(n_3985)
);

AO32x2_ASAP7_75t_L g3986 ( 
.A1(n_3656),
.A2(n_334),
.A3(n_332),
.B1(n_333),
.B2(n_335),
.Y(n_3986)
);

AO31x2_ASAP7_75t_L g3987 ( 
.A1(n_3696),
.A2(n_336),
.A3(n_332),
.B(n_335),
.Y(n_3987)
);

CKINVDCx6p67_ASAP7_75t_R g3988 ( 
.A(n_3830),
.Y(n_3988)
);

INVxp67_ASAP7_75t_L g3989 ( 
.A(n_3654),
.Y(n_3989)
);

OAI21x1_ASAP7_75t_L g3990 ( 
.A1(n_3689),
.A2(n_337),
.B(n_338),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3626),
.A2(n_338),
.B(n_339),
.Y(n_3991)
);

OAI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_3719),
.A2(n_339),
.B(n_340),
.Y(n_3992)
);

NOR2x1_ASAP7_75t_L g3993 ( 
.A(n_3647),
.B(n_3675),
.Y(n_3993)
);

OAI21x1_ASAP7_75t_L g3994 ( 
.A1(n_3730),
.A2(n_341),
.B(n_342),
.Y(n_3994)
);

INVx5_ASAP7_75t_L g3995 ( 
.A(n_3712),
.Y(n_3995)
);

A2O1A1Ixp33_ASAP7_75t_L g3996 ( 
.A1(n_3789),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_3996)
);

O2A1O1Ixp5_ASAP7_75t_SL g3997 ( 
.A1(n_3675),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_3997)
);

BUFx10_ASAP7_75t_L g3998 ( 
.A(n_3790),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3640),
.Y(n_3999)
);

AO31x2_ASAP7_75t_L g4000 ( 
.A1(n_3696),
.A2(n_346),
.A3(n_344),
.B(n_345),
.Y(n_4000)
);

INVxp67_ASAP7_75t_L g4001 ( 
.A(n_3660),
.Y(n_4001)
);

AOI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_3700),
.A2(n_346),
.B(n_347),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3716),
.B(n_347),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3782),
.A2(n_348),
.B(n_349),
.Y(n_4004)
);

OAI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_3645),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3691),
.A2(n_352),
.B(n_353),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3640),
.B(n_352),
.Y(n_4007)
);

OAI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3701),
.A2(n_355),
.B(n_356),
.Y(n_4008)
);

OAI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3690),
.A2(n_355),
.B(n_356),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3729),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_4010)
);

OR2x2_ASAP7_75t_L g4011 ( 
.A(n_3741),
.B(n_357),
.Y(n_4011)
);

CKINVDCx8_ASAP7_75t_R g4012 ( 
.A(n_3784),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3678),
.Y(n_4013)
);

CKINVDCx16_ASAP7_75t_R g4014 ( 
.A(n_3676),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3735),
.A2(n_360),
.B(n_361),
.Y(n_4015)
);

OAI21x1_ASAP7_75t_L g4016 ( 
.A1(n_3720),
.A2(n_360),
.B(n_361),
.Y(n_4016)
);

BUFx2_ASAP7_75t_L g4017 ( 
.A(n_3678),
.Y(n_4017)
);

INVx1_ASAP7_75t_SL g4018 ( 
.A(n_4017),
.Y(n_4018)
);

INVx6_ASAP7_75t_L g4019 ( 
.A(n_3880),
.Y(n_4019)
);

NAND2x1p5_ASAP7_75t_L g4020 ( 
.A(n_3995),
.B(n_3633),
.Y(n_4020)
);

HB1xp67_ASAP7_75t_L g4021 ( 
.A(n_3836),
.Y(n_4021)
);

INVxp67_ASAP7_75t_L g4022 ( 
.A(n_3836),
.Y(n_4022)
);

OAI21x1_ASAP7_75t_SL g4023 ( 
.A1(n_3873),
.A2(n_3780),
.B(n_3733),
.Y(n_4023)
);

OAI33xp33_ASAP7_75t_L g4024 ( 
.A1(n_3908),
.A2(n_3833),
.A3(n_3724),
.B1(n_3787),
.B2(n_3794),
.B3(n_3791),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3977),
.Y(n_4025)
);

OR2x2_ASAP7_75t_L g4026 ( 
.A(n_3879),
.B(n_3741),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3853),
.A2(n_3802),
.B1(n_3798),
.B2(n_3743),
.Y(n_4027)
);

AO31x2_ASAP7_75t_L g4028 ( 
.A1(n_3948),
.A2(n_3656),
.A3(n_3781),
.B(n_3778),
.Y(n_4028)
);

NOR2xp67_ASAP7_75t_L g4029 ( 
.A(n_3995),
.B(n_3679),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3837),
.Y(n_4030)
);

AND2x4_ASAP7_75t_L g4031 ( 
.A(n_3993),
.B(n_3679),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3849),
.Y(n_4032)
);

BUFx2_ASAP7_75t_SL g4033 ( 
.A(n_3934),
.Y(n_4033)
);

OAI21x1_ASAP7_75t_L g4034 ( 
.A1(n_3863),
.A2(n_3786),
.B(n_3693),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3875),
.B(n_3741),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3910),
.B(n_4014),
.Y(n_4036)
);

OAI21x1_ASAP7_75t_L g4037 ( 
.A1(n_3974),
.A2(n_3722),
.B(n_3725),
.Y(n_4037)
);

NAND2x1p5_ASAP7_75t_L g4038 ( 
.A(n_3995),
.B(n_3815),
.Y(n_4038)
);

INVx2_ASAP7_75t_SL g4039 ( 
.A(n_3952),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_4017),
.Y(n_4040)
);

OA21x2_ASAP7_75t_L g4041 ( 
.A1(n_3945),
.A2(n_3615),
.B(n_3634),
.Y(n_4041)
);

AO31x2_ASAP7_75t_L g4042 ( 
.A1(n_3975),
.A2(n_3713),
.A3(n_3668),
.B(n_3670),
.Y(n_4042)
);

OAI21x1_ASAP7_75t_L g4043 ( 
.A1(n_3966),
.A2(n_3745),
.B(n_3765),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_L g4044 ( 
.A(n_3876),
.B(n_3673),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3852),
.Y(n_4045)
);

OA21x2_ASAP7_75t_L g4046 ( 
.A1(n_3960),
.A2(n_3634),
.B(n_3773),
.Y(n_4046)
);

NAND2xp33_ASAP7_75t_SL g4047 ( 
.A(n_3946),
.B(n_3743),
.Y(n_4047)
);

OAI21x1_ASAP7_75t_L g4048 ( 
.A1(n_3862),
.A2(n_3772),
.B(n_3769),
.Y(n_4048)
);

AOI21x1_ASAP7_75t_L g4049 ( 
.A1(n_3872),
.A2(n_3827),
.B(n_3798),
.Y(n_4049)
);

OAI21x1_ASAP7_75t_L g4050 ( 
.A1(n_3978),
.A2(n_3760),
.B(n_3792),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3843),
.B(n_3623),
.Y(n_4051)
);

BUFx6f_ASAP7_75t_L g4052 ( 
.A(n_3858),
.Y(n_4052)
);

AND2x4_ASAP7_75t_L g4053 ( 
.A(n_3941),
.B(n_3815),
.Y(n_4053)
);

OAI221xp5_ASAP7_75t_L g4054 ( 
.A1(n_3893),
.A2(n_3692),
.B1(n_3827),
.B2(n_3805),
.C(n_3801),
.Y(n_4054)
);

NAND3xp33_ASAP7_75t_L g4055 ( 
.A(n_3870),
.B(n_3818),
.C(n_3714),
.Y(n_4055)
);

OAI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3999),
.A2(n_3797),
.B(n_3796),
.Y(n_4056)
);

CKINVDCx5p33_ASAP7_75t_R g4057 ( 
.A(n_3890),
.Y(n_4057)
);

AO21x2_ASAP7_75t_L g4058 ( 
.A1(n_3944),
.A2(n_4004),
.B(n_3868),
.Y(n_4058)
);

OAI22xp33_ASAP7_75t_SL g4059 ( 
.A1(n_3973),
.A2(n_3822),
.B1(n_3744),
.B2(n_3818),
.Y(n_4059)
);

OAI21x1_ASAP7_75t_L g4060 ( 
.A1(n_3917),
.A2(n_3819),
.B(n_3813),
.Y(n_4060)
);

O2A1O1Ixp33_ASAP7_75t_L g4061 ( 
.A1(n_3861),
.A2(n_3766),
.B(n_3774),
.C(n_3822),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3844),
.B(n_3623),
.Y(n_4062)
);

OAI21x1_ASAP7_75t_L g4063 ( 
.A1(n_3897),
.A2(n_3804),
.B(n_3807),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3845),
.Y(n_4064)
);

INVx1_ASAP7_75t_SL g4065 ( 
.A(n_3941),
.Y(n_4065)
);

OR2x6_ASAP7_75t_L g4066 ( 
.A(n_3887),
.B(n_3677),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3922),
.Y(n_4067)
);

INVx3_ASAP7_75t_L g4068 ( 
.A(n_3984),
.Y(n_4068)
);

AOI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_3847),
.A2(n_3785),
.B1(n_3757),
.B2(n_3828),
.Y(n_4069)
);

NAND2xp33_ASAP7_75t_L g4070 ( 
.A(n_3946),
.B(n_3762),
.Y(n_4070)
);

OA21x2_ASAP7_75t_L g4071 ( 
.A1(n_3953),
.A2(n_3980),
.B(n_3903),
.Y(n_4071)
);

OAI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_3894),
.A2(n_3812),
.B(n_3811),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3851),
.Y(n_4073)
);

OAI21x1_ASAP7_75t_L g4074 ( 
.A1(n_3878),
.A2(n_3623),
.B(n_3762),
.Y(n_4074)
);

OA21x2_ASAP7_75t_L g4075 ( 
.A1(n_3981),
.A2(n_3762),
.B(n_3744),
.Y(n_4075)
);

OAI21x1_ASAP7_75t_SL g4076 ( 
.A1(n_3932),
.A2(n_362),
.B(n_363),
.Y(n_4076)
);

O2A1O1Ixp33_ASAP7_75t_SL g4077 ( 
.A1(n_3983),
.A2(n_690),
.B(n_364),
.C(n_362),
.Y(n_4077)
);

BUFx6f_ASAP7_75t_L g4078 ( 
.A(n_3882),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3857),
.Y(n_4079)
);

NOR2xp33_ASAP7_75t_L g4080 ( 
.A(n_3841),
.B(n_363),
.Y(n_4080)
);

OA21x2_ASAP7_75t_L g4081 ( 
.A1(n_3856),
.A2(n_364),
.B(n_365),
.Y(n_4081)
);

OAI21x1_ASAP7_75t_L g4082 ( 
.A1(n_3970),
.A2(n_365),
.B(n_366),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_3928),
.A2(n_690),
.B(n_366),
.Y(n_4083)
);

OAI21x1_ASAP7_75t_L g4084 ( 
.A1(n_3871),
.A2(n_3920),
.B(n_3913),
.Y(n_4084)
);

OA21x2_ASAP7_75t_L g4085 ( 
.A1(n_3867),
.A2(n_367),
.B(n_368),
.Y(n_4085)
);

O2A1O1Ixp33_ASAP7_75t_SL g4086 ( 
.A1(n_3840),
.A2(n_370),
.B(n_367),
.C(n_369),
.Y(n_4086)
);

NAND3x1_ASAP7_75t_L g4087 ( 
.A(n_3923),
.B(n_370),
.C(n_371),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3883),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3888),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_4013),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3989),
.Y(n_4091)
);

A2O1A1Ixp33_ASAP7_75t_L g4092 ( 
.A1(n_3965),
.A2(n_689),
.B(n_373),
.C(n_371),
.Y(n_4092)
);

BUFx3_ASAP7_75t_L g4093 ( 
.A(n_3855),
.Y(n_4093)
);

CKINVDCx12_ASAP7_75t_R g4094 ( 
.A(n_3859),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4001),
.B(n_372),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4007),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3901),
.B(n_372),
.Y(n_4097)
);

OAI21x1_ASAP7_75t_L g4098 ( 
.A1(n_3911),
.A2(n_373),
.B(n_374),
.Y(n_4098)
);

OAI21x1_ASAP7_75t_L g4099 ( 
.A1(n_3950),
.A2(n_374),
.B(n_375),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4011),
.Y(n_4100)
);

AOI22xp33_ASAP7_75t_L g4101 ( 
.A1(n_3926),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4101)
);

OA21x2_ASAP7_75t_L g4102 ( 
.A1(n_3842),
.A2(n_376),
.B(n_377),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3912),
.B(n_379),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3909),
.B(n_379),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3898),
.B(n_380),
.Y(n_4105)
);

INVx3_ASAP7_75t_L g4106 ( 
.A(n_3927),
.Y(n_4106)
);

AND2x4_ASAP7_75t_L g4107 ( 
.A(n_3972),
.B(n_381),
.Y(n_4107)
);

AOI21xp33_ASAP7_75t_L g4108 ( 
.A1(n_3906),
.A2(n_382),
.B(n_383),
.Y(n_4108)
);

OAI21x1_ASAP7_75t_L g4109 ( 
.A1(n_3979),
.A2(n_382),
.B(n_384),
.Y(n_4109)
);

AND2x4_ASAP7_75t_L g4110 ( 
.A(n_3880),
.B(n_385),
.Y(n_4110)
);

BUFx2_ASAP7_75t_L g4111 ( 
.A(n_3882),
.Y(n_4111)
);

BUFx3_ASAP7_75t_L g4112 ( 
.A(n_3880),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3864),
.B(n_385),
.Y(n_4113)
);

OR2x2_ASAP7_75t_L g4114 ( 
.A(n_3848),
.B(n_689),
.Y(n_4114)
);

NOR2x1_ASAP7_75t_SL g4115 ( 
.A(n_3859),
.B(n_386),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3930),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3982),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_3963),
.B(n_388),
.Y(n_4118)
);

OA21x2_ASAP7_75t_L g4119 ( 
.A1(n_3850),
.A2(n_388),
.B(n_389),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3964),
.B(n_390),
.Y(n_4120)
);

BUFx6f_ASAP7_75t_L g4121 ( 
.A(n_3914),
.Y(n_4121)
);

NAND3xp33_ASAP7_75t_L g4122 ( 
.A(n_3929),
.B(n_391),
.C(n_392),
.Y(n_4122)
);

OAI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3860),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3982),
.B(n_393),
.Y(n_4124)
);

OAI21x1_ASAP7_75t_L g4125 ( 
.A1(n_3990),
.A2(n_394),
.B(n_396),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3987),
.Y(n_4126)
);

BUFx3_ASAP7_75t_L g4127 ( 
.A(n_3988),
.Y(n_4127)
);

INVx3_ASAP7_75t_L g4128 ( 
.A(n_4012),
.Y(n_4128)
);

NAND2x1p5_ASAP7_75t_L g4129 ( 
.A(n_3914),
.B(n_394),
.Y(n_4129)
);

OAI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3889),
.A2(n_397),
.B(n_398),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3987),
.B(n_398),
.Y(n_4131)
);

OAI21x1_ASAP7_75t_L g4132 ( 
.A1(n_3985),
.A2(n_399),
.B(n_400),
.Y(n_4132)
);

OAI21xp5_ASAP7_75t_L g4133 ( 
.A1(n_3869),
.A2(n_400),
.B(n_401),
.Y(n_4133)
);

OAI21x1_ASAP7_75t_SL g4134 ( 
.A1(n_3886),
.A2(n_401),
.B(n_402),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4000),
.B(n_402),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_3958),
.A2(n_406),
.B1(n_403),
.B2(n_405),
.Y(n_4136)
);

HB1xp67_ASAP7_75t_L g4137 ( 
.A(n_4000),
.Y(n_4137)
);

INVx2_ASAP7_75t_SL g4138 ( 
.A(n_3931),
.Y(n_4138)
);

INVx3_ASAP7_75t_L g4139 ( 
.A(n_3931),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_L g4140 ( 
.A1(n_4005),
.A2(n_408),
.B1(n_403),
.B2(n_406),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3838),
.Y(n_4141)
);

OAI21xp33_ASAP7_75t_SL g4142 ( 
.A1(n_3915),
.A2(n_409),
.B(n_410),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3904),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3967),
.B(n_409),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3884),
.B(n_411),
.Y(n_4145)
);

OAI21x1_ASAP7_75t_L g4146 ( 
.A1(n_4002),
.A2(n_411),
.B(n_412),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_3943),
.A2(n_3839),
.B1(n_3854),
.B2(n_4010),
.Y(n_4147)
);

OAI21x1_ASAP7_75t_L g4148 ( 
.A1(n_4006),
.A2(n_412),
.B(n_413),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3846),
.Y(n_4149)
);

INVx3_ASAP7_75t_L g4150 ( 
.A(n_3998),
.Y(n_4150)
);

OAI21x1_ASAP7_75t_L g4151 ( 
.A1(n_3971),
.A2(n_413),
.B(n_414),
.Y(n_4151)
);

OA21x2_ASAP7_75t_L g4152 ( 
.A1(n_4008),
.A2(n_3951),
.B(n_3992),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3846),
.Y(n_4153)
);

BUFx3_ASAP7_75t_L g4154 ( 
.A(n_3968),
.Y(n_4154)
);

INVx2_ASAP7_75t_SL g4155 ( 
.A(n_3925),
.Y(n_4155)
);

BUFx3_ASAP7_75t_L g4156 ( 
.A(n_3933),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3969),
.Y(n_4157)
);

NAND3xp33_ASAP7_75t_L g4158 ( 
.A(n_3891),
.B(n_414),
.C(n_415),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3969),
.Y(n_4159)
);

NAND2x1_ASAP7_75t_L g4160 ( 
.A(n_3940),
.B(n_416),
.Y(n_4160)
);

A2O1A1Ixp33_ASAP7_75t_L g4161 ( 
.A1(n_3956),
.A2(n_419),
.B(n_416),
.C(n_418),
.Y(n_4161)
);

A2O1A1Ixp33_ASAP7_75t_L g4162 ( 
.A1(n_3892),
.A2(n_685),
.B(n_420),
.C(n_418),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3986),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3986),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3938),
.Y(n_4165)
);

OA21x2_ASAP7_75t_L g4166 ( 
.A1(n_4009),
.A2(n_419),
.B(n_420),
.Y(n_4166)
);

CKINVDCx5p33_ASAP7_75t_R g4167 ( 
.A(n_3935),
.Y(n_4167)
);

OA21x2_ASAP7_75t_L g4168 ( 
.A1(n_3961),
.A2(n_421),
.B(n_422),
.Y(n_4168)
);

O2A1O1Ixp33_ASAP7_75t_L g4169 ( 
.A1(n_3916),
.A2(n_424),
.B(n_421),
.C(n_423),
.Y(n_4169)
);

NAND3xp33_ASAP7_75t_L g4170 ( 
.A(n_3959),
.B(n_425),
.C(n_426),
.Y(n_4170)
);

AO21x2_ASAP7_75t_L g4171 ( 
.A1(n_3881),
.A2(n_425),
.B(n_426),
.Y(n_4171)
);

AO31x2_ASAP7_75t_L g4172 ( 
.A1(n_4153),
.A2(n_3955),
.A3(n_3921),
.B(n_3962),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_4133),
.A2(n_3918),
.B(n_3877),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_4152),
.A2(n_3885),
.B1(n_3874),
.B2(n_3991),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_4031),
.Y(n_4175)
);

AOI21x1_ASAP7_75t_L g4176 ( 
.A1(n_4124),
.A2(n_3939),
.B(n_4003),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4031),
.Y(n_4177)
);

OR2x2_ASAP7_75t_L g4178 ( 
.A(n_4100),
.B(n_3937),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4051),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4051),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4040),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4062),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4096),
.B(n_3937),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4062),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4030),
.Y(n_4185)
);

OAI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_4147),
.A2(n_3976),
.B1(n_3954),
.B2(n_3996),
.Y(n_4186)
);

AO31x2_ASAP7_75t_L g4187 ( 
.A1(n_4117),
.A2(n_3997),
.A3(n_3942),
.B(n_3949),
.Y(n_4187)
);

OA21x2_ASAP7_75t_L g4188 ( 
.A1(n_4035),
.A2(n_3957),
.B(n_4016),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4042),
.B(n_3938),
.Y(n_4189)
);

BUFx4f_ASAP7_75t_SL g4190 ( 
.A(n_4052),
.Y(n_4190)
);

OAI21x1_ASAP7_75t_L g4191 ( 
.A1(n_4020),
.A2(n_4015),
.B(n_3994),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4042),
.B(n_3899),
.Y(n_4192)
);

AO31x2_ASAP7_75t_L g4193 ( 
.A1(n_4126),
.A2(n_3997),
.A3(n_3949),
.B(n_3924),
.Y(n_4193)
);

AND2x4_ASAP7_75t_L g4194 ( 
.A(n_4036),
.B(n_4029),
.Y(n_4194)
);

OAI21x1_ASAP7_75t_L g4195 ( 
.A1(n_4020),
.A2(n_3924),
.B(n_3866),
.Y(n_4195)
);

AOI21x1_ASAP7_75t_L g4196 ( 
.A1(n_4124),
.A2(n_3936),
.B(n_3919),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4068),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4068),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4032),
.Y(n_4199)
);

AND2x4_ASAP7_75t_L g4200 ( 
.A(n_4029),
.B(n_3905),
.Y(n_4200)
);

NAND2x1p5_ASAP7_75t_L g4201 ( 
.A(n_4053),
.B(n_3907),
.Y(n_4201)
);

AND2x4_ASAP7_75t_L g4202 ( 
.A(n_4112),
.B(n_3905),
.Y(n_4202)
);

OR2x2_ASAP7_75t_L g4203 ( 
.A(n_4091),
.B(n_3895),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4045),
.Y(n_4204)
);

OAI21x1_ASAP7_75t_SL g4205 ( 
.A1(n_4115),
.A2(n_3919),
.B(n_3902),
.Y(n_4205)
);

INVx4_ASAP7_75t_L g4206 ( 
.A(n_4052),
.Y(n_4206)
);

OAI21x1_ASAP7_75t_L g4207 ( 
.A1(n_4074),
.A2(n_3947),
.B(n_3896),
.Y(n_4207)
);

HB1xp67_ASAP7_75t_L g4208 ( 
.A(n_4021),
.Y(n_4208)
);

A2O1A1Ixp33_ASAP7_75t_L g4209 ( 
.A1(n_4169),
.A2(n_3900),
.B(n_3899),
.C(n_3865),
.Y(n_4209)
);

BUFx3_ASAP7_75t_L g4210 ( 
.A(n_4052),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_4133),
.A2(n_3865),
.B(n_3900),
.Y(n_4211)
);

OAI21x1_ASAP7_75t_L g4212 ( 
.A1(n_4038),
.A2(n_3896),
.B(n_3895),
.Y(n_4212)
);

CKINVDCx20_ASAP7_75t_R g4213 ( 
.A(n_4057),
.Y(n_4213)
);

OAI21xp5_ASAP7_75t_L g4214 ( 
.A1(n_4170),
.A2(n_4158),
.B(n_4122),
.Y(n_4214)
);

AOI21xp33_ASAP7_75t_SL g4215 ( 
.A1(n_4152),
.A2(n_4168),
.B(n_4130),
.Y(n_4215)
);

A2O1A1Ixp33_ASAP7_75t_L g4216 ( 
.A1(n_4130),
.A2(n_4070),
.B(n_4142),
.C(n_4170),
.Y(n_4216)
);

AND2x4_ASAP7_75t_L g4217 ( 
.A(n_4106),
.B(n_428),
.Y(n_4217)
);

AOI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_4122),
.A2(n_428),
.B(n_429),
.Y(n_4218)
);

BUFx3_ASAP7_75t_L g4219 ( 
.A(n_4093),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4079),
.Y(n_4220)
);

AOI22xp5_ASAP7_75t_L g4221 ( 
.A1(n_4087),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_4221)
);

BUFx12f_ASAP7_75t_L g4222 ( 
.A(n_4097),
.Y(n_4222)
);

CKINVDCx12_ASAP7_75t_R g4223 ( 
.A(n_4103),
.Y(n_4223)
);

BUFx2_ASAP7_75t_L g4224 ( 
.A(n_4038),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_4150),
.B(n_432),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4088),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4042),
.B(n_432),
.Y(n_4227)
);

AO21x2_ASAP7_75t_L g4228 ( 
.A1(n_4165),
.A2(n_4149),
.B(n_4137),
.Y(n_4228)
);

OAI21x1_ASAP7_75t_L g4229 ( 
.A1(n_4056),
.A2(n_433),
.B(n_434),
.Y(n_4229)
);

HB1xp67_ASAP7_75t_L g4230 ( 
.A(n_4065),
.Y(n_4230)
);

AOI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_4158),
.A2(n_685),
.B(n_433),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4053),
.Y(n_4232)
);

AND2x4_ASAP7_75t_L g4233 ( 
.A(n_4106),
.B(n_434),
.Y(n_4233)
);

AOI22xp5_ASAP7_75t_L g4234 ( 
.A1(n_4094),
.A2(n_4168),
.B1(n_4055),
.B2(n_4123),
.Y(n_4234)
);

A2O1A1Ixp33_ASAP7_75t_L g4235 ( 
.A1(n_4142),
.A2(n_4083),
.B(n_4092),
.C(n_4161),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_4102),
.A2(n_435),
.B(n_436),
.Y(n_4236)
);

OAI21xp5_ASAP7_75t_L g4237 ( 
.A1(n_4034),
.A2(n_437),
.B(n_438),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_4102),
.A2(n_684),
.B(n_438),
.Y(n_4238)
);

OAI21x1_ASAP7_75t_L g4239 ( 
.A1(n_4050),
.A2(n_439),
.B(n_440),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4025),
.Y(n_4240)
);

AND2x2_ASAP7_75t_SL g4241 ( 
.A(n_4081),
.B(n_439),
.Y(n_4241)
);

OAI21x1_ASAP7_75t_L g4242 ( 
.A1(n_4043),
.A2(n_440),
.B(n_441),
.Y(n_4242)
);

CKINVDCx16_ASAP7_75t_R g4243 ( 
.A(n_4033),
.Y(n_4243)
);

AO21x2_ASAP7_75t_L g4244 ( 
.A1(n_4131),
.A2(n_443),
.B(n_444),
.Y(n_4244)
);

OAI21x1_ASAP7_75t_L g4245 ( 
.A1(n_4037),
.A2(n_444),
.B(n_445),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4116),
.B(n_446),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4089),
.Y(n_4247)
);

OA21x2_ASAP7_75t_L g4248 ( 
.A1(n_4035),
.A2(n_447),
.B(n_448),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4027),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_4249)
);

OAI21x1_ASAP7_75t_L g4250 ( 
.A1(n_4060),
.A2(n_449),
.B(n_450),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4064),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_4067),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4065),
.B(n_4111),
.Y(n_4253)
);

OR2x2_ASAP7_75t_L g4254 ( 
.A(n_4026),
.B(n_684),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4073),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_4141),
.B(n_451),
.Y(n_4256)
);

OAI21x1_ASAP7_75t_L g4257 ( 
.A1(n_4084),
.A2(n_451),
.B(n_452),
.Y(n_4257)
);

INVx3_ASAP7_75t_L g4258 ( 
.A(n_4019),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4090),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4119),
.A2(n_4058),
.B(n_4055),
.Y(n_4260)
);

AO31x2_ASAP7_75t_L g4261 ( 
.A1(n_4143),
.A2(n_454),
.A3(n_452),
.B(n_453),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4081),
.Y(n_4262)
);

OR2x2_ASAP7_75t_L g4263 ( 
.A(n_4022),
.B(n_453),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4157),
.B(n_454),
.Y(n_4264)
);

AOI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_4119),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4159),
.B(n_456),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4018),
.Y(n_4267)
);

OA21x2_ASAP7_75t_L g4268 ( 
.A1(n_4163),
.A2(n_457),
.B(n_458),
.Y(n_4268)
);

OAI21x1_ASAP7_75t_L g4269 ( 
.A1(n_4041),
.A2(n_458),
.B(n_459),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_4164),
.B(n_459),
.Y(n_4270)
);

AOI21x1_ASAP7_75t_L g4271 ( 
.A1(n_4131),
.A2(n_460),
.B(n_461),
.Y(n_4271)
);

OA21x2_ASAP7_75t_L g4272 ( 
.A1(n_4135),
.A2(n_461),
.B(n_462),
.Y(n_4272)
);

OAI21x1_ASAP7_75t_L g4273 ( 
.A1(n_4041),
.A2(n_462),
.B(n_463),
.Y(n_4273)
);

AOI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_4058),
.A2(n_463),
.B(n_464),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4018),
.Y(n_4275)
);

OA21x2_ASAP7_75t_L g4276 ( 
.A1(n_4135),
.A2(n_464),
.B(n_465),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4075),
.Y(n_4277)
);

OA21x2_ASAP7_75t_L g4278 ( 
.A1(n_4095),
.A2(n_465),
.B(n_466),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4075),
.Y(n_4279)
);

OAI21x1_ASAP7_75t_L g4280 ( 
.A1(n_4063),
.A2(n_466),
.B(n_467),
.Y(n_4280)
);

HB1xp67_ASAP7_75t_L g4281 ( 
.A(n_4071),
.Y(n_4281)
);

BUFx8_ASAP7_75t_L g4282 ( 
.A(n_4110),
.Y(n_4282)
);

AOI21xp5_ASAP7_75t_SL g4283 ( 
.A1(n_4166),
.A2(n_467),
.B(n_468),
.Y(n_4283)
);

AO21x2_ASAP7_75t_L g4284 ( 
.A1(n_4095),
.A2(n_468),
.B(n_469),
.Y(n_4284)
);

OA21x2_ASAP7_75t_L g4285 ( 
.A1(n_4072),
.A2(n_469),
.B(n_470),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4046),
.Y(n_4286)
);

OAI21x1_ASAP7_75t_SL g4287 ( 
.A1(n_4049),
.A2(n_470),
.B(n_471),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4046),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_L g4289 ( 
.A(n_4150),
.B(n_471),
.Y(n_4289)
);

AO31x2_ASAP7_75t_L g4290 ( 
.A1(n_4162),
.A2(n_4044),
.A3(n_4104),
.B(n_4080),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_4072),
.A2(n_683),
.B(n_472),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4156),
.B(n_472),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4071),
.Y(n_4293)
);

OR2x2_ASAP7_75t_L g4294 ( 
.A(n_4114),
.B(n_682),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4127),
.B(n_473),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4085),
.Y(n_4296)
);

INVx2_ASAP7_75t_SL g4297 ( 
.A(n_4019),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_4144),
.B(n_681),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4085),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4048),
.Y(n_4300)
);

INVx3_ASAP7_75t_L g4301 ( 
.A(n_4078),
.Y(n_4301)
);

AO21x2_ASAP7_75t_L g4302 ( 
.A1(n_4023),
.A2(n_474),
.B(n_475),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4139),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4028),
.Y(n_4304)
);

AND2x4_ASAP7_75t_L g4305 ( 
.A(n_4128),
.B(n_474),
.Y(n_4305)
);

OR2x6_ASAP7_75t_L g4306 ( 
.A(n_4066),
.B(n_4128),
.Y(n_4306)
);

OR2x6_ASAP7_75t_L g4307 ( 
.A(n_4066),
.B(n_475),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4139),
.Y(n_4308)
);

BUFx12f_ASAP7_75t_L g4309 ( 
.A(n_4110),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4108),
.A2(n_476),
.B(n_477),
.Y(n_4310)
);

HB1xp67_ASAP7_75t_L g4311 ( 
.A(n_4066),
.Y(n_4311)
);

CKINVDCx8_ASAP7_75t_R g4312 ( 
.A(n_4167),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4028),
.Y(n_4313)
);

NOR2xp33_ASAP7_75t_L g4314 ( 
.A(n_4154),
.B(n_4024),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4078),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_4166),
.Y(n_4316)
);

AOI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_4108),
.A2(n_678),
.B(n_476),
.Y(n_4317)
);

INVx2_ASAP7_75t_SL g4318 ( 
.A(n_4039),
.Y(n_4318)
);

OA21x2_ASAP7_75t_L g4319 ( 
.A1(n_4082),
.A2(n_478),
.B(n_479),
.Y(n_4319)
);

OA21x2_ASAP7_75t_L g4320 ( 
.A1(n_4098),
.A2(n_478),
.B(n_480),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4078),
.Y(n_4321)
);

BUFx4f_ASAP7_75t_L g4322 ( 
.A(n_4129),
.Y(n_4322)
);

AO21x2_ASAP7_75t_L g4323 ( 
.A1(n_4144),
.A2(n_481),
.B(n_482),
.Y(n_4323)
);

BUFx3_ASAP7_75t_L g4324 ( 
.A(n_4190),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4185),
.Y(n_4325)
);

AOI22xp33_ASAP7_75t_L g4326 ( 
.A1(n_4214),
.A2(n_4101),
.B1(n_4171),
.B2(n_4047),
.Y(n_4326)
);

BUFx4f_ASAP7_75t_SL g4327 ( 
.A(n_4213),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4314),
.B(n_4028),
.Y(n_4328)
);

INVx2_ASAP7_75t_SL g4329 ( 
.A(n_4210),
.Y(n_4329)
);

OAI22xp5_ASAP7_75t_L g4330 ( 
.A1(n_4216),
.A2(n_4234),
.B1(n_4241),
.B2(n_4221),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4185),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_4235),
.A2(n_4069),
.B1(n_4140),
.B2(n_4136),
.Y(n_4332)
);

AOI22xp33_ASAP7_75t_SL g4333 ( 
.A1(n_4186),
.A2(n_4059),
.B1(n_4054),
.B2(n_4076),
.Y(n_4333)
);

AOI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_4291),
.A2(n_4171),
.B1(n_4059),
.B2(n_4134),
.Y(n_4334)
);

INVxp67_ASAP7_75t_L g4335 ( 
.A(n_4316),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4304),
.B(n_4120),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4215),
.B(n_4120),
.Y(n_4337)
);

AOI222xp33_ASAP7_75t_L g4338 ( 
.A1(n_4249),
.A2(n_4145),
.B1(n_4113),
.B2(n_4105),
.C1(n_4148),
.C2(n_4146),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4301),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4304),
.B(n_4105),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4220),
.Y(n_4341)
);

OAI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_4173),
.A2(n_4160),
.B(n_4132),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4201),
.A2(n_4129),
.B1(n_4061),
.B2(n_4113),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_4202),
.B(n_4145),
.Y(n_4344)
);

OAI21xp5_ASAP7_75t_SL g4345 ( 
.A1(n_4174),
.A2(n_4118),
.B(n_4107),
.Y(n_4345)
);

OAI21xp33_ASAP7_75t_L g4346 ( 
.A1(n_4260),
.A2(n_4107),
.B(n_4125),
.Y(n_4346)
);

AOI22xp33_ASAP7_75t_L g4347 ( 
.A1(n_4285),
.A2(n_4155),
.B1(n_4099),
.B2(n_4109),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4301),
.Y(n_4348)
);

AOI222xp33_ASAP7_75t_L g4349 ( 
.A1(n_4237),
.A2(n_4151),
.B1(n_4077),
.B2(n_4086),
.C1(n_485),
.C2(n_486),
.Y(n_4349)
);

AOI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4285),
.A2(n_4138),
.B1(n_4121),
.B2(n_484),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4194),
.B(n_4121),
.Y(n_4351)
);

AOI22xp33_ASAP7_75t_L g4352 ( 
.A1(n_4274),
.A2(n_4121),
.B1(n_486),
.B2(n_482),
.Y(n_4352)
);

AND2x2_ASAP7_75t_L g4353 ( 
.A(n_4194),
.B(n_483),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4209),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4220),
.Y(n_4355)
);

OAI21xp5_ASAP7_75t_SL g4356 ( 
.A1(n_4231),
.A2(n_489),
.B(n_492),
.Y(n_4356)
);

OAI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_4307),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.Y(n_4357)
);

OAI21xp5_ASAP7_75t_SL g4358 ( 
.A1(n_4218),
.A2(n_494),
.B(n_495),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4226),
.Y(n_4359)
);

OAI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4307),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_4360)
);

NOR2xp33_ASAP7_75t_L g4361 ( 
.A(n_4206),
.B(n_498),
.Y(n_4361)
);

AOI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_4297),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4226),
.Y(n_4363)
);

AOI22xp33_ASAP7_75t_L g4364 ( 
.A1(n_4211),
.A2(n_499),
.B1(n_500),
.B2(n_502),
.Y(n_4364)
);

AOI222xp33_ASAP7_75t_L g4365 ( 
.A1(n_4287),
.A2(n_503),
.B1(n_505),
.B2(n_506),
.C1(n_507),
.C2(n_508),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4175),
.Y(n_4366)
);

OAI22xp33_ASAP7_75t_L g4367 ( 
.A1(n_4306),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_4367)
);

OAI22xp33_ASAP7_75t_L g4368 ( 
.A1(n_4306),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_4368)
);

AND2x2_ASAP7_75t_L g4369 ( 
.A(n_4253),
.B(n_509),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_4202),
.B(n_510),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4251),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_4254),
.B(n_511),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4199),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4204),
.Y(n_4374)
);

BUFx3_ASAP7_75t_L g4375 ( 
.A(n_4282),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_4313),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_SL g4377 ( 
.A1(n_4243),
.A2(n_512),
.B1(n_515),
.B2(n_516),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4177),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4302),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_4206),
.B(n_517),
.Y(n_4380)
);

AOI22xp33_ASAP7_75t_L g4381 ( 
.A1(n_4188),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_SL g4382 ( 
.A1(n_4322),
.A2(n_4222),
.B1(n_4276),
.B2(n_4272),
.Y(n_4382)
);

NOR2xp33_ASAP7_75t_L g4383 ( 
.A(n_4312),
.B(n_521),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_SL g4384 ( 
.A1(n_4322),
.A2(n_522),
.B1(n_523),
.B2(n_524),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_SL g4385 ( 
.A1(n_4272),
.A2(n_523),
.B1(n_525),
.B2(n_526),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_SL g4386 ( 
.A(n_4258),
.B(n_526),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4262),
.B(n_527),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4232),
.Y(n_4388)
);

OAI21xp5_ASAP7_75t_SL g4389 ( 
.A1(n_4265),
.A2(n_527),
.B(n_528),
.Y(n_4389)
);

AO22x1_ASAP7_75t_L g4390 ( 
.A1(n_4262),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_4390)
);

OAI22xp33_ASAP7_75t_L g4391 ( 
.A1(n_4227),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4247),
.Y(n_4392)
);

BUFx6f_ASAP7_75t_L g4393 ( 
.A(n_4305),
.Y(n_4393)
);

HB1xp67_ASAP7_75t_L g4394 ( 
.A(n_4230),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4255),
.Y(n_4395)
);

OAI21xp5_ASAP7_75t_SL g4396 ( 
.A1(n_4310),
.A2(n_531),
.B(n_532),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4258),
.B(n_532),
.Y(n_4397)
);

AOI22xp33_ASAP7_75t_L g4398 ( 
.A1(n_4188),
.A2(n_533),
.B1(n_534),
.B2(n_535),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_L g4399 ( 
.A1(n_4317),
.A2(n_535),
.B1(n_536),
.B2(n_537),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4228),
.Y(n_4400)
);

AOI22xp33_ASAP7_75t_L g4401 ( 
.A1(n_4183),
.A2(n_536),
.B1(n_538),
.B2(n_539),
.Y(n_4401)
);

OAI21xp33_ASAP7_75t_L g4402 ( 
.A1(n_4283),
.A2(n_540),
.B(n_542),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_4236),
.A2(n_543),
.B1(n_544),
.B2(n_545),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_L g4404 ( 
.A1(n_4238),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_4404)
);

AOI222xp33_ASAP7_75t_L g4405 ( 
.A1(n_4264),
.A2(n_4270),
.B1(n_4266),
.B2(n_4299),
.C1(n_4296),
.C2(n_4205),
.Y(n_4405)
);

BUFx2_ASAP7_75t_L g4406 ( 
.A(n_4309),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4268),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_SL g4408 ( 
.A1(n_4276),
.A2(n_678),
.B1(n_549),
.B2(n_550),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4311),
.B(n_546),
.Y(n_4409)
);

OR2x2_ASAP7_75t_L g4410 ( 
.A(n_4203),
.B(n_550),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4244),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.Y(n_4411)
);

HB1xp67_ASAP7_75t_L g4412 ( 
.A(n_4208),
.Y(n_4412)
);

AOI22xp33_ASAP7_75t_SL g4413 ( 
.A1(n_4278),
.A2(n_677),
.B1(n_552),
.B2(n_553),
.Y(n_4413)
);

AOI21xp5_ASAP7_75t_L g4414 ( 
.A1(n_4189),
.A2(n_551),
.B(n_554),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4176),
.A2(n_4196),
.B1(n_4268),
.B2(n_4278),
.Y(n_4415)
);

OAI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4248),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4197),
.Y(n_4417)
);

AOI22xp33_ASAP7_75t_L g4418 ( 
.A1(n_4224),
.A2(n_555),
.B1(n_556),
.B2(n_557),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4284),
.B(n_557),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_4198),
.Y(n_4420)
);

AND2x2_ASAP7_75t_L g4421 ( 
.A(n_4315),
.B(n_558),
.Y(n_4421)
);

BUFx4f_ASAP7_75t_SL g4422 ( 
.A(n_4282),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4248),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_4219),
.Y(n_4424)
);

BUFx2_ASAP7_75t_L g4425 ( 
.A(n_4200),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4321),
.B(n_558),
.Y(n_4426)
);

AOI211xp5_ASAP7_75t_L g4427 ( 
.A1(n_4281),
.A2(n_560),
.B(n_561),
.C(n_563),
.Y(n_4427)
);

BUFx6f_ASAP7_75t_L g4428 ( 
.A(n_4305),
.Y(n_4428)
);

CKINVDCx20_ASAP7_75t_R g4429 ( 
.A(n_4223),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4240),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4252),
.Y(n_4431)
);

OAI22xp5_ASAP7_75t_SL g4432 ( 
.A1(n_4225),
.A2(n_560),
.B1(n_561),
.B2(n_563),
.Y(n_4432)
);

AOI22xp33_ASAP7_75t_L g4433 ( 
.A1(n_4178),
.A2(n_565),
.B1(n_566),
.B2(n_567),
.Y(n_4433)
);

AOI22xp33_ASAP7_75t_SL g4434 ( 
.A1(n_4323),
.A2(n_565),
.B1(n_566),
.B2(n_567),
.Y(n_4434)
);

AOI22xp33_ASAP7_75t_L g4435 ( 
.A1(n_4319),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.Y(n_4435)
);

AOI22xp33_ASAP7_75t_L g4436 ( 
.A1(n_4319),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.Y(n_4436)
);

OAI222xp33_ASAP7_75t_L g4437 ( 
.A1(n_4271),
.A2(n_571),
.B1(n_572),
.B2(n_573),
.C1(n_574),
.C2(n_575),
.Y(n_4437)
);

OAI22xp5_ASAP7_75t_L g4438 ( 
.A1(n_4298),
.A2(n_572),
.B1(n_573),
.B2(n_577),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4179),
.B(n_4180),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4192),
.Y(n_4440)
);

AOI22xp33_ASAP7_75t_L g4441 ( 
.A1(n_4320),
.A2(n_577),
.B1(n_578),
.B2(n_579),
.Y(n_4441)
);

AOI22xp33_ASAP7_75t_L g4442 ( 
.A1(n_4320),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4303),
.B(n_580),
.Y(n_4443)
);

AOI22xp33_ASAP7_75t_L g4444 ( 
.A1(n_4300),
.A2(n_581),
.B1(n_582),
.B2(n_584),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4259),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4179),
.B(n_581),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4269),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4273),
.Y(n_4448)
);

AND2x4_ASAP7_75t_L g4449 ( 
.A(n_4200),
.B(n_582),
.Y(n_4449)
);

AOI22xp33_ASAP7_75t_L g4450 ( 
.A1(n_4300),
.A2(n_4207),
.B1(n_4289),
.B2(n_4318),
.Y(n_4450)
);

HB1xp67_ASAP7_75t_L g4451 ( 
.A(n_4212),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4308),
.B(n_584),
.Y(n_4452)
);

BUFx2_ASAP7_75t_L g4453 ( 
.A(n_4217),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4181),
.Y(n_4454)
);

NAND3xp33_ASAP7_75t_L g4455 ( 
.A(n_4293),
.B(n_585),
.C(n_586),
.Y(n_4455)
);

OAI22xp5_ASAP7_75t_L g4456 ( 
.A1(n_4263),
.A2(n_585),
.B1(n_586),
.B2(n_587),
.Y(n_4456)
);

BUFx6f_ASAP7_75t_L g4457 ( 
.A(n_4217),
.Y(n_4457)
);

INVx3_ASAP7_75t_L g4458 ( 
.A(n_4233),
.Y(n_4458)
);

OAI21xp33_ASAP7_75t_L g4459 ( 
.A1(n_4293),
.A2(n_587),
.B(n_588),
.Y(n_4459)
);

OAI21xp5_ASAP7_75t_SL g4460 ( 
.A1(n_4292),
.A2(n_588),
.B(n_589),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_4246),
.B(n_589),
.Y(n_4461)
);

AOI222xp33_ASAP7_75t_L g4462 ( 
.A1(n_4256),
.A2(n_590),
.B1(n_591),
.B2(n_592),
.C1(n_593),
.C2(n_595),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4267),
.B(n_590),
.Y(n_4463)
);

OAI21xp33_ASAP7_75t_L g4464 ( 
.A1(n_4286),
.A2(n_591),
.B(n_593),
.Y(n_4464)
);

OAI22xp5_ASAP7_75t_L g4465 ( 
.A1(n_4294),
.A2(n_595),
.B1(n_596),
.B2(n_598),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4267),
.Y(n_4466)
);

AOI22xp33_ASAP7_75t_L g4467 ( 
.A1(n_4195),
.A2(n_599),
.B1(n_600),
.B2(n_601),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4275),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4275),
.Y(n_4469)
);

NOR2xp33_ASAP7_75t_L g4470 ( 
.A(n_4295),
.B(n_599),
.Y(n_4470)
);

HB1xp67_ASAP7_75t_L g4471 ( 
.A(n_4245),
.Y(n_4471)
);

AOI22xp33_ASAP7_75t_L g4472 ( 
.A1(n_4191),
.A2(n_601),
.B1(n_602),
.B2(n_604),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4277),
.Y(n_4473)
);

OAI22xp33_ASAP7_75t_L g4474 ( 
.A1(n_4286),
.A2(n_4288),
.B1(n_4277),
.B2(n_4279),
.Y(n_4474)
);

BUFx2_ASAP7_75t_L g4475 ( 
.A(n_4429),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4449),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4325),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4449),
.Y(n_4478)
);

AO21x2_ASAP7_75t_L g4479 ( 
.A1(n_4400),
.A2(n_4474),
.B(n_4407),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4425),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4453),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4473),
.Y(n_4482)
);

AOI21x1_ASAP7_75t_L g4483 ( 
.A1(n_4406),
.A2(n_4288),
.B(n_4233),
.Y(n_4483)
);

AO21x2_ASAP7_75t_L g4484 ( 
.A1(n_4415),
.A2(n_4279),
.B(n_4242),
.Y(n_4484)
);

OR2x6_ASAP7_75t_L g4485 ( 
.A(n_4354),
.B(n_4280),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4331),
.Y(n_4486)
);

HB1xp67_ASAP7_75t_L g4487 ( 
.A(n_4394),
.Y(n_4487)
);

OR2x2_ASAP7_75t_L g4488 ( 
.A(n_4336),
.B(n_4180),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4393),
.Y(n_4489)
);

INVxp33_ASAP7_75t_L g4490 ( 
.A(n_4382),
.Y(n_4490)
);

HB1xp67_ASAP7_75t_L g4491 ( 
.A(n_4412),
.Y(n_4491)
);

OR2x2_ASAP7_75t_L g4492 ( 
.A(n_4336),
.B(n_4182),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_4422),
.B(n_4229),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_4341),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4393),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4355),
.Y(n_4496)
);

OAI21xp5_ASAP7_75t_L g4497 ( 
.A1(n_4330),
.A2(n_4250),
.B(n_4239),
.Y(n_4497)
);

OA21x2_ASAP7_75t_L g4498 ( 
.A1(n_4328),
.A2(n_4182),
.B(n_4184),
.Y(n_4498)
);

NOR2xp33_ASAP7_75t_L g4499 ( 
.A(n_4375),
.B(n_4257),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4393),
.Y(n_4500)
);

AOI22xp33_ASAP7_75t_L g4501 ( 
.A1(n_4330),
.A2(n_4184),
.B1(n_4290),
.B2(n_4172),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4359),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4363),
.Y(n_4503)
);

HB1xp67_ASAP7_75t_L g4504 ( 
.A(n_4335),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4371),
.Y(n_4505)
);

BUFx6f_ASAP7_75t_L g4506 ( 
.A(n_4324),
.Y(n_4506)
);

AO21x2_ASAP7_75t_L g4507 ( 
.A1(n_4415),
.A2(n_4387),
.B(n_4423),
.Y(n_4507)
);

INVxp67_ASAP7_75t_SL g4508 ( 
.A(n_4428),
.Y(n_4508)
);

AO21x2_ASAP7_75t_L g4509 ( 
.A1(n_4387),
.A2(n_4261),
.B(n_4187),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4351),
.B(n_4172),
.Y(n_4510)
);

AO21x2_ASAP7_75t_L g4511 ( 
.A1(n_4354),
.A2(n_4261),
.B(n_4187),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4428),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4339),
.B(n_4172),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4348),
.B(n_4290),
.Y(n_4514)
);

AND2x4_ASAP7_75t_L g4515 ( 
.A(n_4458),
.B(n_4261),
.Y(n_4515)
);

OA21x2_ASAP7_75t_L g4516 ( 
.A1(n_4450),
.A2(n_4187),
.B(n_4290),
.Y(n_4516)
);

HB1xp67_ASAP7_75t_L g4517 ( 
.A(n_4471),
.Y(n_4517)
);

INVx2_ASAP7_75t_L g4518 ( 
.A(n_4428),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4373),
.Y(n_4519)
);

INVx3_ASAP7_75t_L g4520 ( 
.A(n_4457),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4458),
.Y(n_4521)
);

HB1xp67_ASAP7_75t_L g4522 ( 
.A(n_4447),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4457),
.Y(n_4523)
);

AND2x4_ASAP7_75t_L g4524 ( 
.A(n_4466),
.B(n_4469),
.Y(n_4524)
);

AOI21xp5_ASAP7_75t_SL g4525 ( 
.A1(n_4402),
.A2(n_4193),
.B(n_606),
.Y(n_4525)
);

INVxp67_ASAP7_75t_L g4526 ( 
.A(n_4370),
.Y(n_4526)
);

AOI22xp33_ASAP7_75t_L g4527 ( 
.A1(n_4333),
.A2(n_4193),
.B1(n_606),
.B2(n_607),
.Y(n_4527)
);

BUFx2_ASAP7_75t_L g4528 ( 
.A(n_4457),
.Y(n_4528)
);

INVxp33_ASAP7_75t_L g4529 ( 
.A(n_4337),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4374),
.Y(n_4530)
);

INVx1_ASAP7_75t_SL g4531 ( 
.A(n_4327),
.Y(n_4531)
);

OR2x2_ASAP7_75t_L g4532 ( 
.A(n_4340),
.B(n_4193),
.Y(n_4532)
);

BUFx3_ASAP7_75t_L g4533 ( 
.A(n_4329),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4405),
.B(n_605),
.Y(n_4534)
);

INVxp33_ASAP7_75t_L g4535 ( 
.A(n_4343),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4392),
.Y(n_4536)
);

AO21x2_ASAP7_75t_L g4537 ( 
.A1(n_4451),
.A2(n_608),
.B(n_609),
.Y(n_4537)
);

INVx3_ASAP7_75t_L g4538 ( 
.A(n_4468),
.Y(n_4538)
);

AO21x2_ASAP7_75t_L g4539 ( 
.A1(n_4419),
.A2(n_608),
.B(n_610),
.Y(n_4539)
);

BUFx8_ASAP7_75t_SL g4540 ( 
.A(n_4397),
.Y(n_4540)
);

AO31x2_ASAP7_75t_L g4541 ( 
.A1(n_4416),
.A2(n_610),
.A3(n_611),
.B(n_612),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4366),
.B(n_4378),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4388),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4417),
.Y(n_4544)
);

BUFx3_ASAP7_75t_L g4545 ( 
.A(n_4424),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4420),
.B(n_611),
.Y(n_4546)
);

HB1xp67_ASAP7_75t_L g4547 ( 
.A(n_4448),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4454),
.B(n_612),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4395),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4430),
.Y(n_4550)
);

HB1xp67_ASAP7_75t_L g4551 ( 
.A(n_4410),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4338),
.B(n_613),
.Y(n_4552)
);

CKINVDCx6p67_ASAP7_75t_R g4553 ( 
.A(n_4386),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4344),
.B(n_613),
.Y(n_4554)
);

BUFx3_ASAP7_75t_L g4555 ( 
.A(n_4353),
.Y(n_4555)
);

INVxp67_ASAP7_75t_L g4556 ( 
.A(n_4343),
.Y(n_4556)
);

INVx3_ASAP7_75t_L g4557 ( 
.A(n_4431),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4445),
.Y(n_4558)
);

NOR2xp33_ASAP7_75t_L g4559 ( 
.A(n_4345),
.B(n_614),
.Y(n_4559)
);

NOR2xp33_ASAP7_75t_L g4560 ( 
.A(n_4361),
.B(n_615),
.Y(n_4560)
);

OR2x6_ASAP7_75t_L g4561 ( 
.A(n_4390),
.B(n_616),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4446),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4440),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4446),
.Y(n_4564)
);

AND2x4_ASAP7_75t_L g4565 ( 
.A(n_4342),
.B(n_616),
.Y(n_4565)
);

AO21x2_ASAP7_75t_L g4566 ( 
.A1(n_4416),
.A2(n_4414),
.B(n_4391),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4340),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4439),
.Y(n_4568)
);

INVx2_ASAP7_75t_L g4569 ( 
.A(n_4439),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4443),
.Y(n_4570)
);

BUFx2_ASAP7_75t_L g4571 ( 
.A(n_4342),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4452),
.Y(n_4572)
);

AO21x2_ASAP7_75t_L g4573 ( 
.A1(n_4455),
.A2(n_617),
.B(n_618),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_4346),
.B(n_617),
.Y(n_4574)
);

AOI21x1_ASAP7_75t_L g4575 ( 
.A1(n_4409),
.A2(n_618),
.B(n_619),
.Y(n_4575)
);

BUFx6f_ASAP7_75t_L g4576 ( 
.A(n_4421),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4426),
.Y(n_4577)
);

CKINVDCx5p33_ASAP7_75t_R g4578 ( 
.A(n_4432),
.Y(n_4578)
);

INVxp33_ASAP7_75t_L g4579 ( 
.A(n_4380),
.Y(n_4579)
);

AO21x2_ASAP7_75t_L g4580 ( 
.A1(n_4367),
.A2(n_619),
.B(n_620),
.Y(n_4580)
);

BUFx6f_ASAP7_75t_L g4581 ( 
.A(n_4463),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4369),
.Y(n_4582)
);

AO21x2_ASAP7_75t_L g4583 ( 
.A1(n_4368),
.A2(n_620),
.B(n_621),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4372),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_4350),
.Y(n_4585)
);

AND2x4_ASAP7_75t_L g4586 ( 
.A(n_4347),
.B(n_621),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4461),
.Y(n_4587)
);

NOR2xp33_ASAP7_75t_L g4588 ( 
.A(n_4460),
.B(n_622),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4470),
.Y(n_4589)
);

OR2x2_ASAP7_75t_L g4590 ( 
.A(n_4334),
.B(n_4467),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4456),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4456),
.Y(n_4592)
);

INVx2_ASAP7_75t_SL g4593 ( 
.A(n_4357),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4465),
.Y(n_4594)
);

BUFx3_ASAP7_75t_L g4595 ( 
.A(n_4383),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4465),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_4326),
.B(n_4381),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4438),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4398),
.B(n_623),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4438),
.Y(n_4600)
);

INVx4_ASAP7_75t_L g4601 ( 
.A(n_4437),
.Y(n_4601)
);

BUFx3_ASAP7_75t_L g4602 ( 
.A(n_4362),
.Y(n_4602)
);

OA21x2_ASAP7_75t_L g4603 ( 
.A1(n_4389),
.A2(n_624),
.B(n_625),
.Y(n_4603)
);

HB1xp67_ASAP7_75t_L g4604 ( 
.A(n_4357),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4413),
.Y(n_4605)
);

OA21x2_ASAP7_75t_L g4606 ( 
.A1(n_4459),
.A2(n_624),
.B(n_625),
.Y(n_4606)
);

INVx2_ASAP7_75t_L g4607 ( 
.A(n_4332),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4385),
.B(n_626),
.Y(n_4608)
);

AO21x2_ASAP7_75t_L g4609 ( 
.A1(n_4360),
.A2(n_626),
.B(n_627),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4408),
.Y(n_4610)
);

OR2x2_ASAP7_75t_L g4611 ( 
.A(n_4435),
.B(n_628),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4472),
.B(n_628),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4545),
.Y(n_4613)
);

INVx1_ASAP7_75t_SL g4614 ( 
.A(n_4540),
.Y(n_4614)
);

HB1xp67_ASAP7_75t_L g4615 ( 
.A(n_4487),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4545),
.Y(n_4616)
);

NOR2x1_ASAP7_75t_L g4617 ( 
.A(n_4537),
.B(n_4360),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4508),
.B(n_4434),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4479),
.Y(n_4619)
);

OR2x6_ASAP7_75t_L g4620 ( 
.A(n_4525),
.B(n_4356),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4479),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4528),
.B(n_4349),
.Y(n_4622)
);

BUFx2_ASAP7_75t_L g4623 ( 
.A(n_4479),
.Y(n_4623)
);

AOI22xp5_ASAP7_75t_L g4624 ( 
.A1(n_4601),
.A2(n_4332),
.B1(n_4358),
.B2(n_4427),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4520),
.B(n_4436),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4520),
.B(n_4441),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4491),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4482),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4520),
.B(n_4442),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4533),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4533),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4601),
.B(n_4574),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4481),
.B(n_4364),
.Y(n_4633)
);

INVx2_ASAP7_75t_SL g4634 ( 
.A(n_4506),
.Y(n_4634)
);

INVx3_ASAP7_75t_L g4635 ( 
.A(n_4506),
.Y(n_4635)
);

AND2x4_ASAP7_75t_L g4636 ( 
.A(n_4521),
.B(n_4379),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4482),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4481),
.B(n_4411),
.Y(n_4638)
);

HB1xp67_ASAP7_75t_L g4639 ( 
.A(n_4581),
.Y(n_4639)
);

HB1xp67_ASAP7_75t_L g4640 ( 
.A(n_4581),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4581),
.Y(n_4641)
);

BUFx2_ASAP7_75t_L g4642 ( 
.A(n_4561),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4581),
.Y(n_4643)
);

INVx3_ASAP7_75t_L g4644 ( 
.A(n_4506),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4489),
.B(n_4418),
.Y(n_4645)
);

INVx3_ASAP7_75t_L g4646 ( 
.A(n_4506),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4477),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4576),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4486),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4489),
.B(n_4433),
.Y(n_4650)
);

INVx1_ASAP7_75t_SL g4651 ( 
.A(n_4540),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_L g4652 ( 
.A(n_4601),
.B(n_4462),
.Y(n_4652)
);

AND2x4_ASAP7_75t_L g4653 ( 
.A(n_4521),
.B(n_4401),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4576),
.Y(n_4654)
);

NOR2xp33_ASAP7_75t_L g4655 ( 
.A(n_4475),
.B(n_4396),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4574),
.B(n_4365),
.Y(n_4656)
);

AND2x2_ASAP7_75t_L g4657 ( 
.A(n_4495),
.B(n_4500),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4495),
.B(n_4377),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4494),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4600),
.B(n_4464),
.Y(n_4660)
);

BUFx6f_ASAP7_75t_L g4661 ( 
.A(n_4537),
.Y(n_4661)
);

HB1xp67_ASAP7_75t_L g4662 ( 
.A(n_4517),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4500),
.B(n_4352),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4600),
.B(n_4403),
.Y(n_4664)
);

HB1xp67_ASAP7_75t_L g4665 ( 
.A(n_4551),
.Y(n_4665)
);

HB1xp67_ASAP7_75t_L g4666 ( 
.A(n_4480),
.Y(n_4666)
);

INVx2_ASAP7_75t_SL g4667 ( 
.A(n_4515),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4512),
.B(n_4404),
.Y(n_4668)
);

HB1xp67_ASAP7_75t_L g4669 ( 
.A(n_4480),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4576),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4512),
.B(n_4384),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4518),
.B(n_4399),
.Y(n_4672)
);

HB1xp67_ASAP7_75t_L g4673 ( 
.A(n_4504),
.Y(n_4673)
);

OR2x2_ASAP7_75t_L g4674 ( 
.A(n_4593),
.B(n_4511),
.Y(n_4674)
);

INVxp67_ASAP7_75t_SL g4675 ( 
.A(n_4576),
.Y(n_4675)
);

INVx2_ASAP7_75t_L g4676 ( 
.A(n_4483),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4518),
.B(n_4523),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4523),
.B(n_4376),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4510),
.B(n_4444),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4496),
.Y(n_4680)
);

AND2x4_ASAP7_75t_L g4681 ( 
.A(n_4515),
.B(n_629),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4510),
.B(n_630),
.Y(n_4682)
);

INVx2_ASAP7_75t_L g4683 ( 
.A(n_4555),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4502),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4503),
.Y(n_4685)
);

INVxp67_ASAP7_75t_L g4686 ( 
.A(n_4561),
.Y(n_4686)
);

OR2x2_ASAP7_75t_L g4687 ( 
.A(n_4593),
.B(n_631),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4565),
.B(n_631),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4511),
.B(n_633),
.Y(n_4689)
);

OR2x2_ASAP7_75t_L g4690 ( 
.A(n_4511),
.B(n_633),
.Y(n_4690)
);

INVx3_ASAP7_75t_L g4691 ( 
.A(n_4537),
.Y(n_4691)
);

HB1xp67_ASAP7_75t_L g4692 ( 
.A(n_4476),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4565),
.B(n_634),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4505),
.Y(n_4694)
);

BUFx6f_ASAP7_75t_L g4695 ( 
.A(n_4609),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4565),
.B(n_635),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_4605),
.B(n_636),
.Y(n_4697)
);

BUFx3_ASAP7_75t_L g4698 ( 
.A(n_4561),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4519),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4476),
.B(n_636),
.Y(n_4700)
);

NOR2x1_ASAP7_75t_L g4701 ( 
.A(n_4534),
.B(n_637),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4478),
.B(n_637),
.Y(n_4702)
);

AND2x2_ASAP7_75t_SL g4703 ( 
.A(n_4571),
.B(n_638),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4530),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4478),
.B(n_638),
.Y(n_4705)
);

BUFx2_ASAP7_75t_L g4706 ( 
.A(n_4561),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4542),
.B(n_639),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4536),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4542),
.B(n_639),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4514),
.B(n_640),
.Y(n_4710)
);

OA21x2_ASAP7_75t_L g4711 ( 
.A1(n_4527),
.A2(n_640),
.B(n_641),
.Y(n_4711)
);

INVx2_ASAP7_75t_L g4712 ( 
.A(n_4555),
.Y(n_4712)
);

BUFx6f_ASAP7_75t_L g4713 ( 
.A(n_4609),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4549),
.Y(n_4714)
);

HB1xp67_ASAP7_75t_L g4715 ( 
.A(n_4538),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4515),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4538),
.Y(n_4717)
);

INVxp67_ASAP7_75t_L g4718 ( 
.A(n_4595),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4538),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4507),
.Y(n_4720)
);

INVx3_ASAP7_75t_L g4721 ( 
.A(n_4507),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_4507),
.Y(n_4722)
);

AO31x2_ASAP7_75t_L g4723 ( 
.A1(n_4552),
.A2(n_643),
.A3(n_644),
.B(n_645),
.Y(n_4723)
);

HB1xp67_ASAP7_75t_L g4724 ( 
.A(n_4698),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4665),
.Y(n_4725)
);

AND2x4_ASAP7_75t_L g4726 ( 
.A(n_4635),
.B(n_4524),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4673),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4623),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_4624),
.B(n_4490),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4623),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4642),
.B(n_4514),
.Y(n_4731)
);

OR2x2_ASAP7_75t_L g4732 ( 
.A(n_4689),
.B(n_4604),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4642),
.B(n_4513),
.Y(n_4733)
);

OR2x2_ASAP7_75t_L g4734 ( 
.A(n_4689),
.B(n_4607),
.Y(n_4734)
);

INVx2_ASAP7_75t_L g4735 ( 
.A(n_4721),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_L g4736 ( 
.A(n_4614),
.B(n_4579),
.Y(n_4736)
);

AND2x4_ASAP7_75t_L g4737 ( 
.A(n_4635),
.B(n_4524),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4706),
.B(n_4613),
.Y(n_4738)
);

INVx2_ASAP7_75t_L g4739 ( 
.A(n_4721),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4703),
.B(n_4597),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4721),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4703),
.B(n_4597),
.Y(n_4742)
);

AND2x4_ASAP7_75t_L g4743 ( 
.A(n_4635),
.B(n_4524),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4619),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4706),
.B(n_4613),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4616),
.B(n_4513),
.Y(n_4746)
);

HB1xp67_ASAP7_75t_L g4747 ( 
.A(n_4698),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4616),
.B(n_4556),
.Y(n_4748)
);

INVxp67_ASAP7_75t_SL g4749 ( 
.A(n_4644),
.Y(n_4749)
);

AND2x2_ASAP7_75t_L g4750 ( 
.A(n_4630),
.B(n_4535),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4703),
.B(n_4585),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4615),
.Y(n_4752)
);

INVxp67_ASAP7_75t_SL g4753 ( 
.A(n_4644),
.Y(n_4753)
);

BUFx2_ASAP7_75t_L g4754 ( 
.A(n_4620),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4630),
.B(n_4535),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4692),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4619),
.Y(n_4757)
);

INVx2_ASAP7_75t_L g4758 ( 
.A(n_4621),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4621),
.Y(n_4759)
);

INVx3_ASAP7_75t_L g4760 ( 
.A(n_4695),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4715),
.Y(n_4761)
);

BUFx6f_ASAP7_75t_L g4762 ( 
.A(n_4690),
.Y(n_4762)
);

HB1xp67_ASAP7_75t_L g4763 ( 
.A(n_4698),
.Y(n_4763)
);

AND2x4_ASAP7_75t_L g4764 ( 
.A(n_4644),
.B(n_4582),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4686),
.B(n_4585),
.Y(n_4765)
);

BUFx6f_ASAP7_75t_L g4766 ( 
.A(n_4690),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4675),
.B(n_4578),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4661),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4631),
.B(n_4562),
.Y(n_4769)
);

AOI22xp33_ASAP7_75t_L g4770 ( 
.A1(n_4652),
.A2(n_4490),
.B1(n_4607),
.B2(n_4566),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4720),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4720),
.Y(n_4772)
);

INVxp67_ASAP7_75t_L g4773 ( 
.A(n_4614),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4631),
.B(n_4564),
.Y(n_4774)
);

AND2x2_ASAP7_75t_L g4775 ( 
.A(n_4651),
.B(n_4589),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_4651),
.B(n_4589),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4722),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4624),
.B(n_4578),
.Y(n_4778)
);

NAND2xp5_ASAP7_75t_L g4779 ( 
.A(n_4658),
.B(n_4634),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4666),
.Y(n_4780)
);

CKINVDCx14_ASAP7_75t_R g4781 ( 
.A(n_4646),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4661),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4661),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4634),
.B(n_4543),
.Y(n_4784)
);

INVx1_ASAP7_75t_SL g4785 ( 
.A(n_4687),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4669),
.Y(n_4786)
);

OR2x2_ASAP7_75t_L g4787 ( 
.A(n_4674),
.B(n_4509),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4618),
.B(n_4543),
.Y(n_4788)
);

OR2x2_ASAP7_75t_L g4789 ( 
.A(n_4674),
.B(n_4509),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4662),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4775),
.B(n_4646),
.Y(n_4791)
);

OR2x2_ASAP7_75t_L g4792 ( 
.A(n_4732),
.B(n_4695),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4730),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4773),
.B(n_4658),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4730),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4760),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4724),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4747),
.Y(n_4798)
);

INVxp67_ASAP7_75t_L g4799 ( 
.A(n_4736),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4775),
.B(n_4646),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4763),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4762),
.Y(n_4802)
);

NAND3xp33_ASAP7_75t_L g4803 ( 
.A(n_4770),
.B(n_4713),
.C(n_4695),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4760),
.Y(n_4804)
);

AND2x2_ASAP7_75t_L g4805 ( 
.A(n_4776),
.B(n_4618),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4776),
.B(n_4738),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4762),
.Y(n_4807)
);

NAND2xp33_ASAP7_75t_SL g4808 ( 
.A(n_4762),
.B(n_4695),
.Y(n_4808)
);

AND2x2_ASAP7_75t_L g4809 ( 
.A(n_4738),
.B(n_4657),
.Y(n_4809)
);

INVx2_ASAP7_75t_L g4810 ( 
.A(n_4760),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4762),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4762),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4766),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4741),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4741),
.Y(n_4815)
);

AND2x2_ASAP7_75t_L g4816 ( 
.A(n_4745),
.B(n_4657),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4745),
.B(n_4750),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4750),
.B(n_4677),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4755),
.B(n_4671),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4766),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4735),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4755),
.B(n_4671),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4735),
.Y(n_4823)
);

AND2x2_ASAP7_75t_L g4824 ( 
.A(n_4788),
.B(n_4781),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4785),
.B(n_4718),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4739),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4739),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4788),
.B(n_4682),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4766),
.Y(n_4829)
);

INVx2_ASAP7_75t_L g4830 ( 
.A(n_4766),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4766),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4726),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_SL g4833 ( 
.A(n_4740),
.B(n_4695),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4749),
.Y(n_4834)
);

HB1xp67_ASAP7_75t_L g4835 ( 
.A(n_4726),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4748),
.B(n_4682),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4748),
.B(n_4639),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4746),
.B(n_4677),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4754),
.B(n_4640),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4753),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4728),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4746),
.B(n_4683),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4754),
.B(n_4683),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4728),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4733),
.B(n_4712),
.Y(n_4845)
);

AND2x2_ASAP7_75t_L g4846 ( 
.A(n_4733),
.B(n_4712),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_4806),
.B(n_4641),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4812),
.Y(n_4848)
);

AND2x4_ASAP7_75t_L g4849 ( 
.A(n_4812),
.B(n_4726),
.Y(n_4849)
);

NAND4xp25_ASAP7_75t_SL g4850 ( 
.A(n_4803),
.B(n_4632),
.C(n_4778),
.D(n_4617),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4830),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4830),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4806),
.B(n_4641),
.Y(n_4853)
);

INVxp67_ASAP7_75t_SL g4854 ( 
.A(n_4835),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_4805),
.B(n_4791),
.Y(n_4855)
);

INVx1_ASAP7_75t_SL g4856 ( 
.A(n_4805),
.Y(n_4856)
);

AND2x2_ASAP7_75t_L g4857 ( 
.A(n_4791),
.B(n_4643),
.Y(n_4857)
);

HB1xp67_ASAP7_75t_L g4858 ( 
.A(n_4800),
.Y(n_4858)
);

AND2x2_ASAP7_75t_L g4859 ( 
.A(n_4800),
.B(n_4643),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4792),
.Y(n_4860)
);

BUFx3_ASAP7_75t_L g4861 ( 
.A(n_4802),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4809),
.B(n_4622),
.Y(n_4862)
);

AND2x2_ASAP7_75t_L g4863 ( 
.A(n_4809),
.B(n_4648),
.Y(n_4863)
);

INVx1_ASAP7_75t_SL g4864 ( 
.A(n_4816),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4802),
.Y(n_4865)
);

HB1xp67_ASAP7_75t_L g4866 ( 
.A(n_4816),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4824),
.B(n_4648),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4792),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4807),
.Y(n_4869)
);

AND2x4_ASAP7_75t_L g4870 ( 
.A(n_4807),
.B(n_4737),
.Y(n_4870)
);

OR2x2_ASAP7_75t_L g4871 ( 
.A(n_4811),
.B(n_4732),
.Y(n_4871)
);

AND2x2_ASAP7_75t_L g4872 ( 
.A(n_4824),
.B(n_4654),
.Y(n_4872)
);

INVx1_ASAP7_75t_SL g4873 ( 
.A(n_4818),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4811),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4818),
.B(n_4654),
.Y(n_4875)
);

INVx2_ASAP7_75t_L g4876 ( 
.A(n_4813),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_4845),
.B(n_4670),
.Y(n_4877)
);

OR2x2_ASAP7_75t_L g4878 ( 
.A(n_4813),
.B(n_4661),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4820),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_4845),
.B(n_4622),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4846),
.B(n_4670),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4820),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4829),
.Y(n_4883)
);

AND2x2_ASAP7_75t_L g4884 ( 
.A(n_4846),
.B(n_4731),
.Y(n_4884)
);

OR2x6_ASAP7_75t_SL g4885 ( 
.A(n_4794),
.B(n_4767),
.Y(n_4885)
);

OR2x2_ASAP7_75t_L g4886 ( 
.A(n_4831),
.B(n_4661),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4838),
.Y(n_4887)
);

HB1xp67_ASAP7_75t_L g4888 ( 
.A(n_4832),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4838),
.Y(n_4889)
);

INVx2_ASAP7_75t_L g4890 ( 
.A(n_4832),
.Y(n_4890)
);

OR2x2_ASAP7_75t_L g4891 ( 
.A(n_4828),
.B(n_4713),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4842),
.B(n_4731),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4842),
.B(n_4638),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4844),
.Y(n_4894)
);

AND2x4_ASAP7_75t_L g4895 ( 
.A(n_4843),
.B(n_4737),
.Y(n_4895)
);

NAND2x1p5_ASAP7_75t_L g4896 ( 
.A(n_4860),
.B(n_4617),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4893),
.B(n_4799),
.Y(n_4897)
);

BUFx2_ASAP7_75t_L g4898 ( 
.A(n_4895),
.Y(n_4898)
);

NAND2x1_ASAP7_75t_L g4899 ( 
.A(n_4895),
.B(n_4737),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4893),
.B(n_4817),
.Y(n_4900)
);

INVx3_ASAP7_75t_L g4901 ( 
.A(n_4895),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4858),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4866),
.Y(n_4903)
);

OR2x2_ASAP7_75t_L g4904 ( 
.A(n_4856),
.B(n_4819),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4861),
.Y(n_4905)
);

OR2x2_ASAP7_75t_L g4906 ( 
.A(n_4864),
.B(n_4822),
.Y(n_4906)
);

INVx2_ASAP7_75t_SL g4907 ( 
.A(n_4895),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4854),
.B(n_4729),
.Y(n_4908)
);

OAI22xp5_ASAP7_75t_L g4909 ( 
.A1(n_4885),
.A2(n_4620),
.B1(n_4553),
.B2(n_4713),
.Y(n_4909)
);

BUFx6f_ASAP7_75t_L g4910 ( 
.A(n_4861),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4861),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4855),
.Y(n_4912)
);

OR2x2_ASAP7_75t_L g4913 ( 
.A(n_4864),
.B(n_4751),
.Y(n_4913)
);

OR2x2_ASAP7_75t_L g4914 ( 
.A(n_4880),
.B(n_4836),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4855),
.B(n_4843),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_L g4916 ( 
.A(n_4884),
.B(n_4892),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4888),
.Y(n_4917)
);

NOR2x1_ASAP7_75t_L g4918 ( 
.A(n_4850),
.B(n_4620),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4871),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4871),
.Y(n_4920)
);

AND2x2_ASAP7_75t_L g4921 ( 
.A(n_4884),
.B(n_4779),
.Y(n_4921)
);

AND2x2_ASAP7_75t_L g4922 ( 
.A(n_4867),
.B(n_4872),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4890),
.Y(n_4923)
);

AND2x2_ASAP7_75t_L g4924 ( 
.A(n_4867),
.B(n_4663),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4849),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4890),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4890),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_4892),
.B(n_4797),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4872),
.B(n_4873),
.Y(n_4929)
);

BUFx2_ASAP7_75t_L g4930 ( 
.A(n_4849),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4847),
.Y(n_4931)
);

AND2x4_ASAP7_75t_L g4932 ( 
.A(n_4849),
.B(n_4798),
.Y(n_4932)
);

AND2x4_ASAP7_75t_L g4933 ( 
.A(n_4849),
.B(n_4870),
.Y(n_4933)
);

INVx3_ASAP7_75t_L g4934 ( 
.A(n_4870),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4930),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4922),
.B(n_4915),
.Y(n_4936)
);

OR2x2_ASAP7_75t_L g4937 ( 
.A(n_4896),
.B(n_4860),
.Y(n_4937)
);

INVx1_ASAP7_75t_SL g4938 ( 
.A(n_4924),
.Y(n_4938)
);

OR2x2_ASAP7_75t_L g4939 ( 
.A(n_4916),
.B(n_4862),
.Y(n_4939)
);

INVx2_ASAP7_75t_L g4940 ( 
.A(n_4896),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4929),
.B(n_4877),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4910),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4932),
.B(n_4877),
.Y(n_4943)
);

OR2x2_ASAP7_75t_L g4944 ( 
.A(n_4916),
.B(n_4734),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4910),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4910),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4910),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4898),
.B(n_4881),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4934),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4934),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4933),
.Y(n_4951)
);

OR2x2_ASAP7_75t_L g4952 ( 
.A(n_4907),
.B(n_4734),
.Y(n_4952)
);

OR2x6_ASAP7_75t_L g4953 ( 
.A(n_4905),
.B(n_4911),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4933),
.B(n_4881),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4933),
.Y(n_4955)
);

OR2x2_ASAP7_75t_L g4956 ( 
.A(n_4907),
.B(n_4742),
.Y(n_4956)
);

OR2x2_ASAP7_75t_L g4957 ( 
.A(n_4913),
.B(n_4837),
.Y(n_4957)
);

INVx2_ASAP7_75t_L g4958 ( 
.A(n_4901),
.Y(n_4958)
);

AND2x2_ASAP7_75t_L g4959 ( 
.A(n_4921),
.B(n_4847),
.Y(n_4959)
);

INVxp67_ASAP7_75t_L g4960 ( 
.A(n_4899),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4900),
.B(n_4853),
.Y(n_4961)
);

AND2x2_ASAP7_75t_L g4962 ( 
.A(n_4901),
.B(n_4853),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4925),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4931),
.B(n_4857),
.Y(n_4964)
);

INVx3_ASAP7_75t_L g4965 ( 
.A(n_4932),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4925),
.Y(n_4966)
);

NAND2x1p5_ASAP7_75t_L g4967 ( 
.A(n_4917),
.B(n_4860),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4912),
.B(n_4857),
.Y(n_4968)
);

AND2x2_ASAP7_75t_L g4969 ( 
.A(n_4897),
.B(n_4859),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4919),
.B(n_4859),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4969),
.B(n_4875),
.Y(n_4971)
);

OAI22xp5_ASAP7_75t_L g4972 ( 
.A1(n_4967),
.A2(n_4885),
.B1(n_4620),
.B2(n_4909),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4965),
.Y(n_4973)
);

AOI211x1_ASAP7_75t_SL g4974 ( 
.A1(n_4943),
.A2(n_4909),
.B(n_4833),
.C(n_4839),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4965),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4965),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4937),
.Y(n_4977)
);

OR2x2_ASAP7_75t_L g4978 ( 
.A(n_4952),
.B(n_4928),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4969),
.B(n_4875),
.Y(n_4979)
);

INVxp67_ASAP7_75t_L g4980 ( 
.A(n_4948),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4948),
.B(n_4863),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4937),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4967),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4962),
.Y(n_4984)
);

OR2x2_ASAP7_75t_L g4985 ( 
.A(n_4956),
.B(n_4928),
.Y(n_4985)
);

HB1xp67_ASAP7_75t_L g4986 ( 
.A(n_4962),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4954),
.B(n_4961),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4954),
.B(n_4863),
.Y(n_4988)
);

AOI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4938),
.A2(n_4713),
.B1(n_4620),
.B2(n_4918),
.Y(n_4989)
);

INVx1_ASAP7_75t_SL g4990 ( 
.A(n_4959),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4951),
.Y(n_4991)
);

INVx2_ASAP7_75t_SL g4992 ( 
.A(n_4955),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4961),
.Y(n_4993)
);

INVx1_ASAP7_75t_SL g4994 ( 
.A(n_4959),
.Y(n_4994)
);

AND2x2_ASAP7_75t_L g4995 ( 
.A(n_4941),
.B(n_4887),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4941),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4958),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4958),
.Y(n_4998)
);

AOI322xp5_ASAP7_75t_L g4999 ( 
.A1(n_4936),
.A2(n_4808),
.A3(n_4908),
.B1(n_4727),
.B2(n_4701),
.C1(n_4725),
.C2(n_4752),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4971),
.B(n_4968),
.Y(n_5000)
);

OAI33xp33_ASAP7_75t_L g5001 ( 
.A1(n_4972),
.A2(n_4908),
.A3(n_4935),
.B1(n_4852),
.B2(n_4851),
.B3(n_4848),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4979),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4995),
.B(n_4968),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4996),
.B(n_4970),
.Y(n_5004)
);

INVxp67_ASAP7_75t_SL g5005 ( 
.A(n_4981),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4986),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4988),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4987),
.Y(n_5008)
);

HB1xp67_ASAP7_75t_L g5009 ( 
.A(n_4972),
.Y(n_5009)
);

BUFx2_ASAP7_75t_L g5010 ( 
.A(n_4983),
.Y(n_5010)
);

AND2x2_ASAP7_75t_L g5011 ( 
.A(n_4990),
.B(n_4970),
.Y(n_5011)
);

OAI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4999),
.A2(n_4808),
.B(n_4960),
.Y(n_5012)
);

OR2x2_ASAP7_75t_L g5013 ( 
.A(n_4990),
.B(n_4944),
.Y(n_5013)
);

NAND2x1p5_ASAP7_75t_L g5014 ( 
.A(n_4994),
.B(n_4949),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4977),
.Y(n_5015)
);

AOI32xp33_ASAP7_75t_L g5016 ( 
.A1(n_4994),
.A2(n_4691),
.A3(n_4790),
.B1(n_4887),
.B2(n_4889),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4987),
.Y(n_5017)
);

AND2x2_ASAP7_75t_L g5018 ( 
.A(n_4993),
.B(n_4889),
.Y(n_5018)
);

NOR2xp33_ASAP7_75t_L g5019 ( 
.A(n_4980),
.B(n_4801),
.Y(n_5019)
);

AND2x4_ASAP7_75t_L g5020 ( 
.A(n_4982),
.B(n_4870),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_5020),
.B(n_4964),
.Y(n_5021)
);

OA21x2_ASAP7_75t_L g5022 ( 
.A1(n_5012),
.A2(n_4926),
.B(n_4923),
.Y(n_5022)
);

INVxp67_ASAP7_75t_L g5023 ( 
.A(n_5020),
.Y(n_5023)
);

AOI22xp5_ASAP7_75t_L g5024 ( 
.A1(n_5002),
.A2(n_4765),
.B1(n_4992),
.B2(n_4825),
.Y(n_5024)
);

AOI21xp33_ASAP7_75t_L g5025 ( 
.A1(n_5013),
.A2(n_4906),
.B(n_4978),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_5014),
.Y(n_5026)
);

HB1xp67_ASAP7_75t_L g5027 ( 
.A(n_5014),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_5003),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_5000),
.B(n_4964),
.Y(n_5029)
);

AOI21xp33_ASAP7_75t_L g5030 ( 
.A1(n_5011),
.A2(n_4985),
.B(n_4904),
.Y(n_5030)
);

INVxp67_ASAP7_75t_L g5031 ( 
.A(n_5004),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_5018),
.Y(n_5032)
);

AOI22xp5_ASAP7_75t_L g5033 ( 
.A1(n_5019),
.A2(n_4903),
.B1(n_4902),
.B2(n_4840),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_5010),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_5001),
.B(n_4939),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_5006),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_5015),
.B(n_4834),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_5029),
.B(n_4920),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_5027),
.Y(n_5039)
);

AND2x2_ASAP7_75t_L g5040 ( 
.A(n_5023),
.B(n_4984),
.Y(n_5040)
);

OAI22xp5_ASAP7_75t_L g5041 ( 
.A1(n_5024),
.A2(n_4989),
.B1(n_4627),
.B2(n_4957),
.Y(n_5041)
);

OAI32xp33_ASAP7_75t_L g5042 ( 
.A1(n_5026),
.A2(n_4974),
.A3(n_4891),
.B1(n_5009),
.B2(n_4991),
.Y(n_5042)
);

AOI22xp5_ASAP7_75t_L g5043 ( 
.A1(n_5028),
.A2(n_4786),
.B1(n_4780),
.B2(n_4870),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_5021),
.Y(n_5044)
);

AOI22xp5_ASAP7_75t_L g5045 ( 
.A1(n_5034),
.A2(n_5007),
.B1(n_4950),
.B2(n_5008),
.Y(n_5045)
);

NOR2xp33_ASAP7_75t_L g5046 ( 
.A(n_5031),
.B(n_5001),
.Y(n_5046)
);

AOI21xp5_ASAP7_75t_L g5047 ( 
.A1(n_5025),
.A2(n_5005),
.B(n_5012),
.Y(n_5047)
);

OAI311xp33_ASAP7_75t_L g5048 ( 
.A1(n_5033),
.A2(n_4891),
.A3(n_5016),
.B1(n_4914),
.C1(n_4886),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_5035),
.B(n_4973),
.Y(n_5049)
);

OAI21x1_ASAP7_75t_SL g5050 ( 
.A1(n_5022),
.A2(n_4868),
.B(n_4946),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_5022),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_5037),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_5032),
.B(n_4975),
.Y(n_5053)
);

OAI22xp5_ASAP7_75t_L g5054 ( 
.A1(n_5036),
.A2(n_4627),
.B1(n_4756),
.B2(n_4761),
.Y(n_5054)
);

OAI21xp5_ASAP7_75t_L g5055 ( 
.A1(n_5030),
.A2(n_5005),
.B(n_5009),
.Y(n_5055)
);

AOI31xp33_ASAP7_75t_L g5056 ( 
.A1(n_5023),
.A2(n_4976),
.A3(n_4942),
.B(n_4945),
.Y(n_5056)
);

NAND2xp33_ASAP7_75t_SL g5057 ( 
.A(n_5027),
.B(n_4868),
.Y(n_5057)
);

OR2x2_ASAP7_75t_L g5058 ( 
.A(n_5038),
.B(n_4953),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_5050),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_5040),
.Y(n_5060)
);

NOR2xp33_ASAP7_75t_L g5061 ( 
.A(n_5056),
.B(n_5017),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5043),
.B(n_4868),
.Y(n_5062)
);

AND2x2_ASAP7_75t_L g5063 ( 
.A(n_5055),
.B(n_4953),
.Y(n_5063)
);

AOI22xp5_ASAP7_75t_SL g5064 ( 
.A1(n_5041),
.A2(n_4966),
.B1(n_4963),
.B2(n_4851),
.Y(n_5064)
);

AOI322xp5_ASAP7_75t_L g5065 ( 
.A1(n_5046),
.A2(n_4997),
.A3(n_4883),
.B1(n_4848),
.B2(n_4852),
.C1(n_4998),
.C2(n_4894),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_5039),
.B(n_4883),
.Y(n_5066)
);

OAI22xp33_ASAP7_75t_SL g5067 ( 
.A1(n_5049),
.A2(n_4886),
.B1(n_4953),
.B2(n_4878),
.Y(n_5067)
);

AOI22xp33_ASAP7_75t_L g5068 ( 
.A1(n_5044),
.A2(n_4722),
.B1(n_4743),
.B2(n_4713),
.Y(n_5068)
);

AND2x2_ASAP7_75t_L g5069 ( 
.A(n_5052),
.B(n_4953),
.Y(n_5069)
);

AOI22xp5_ASAP7_75t_L g5070 ( 
.A1(n_5057),
.A2(n_4841),
.B1(n_4844),
.B2(n_4764),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_5054),
.B(n_4946),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_5051),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_5047),
.B(n_4947),
.Y(n_5073)
);

NOR2xp33_ASAP7_75t_L g5074 ( 
.A(n_5042),
.B(n_4947),
.Y(n_5074)
);

OAI22xp33_ASAP7_75t_SL g5075 ( 
.A1(n_5053),
.A2(n_4878),
.B1(n_4927),
.B2(n_4894),
.Y(n_5075)
);

AOI221x1_ASAP7_75t_SL g5076 ( 
.A1(n_5048),
.A2(n_4879),
.B1(n_4869),
.B2(n_4865),
.C(n_4940),
.Y(n_5076)
);

AOI221xp5_ASAP7_75t_L g5077 ( 
.A1(n_5045),
.A2(n_4879),
.B1(n_4865),
.B2(n_4869),
.C(n_4793),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_5043),
.B(n_4874),
.Y(n_5078)
);

AOI22xp5_ASAP7_75t_L g5079 ( 
.A1(n_5040),
.A2(n_4764),
.B1(n_4823),
.B2(n_4821),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_5050),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_5050),
.Y(n_5081)
);

INVxp67_ASAP7_75t_L g5082 ( 
.A(n_5057),
.Y(n_5082)
);

NAND2xp33_ASAP7_75t_SL g5083 ( 
.A(n_5038),
.B(n_4940),
.Y(n_5083)
);

AOI22xp5_ASAP7_75t_L g5084 ( 
.A1(n_5040),
.A2(n_4764),
.B1(n_4827),
.B2(n_4826),
.Y(n_5084)
);

NAND2x1_ASAP7_75t_L g5085 ( 
.A(n_5050),
.B(n_4874),
.Y(n_5085)
);

AOI211x1_ASAP7_75t_SL g5086 ( 
.A1(n_5054),
.A2(n_4882),
.B(n_4876),
.C(n_4874),
.Y(n_5086)
);

AOI21xp5_ASAP7_75t_L g5087 ( 
.A1(n_5057),
.A2(n_4882),
.B(n_4876),
.Y(n_5087)
);

AND2x2_ASAP7_75t_L g5088 ( 
.A(n_5069),
.B(n_4876),
.Y(n_5088)
);

AOI221xp5_ASAP7_75t_L g5089 ( 
.A1(n_5067),
.A2(n_4793),
.B1(n_4795),
.B2(n_4882),
.C(n_4815),
.Y(n_5089)
);

AOI222xp33_ASAP7_75t_L g5090 ( 
.A1(n_5077),
.A2(n_5082),
.B1(n_4782),
.B2(n_4783),
.C1(n_4768),
.C2(n_4795),
.Y(n_5090)
);

AOI222xp33_ASAP7_75t_L g5091 ( 
.A1(n_5083),
.A2(n_4783),
.B1(n_4782),
.B2(n_4768),
.C1(n_4757),
.C2(n_4744),
.Y(n_5091)
);

OAI22xp33_ASAP7_75t_L g5092 ( 
.A1(n_5070),
.A2(n_4691),
.B1(n_4810),
.B2(n_4804),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_5085),
.Y(n_5093)
);

AOI22xp33_ASAP7_75t_L g5094 ( 
.A1(n_5063),
.A2(n_5060),
.B1(n_5061),
.B2(n_5074),
.Y(n_5094)
);

AOI222xp33_ASAP7_75t_L g5095 ( 
.A1(n_5072),
.A2(n_4744),
.B1(n_4757),
.B2(n_4759),
.C1(n_4758),
.C2(n_4814),
.Y(n_5095)
);

AOI211xp5_ASAP7_75t_L g5096 ( 
.A1(n_5075),
.A2(n_4810),
.B(n_4804),
.C(n_4796),
.Y(n_5096)
);

OAI32xp33_ASAP7_75t_L g5097 ( 
.A1(n_5086),
.A2(n_4796),
.A3(n_4759),
.B1(n_4758),
.B2(n_4772),
.Y(n_5097)
);

AND2x4_ASAP7_75t_L g5098 ( 
.A(n_5079),
.B(n_5084),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_5065),
.B(n_4769),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_5062),
.Y(n_5100)
);

OAI22xp5_ASAP7_75t_L g5101 ( 
.A1(n_5058),
.A2(n_4687),
.B1(n_4743),
.B2(n_4769),
.Y(n_5101)
);

AOI21xp5_ASAP7_75t_L g5102 ( 
.A1(n_5087),
.A2(n_5073),
.B(n_5078),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5064),
.Y(n_5103)
);

OAI221xp5_ASAP7_75t_L g5104 ( 
.A1(n_5076),
.A2(n_4771),
.B1(n_4772),
.B2(n_4777),
.C(n_4697),
.Y(n_5104)
);

OAI211xp5_ASAP7_75t_L g5105 ( 
.A1(n_5068),
.A2(n_4771),
.B(n_4777),
.C(n_4789),
.Y(n_5105)
);

AOI211xp5_ASAP7_75t_L g5106 ( 
.A1(n_5066),
.A2(n_5071),
.B(n_5080),
.C(n_5081),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_SL g5107 ( 
.A(n_5059),
.B(n_4743),
.Y(n_5107)
);

OAI211xp5_ASAP7_75t_SL g5108 ( 
.A1(n_5065),
.A2(n_4701),
.B(n_4787),
.C(n_4789),
.Y(n_5108)
);

INVxp67_ASAP7_75t_L g5109 ( 
.A(n_5062),
.Y(n_5109)
);

NOR2xp33_ASAP7_75t_SL g5110 ( 
.A(n_5069),
.B(n_4710),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5085),
.Y(n_5111)
);

AOI21xp5_ASAP7_75t_L g5112 ( 
.A1(n_5085),
.A2(n_4656),
.B(n_4774),
.Y(n_5112)
);

OAI21xp5_ASAP7_75t_SL g5113 ( 
.A1(n_5079),
.A2(n_4774),
.B(n_4784),
.Y(n_5113)
);

INVx1_ASAP7_75t_SL g5114 ( 
.A(n_5069),
.Y(n_5114)
);

AOI221xp5_ASAP7_75t_L g5115 ( 
.A1(n_5067),
.A2(n_4691),
.B1(n_4784),
.B2(n_4676),
.C(n_4667),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5070),
.B(n_4595),
.Y(n_5116)
);

OA211x2_ASAP7_75t_L g5117 ( 
.A1(n_5074),
.A2(n_4655),
.B(n_4493),
.C(n_4560),
.Y(n_5117)
);

OAI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_5061),
.A2(n_4702),
.B(n_4700),
.Y(n_5118)
);

AOI221xp5_ASAP7_75t_L g5119 ( 
.A1(n_5101),
.A2(n_4667),
.B1(n_4787),
.B2(n_4716),
.C(n_4676),
.Y(n_5119)
);

NAND3xp33_ASAP7_75t_SL g5120 ( 
.A(n_5096),
.B(n_4529),
.C(n_4688),
.Y(n_5120)
);

AOI211xp5_ASAP7_75t_L g5121 ( 
.A1(n_5092),
.A2(n_4681),
.B(n_4700),
.C(n_4702),
.Y(n_5121)
);

AOI22xp5_ASAP7_75t_L g5122 ( 
.A1(n_5110),
.A2(n_4681),
.B1(n_4705),
.B2(n_4710),
.Y(n_5122)
);

AOI21xp33_ASAP7_75t_L g5123 ( 
.A1(n_5114),
.A2(n_4579),
.B(n_4529),
.Y(n_5123)
);

AOI211xp5_ASAP7_75t_L g5124 ( 
.A1(n_5097),
.A2(n_4681),
.B(n_4705),
.C(n_4716),
.Y(n_5124)
);

AND3x1_ASAP7_75t_L g5125 ( 
.A(n_5088),
.B(n_4693),
.C(n_4688),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_5099),
.Y(n_5126)
);

AOI221xp5_ASAP7_75t_L g5127 ( 
.A1(n_5115),
.A2(n_4681),
.B1(n_4704),
.B2(n_4694),
.C(n_4714),
.Y(n_5127)
);

OA211x2_ASAP7_75t_L g5128 ( 
.A1(n_5107),
.A2(n_5089),
.B(n_5116),
.C(n_5109),
.Y(n_5128)
);

AOI211xp5_ASAP7_75t_SL g5129 ( 
.A1(n_5103),
.A2(n_4693),
.B(n_4696),
.C(n_4525),
.Y(n_5129)
);

INVx2_ASAP7_75t_SL g5130 ( 
.A(n_5098),
.Y(n_5130)
);

NOR3xp33_ASAP7_75t_L g5131 ( 
.A(n_5100),
.B(n_5106),
.C(n_5102),
.Y(n_5131)
);

AOI21xp5_ASAP7_75t_L g5132 ( 
.A1(n_5112),
.A2(n_4531),
.B(n_4587),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5118),
.Y(n_5133)
);

NOR4xp25_ASAP7_75t_L g5134 ( 
.A(n_5094),
.B(n_4637),
.C(n_4628),
.D(n_4694),
.Y(n_5134)
);

AOI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_5093),
.A2(n_4584),
.B(n_4699),
.Y(n_5135)
);

AOI222xp33_ASAP7_75t_L g5136 ( 
.A1(n_5108),
.A2(n_4559),
.B1(n_4696),
.B2(n_4704),
.C1(n_4714),
.C2(n_4699),
.Y(n_5136)
);

NOR2x1_ASAP7_75t_L g5137 ( 
.A(n_5111),
.B(n_5098),
.Y(n_5137)
);

AOI322xp5_ASAP7_75t_L g5138 ( 
.A1(n_5117),
.A2(n_4588),
.A3(n_4501),
.B1(n_4610),
.B2(n_4679),
.C1(n_4608),
.C2(n_4638),
.Y(n_5138)
);

NAND4xp25_ASAP7_75t_L g5139 ( 
.A(n_5090),
.B(n_4664),
.C(n_4660),
.D(n_4633),
.Y(n_5139)
);

OAI21xp5_ASAP7_75t_SL g5140 ( 
.A1(n_5113),
.A2(n_4709),
.B(n_4707),
.Y(n_5140)
);

OAI322xp33_ASAP7_75t_L g5141 ( 
.A1(n_5104),
.A2(n_4664),
.A3(n_4637),
.B1(n_4628),
.B2(n_4708),
.C1(n_4660),
.C2(n_4659),
.Y(n_5141)
);

OAI211xp5_ASAP7_75t_SL g5142 ( 
.A1(n_5091),
.A2(n_4526),
.B(n_4590),
.C(n_4708),
.Y(n_5142)
);

AOI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_5105),
.A2(n_4649),
.B(n_4647),
.Y(n_5143)
);

NOR2xp67_ASAP7_75t_L g5144 ( 
.A(n_5095),
.B(n_4707),
.Y(n_5144)
);

AOI221xp5_ASAP7_75t_L g5145 ( 
.A1(n_5101),
.A2(n_4649),
.B1(n_4647),
.B2(n_4659),
.C(n_4680),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_5088),
.Y(n_5146)
);

NAND3xp33_ASAP7_75t_SL g5147 ( 
.A(n_5096),
.B(n_4709),
.C(n_4633),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_5122),
.B(n_4723),
.Y(n_5148)
);

A2O1A1Ixp33_ASAP7_75t_L g5149 ( 
.A1(n_5119),
.A2(n_5144),
.B(n_5130),
.C(n_5132),
.Y(n_5149)
);

AOI221x1_ASAP7_75t_L g5150 ( 
.A1(n_5131),
.A2(n_5126),
.B1(n_5146),
.B2(n_5133),
.C(n_5123),
.Y(n_5150)
);

NAND3xp33_ASAP7_75t_L g5151 ( 
.A(n_5137),
.B(n_4680),
.C(n_4685),
.Y(n_5151)
);

A2O1A1Ixp33_ASAP7_75t_L g5152 ( 
.A1(n_5143),
.A2(n_4684),
.B(n_4685),
.C(n_4717),
.Y(n_5152)
);

OAI211xp5_ASAP7_75t_L g5153 ( 
.A1(n_5134),
.A2(n_5124),
.B(n_5135),
.C(n_5139),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_5138),
.B(n_4723),
.Y(n_5154)
);

O2A1O1Ixp33_ASAP7_75t_L g5155 ( 
.A1(n_5120),
.A2(n_4684),
.B(n_4602),
.C(n_4717),
.Y(n_5155)
);

OAI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_5147),
.A2(n_4672),
.B(n_4668),
.Y(n_5156)
);

AOI21xp5_ASAP7_75t_L g5157 ( 
.A1(n_5125),
.A2(n_4663),
.B(n_4672),
.Y(n_5157)
);

NOR3xp33_ASAP7_75t_L g5158 ( 
.A(n_5142),
.B(n_4499),
.C(n_4590),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_5121),
.B(n_4636),
.Y(n_5159)
);

INVx2_ASAP7_75t_L g5160 ( 
.A(n_5128),
.Y(n_5160)
);

NAND3xp33_ASAP7_75t_L g5161 ( 
.A(n_5127),
.B(n_4719),
.C(n_4625),
.Y(n_5161)
);

AOI322xp5_ASAP7_75t_L g5162 ( 
.A1(n_5145),
.A2(n_4679),
.A3(n_4586),
.B1(n_4592),
.B2(n_4591),
.C1(n_4602),
.C2(n_4598),
.Y(n_5162)
);

INVx2_ASAP7_75t_L g5163 ( 
.A(n_5140),
.Y(n_5163)
);

AOI221xp5_ASAP7_75t_L g5164 ( 
.A1(n_5141),
.A2(n_4719),
.B1(n_4668),
.B2(n_4636),
.C(n_4653),
.Y(n_5164)
);

AOI221xp5_ASAP7_75t_L g5165 ( 
.A1(n_5136),
.A2(n_4668),
.B1(n_4636),
.B2(n_4653),
.C(n_4629),
.Y(n_5165)
);

O2A1O1Ixp5_ASAP7_75t_SL g5166 ( 
.A1(n_5129),
.A2(n_4522),
.B(n_4547),
.C(n_4557),
.Y(n_5166)
);

AOI221xp5_ASAP7_75t_L g5167 ( 
.A1(n_5123),
.A2(n_4668),
.B1(n_4636),
.B2(n_4653),
.C(n_4626),
.Y(n_5167)
);

AOI211xp5_ASAP7_75t_L g5168 ( 
.A1(n_5123),
.A2(n_4625),
.B(n_4626),
.C(n_4629),
.Y(n_5168)
);

NOR2xp33_ASAP7_75t_L g5169 ( 
.A(n_5139),
.B(n_4645),
.Y(n_5169)
);

NAND3xp33_ASAP7_75t_SL g5170 ( 
.A(n_5153),
.B(n_5149),
.C(n_5166),
.Y(n_5170)
);

NOR2x1_ASAP7_75t_SL g5171 ( 
.A(n_5151),
.B(n_4539),
.Y(n_5171)
);

NOR2x1_ASAP7_75t_L g5172 ( 
.A(n_5160),
.B(n_5163),
.Y(n_5172)
);

NAND4xp75_ASAP7_75t_L g5173 ( 
.A(n_5150),
.B(n_4645),
.C(n_4650),
.D(n_4678),
.Y(n_5173)
);

NOR3xp33_ASAP7_75t_L g5174 ( 
.A(n_5169),
.B(n_4497),
.C(n_4678),
.Y(n_5174)
);

NAND3xp33_ASAP7_75t_L g5175 ( 
.A(n_5159),
.B(n_4532),
.C(n_4650),
.Y(n_5175)
);

NOR2xp33_ASAP7_75t_L g5176 ( 
.A(n_5161),
.B(n_4653),
.Y(n_5176)
);

AOI221xp5_ASAP7_75t_L g5177 ( 
.A1(n_5157),
.A2(n_4554),
.B1(n_4594),
.B2(n_4596),
.C(n_4586),
.Y(n_5177)
);

AOI211xp5_ASAP7_75t_L g5178 ( 
.A1(n_5156),
.A2(n_4532),
.B(n_4554),
.C(n_4548),
.Y(n_5178)
);

NOR2xp33_ASAP7_75t_L g5179 ( 
.A(n_5154),
.B(n_4586),
.Y(n_5179)
);

AND2x2_ASAP7_75t_L g5180 ( 
.A(n_5168),
.B(n_4582),
.Y(n_5180)
);

OAI221xp5_ASAP7_75t_SL g5181 ( 
.A1(n_5164),
.A2(n_4553),
.B1(n_4567),
.B2(n_4548),
.C(n_4563),
.Y(n_5181)
);

NAND3xp33_ASAP7_75t_SL g5182 ( 
.A(n_5167),
.B(n_4546),
.C(n_4577),
.Y(n_5182)
);

AOI221xp5_ASAP7_75t_L g5183 ( 
.A1(n_5155),
.A2(n_4546),
.B1(n_4568),
.B2(n_4563),
.C(n_4569),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_5165),
.B(n_4723),
.Y(n_5184)
);

NAND3xp33_ASAP7_75t_SL g5185 ( 
.A(n_5158),
.B(n_4577),
.C(n_4572),
.Y(n_5185)
);

AOI221xp5_ASAP7_75t_L g5186 ( 
.A1(n_5181),
.A2(n_5148),
.B1(n_5152),
.B2(n_5162),
.C(n_4569),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_5170),
.A2(n_4516),
.B(n_4539),
.Y(n_5187)
);

NOR4xp25_ASAP7_75t_L g5188 ( 
.A(n_5175),
.B(n_4557),
.C(n_4550),
.D(n_4558),
.Y(n_5188)
);

NAND4xp25_ASAP7_75t_L g5189 ( 
.A(n_5179),
.B(n_5176),
.C(n_5172),
.D(n_5180),
.Y(n_5189)
);

OAI221xp5_ASAP7_75t_L g5190 ( 
.A1(n_5174),
.A2(n_4516),
.B1(n_4711),
.B2(n_4485),
.C(n_4557),
.Y(n_5190)
);

AND4x1_ASAP7_75t_L g5191 ( 
.A(n_5178),
.B(n_5177),
.C(n_5184),
.D(n_5183),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_5173),
.B(n_5171),
.Y(n_5192)
);

NAND3xp33_ASAP7_75t_L g5193 ( 
.A(n_5185),
.B(n_4516),
.C(n_4498),
.Y(n_5193)
);

OAI21xp33_ASAP7_75t_SL g5194 ( 
.A1(n_5182),
.A2(n_4572),
.B(n_4570),
.Y(n_5194)
);

NOR3xp33_ASAP7_75t_L g5195 ( 
.A(n_5170),
.B(n_4575),
.C(n_4599),
.Y(n_5195)
);

NOR2x1_ASAP7_75t_L g5196 ( 
.A(n_5170),
.B(n_4539),
.Y(n_5196)
);

NOR2x1_ASAP7_75t_L g5197 ( 
.A(n_5170),
.B(n_4484),
.Y(n_5197)
);

AOI21xp33_ASAP7_75t_SL g5198 ( 
.A1(n_5176),
.A2(n_643),
.B(n_644),
.Y(n_5198)
);

NAND4xp25_ASAP7_75t_L g5199 ( 
.A(n_5179),
.B(n_4611),
.C(n_4612),
.D(n_4570),
.Y(n_5199)
);

NAND3xp33_ASAP7_75t_L g5200 ( 
.A(n_5172),
.B(n_4498),
.C(n_4711),
.Y(n_5200)
);

AOI21x1_ASAP7_75t_L g5201 ( 
.A1(n_5172),
.A2(n_4498),
.B(n_4544),
.Y(n_5201)
);

NAND3xp33_ASAP7_75t_SL g5202 ( 
.A(n_5176),
.B(n_4611),
.C(n_4544),
.Y(n_5202)
);

NAND3xp33_ASAP7_75t_L g5203 ( 
.A(n_5172),
.B(n_4711),
.C(n_4485),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_SL g5204 ( 
.A(n_5175),
.B(n_4488),
.Y(n_5204)
);

AOI22xp5_ASAP7_75t_L g5205 ( 
.A1(n_5195),
.A2(n_4484),
.B1(n_4566),
.B2(n_4509),
.Y(n_5205)
);

NOR2xp33_ASAP7_75t_L g5206 ( 
.A(n_5202),
.B(n_4566),
.Y(n_5206)
);

OAI22xp5_ASAP7_75t_L g5207 ( 
.A1(n_5200),
.A2(n_5203),
.B1(n_5190),
.B2(n_5193),
.Y(n_5207)
);

INVx2_ASAP7_75t_L g5208 ( 
.A(n_5201),
.Y(n_5208)
);

BUFx10_ASAP7_75t_L g5209 ( 
.A(n_5189),
.Y(n_5209)
);

NOR2x1_ASAP7_75t_L g5210 ( 
.A(n_5192),
.B(n_4484),
.Y(n_5210)
);

NOR2xp67_ASAP7_75t_L g5211 ( 
.A(n_5198),
.B(n_646),
.Y(n_5211)
);

XNOR2xp5_ASAP7_75t_L g5212 ( 
.A(n_5191),
.B(n_646),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5197),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_5204),
.B(n_4723),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_5196),
.Y(n_5215)
);

AND2x2_ASAP7_75t_L g5216 ( 
.A(n_5194),
.B(n_4723),
.Y(n_5216)
);

AOI22xp5_ASAP7_75t_L g5217 ( 
.A1(n_5186),
.A2(n_4711),
.B1(n_4580),
.B2(n_4583),
.Y(n_5217)
);

AOI22xp5_ASAP7_75t_L g5218 ( 
.A1(n_5199),
.A2(n_4580),
.B1(n_4583),
.B2(n_4609),
.Y(n_5218)
);

AOI22xp5_ASAP7_75t_L g5219 ( 
.A1(n_5187),
.A2(n_4580),
.B1(n_4583),
.B2(n_4573),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5188),
.Y(n_5220)
);

NOR2x1_ASAP7_75t_L g5221 ( 
.A(n_5189),
.B(n_4573),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_5197),
.Y(n_5222)
);

NOR3xp33_ASAP7_75t_L g5223 ( 
.A(n_5220),
.B(n_4612),
.C(n_648),
.Y(n_5223)
);

AOI211xp5_ASAP7_75t_L g5224 ( 
.A1(n_5207),
.A2(n_647),
.B(n_648),
.C(n_649),
.Y(n_5224)
);

NOR3xp33_ASAP7_75t_L g5225 ( 
.A(n_5215),
.B(n_647),
.C(n_649),
.Y(n_5225)
);

NOR3xp33_ASAP7_75t_L g5226 ( 
.A(n_5213),
.B(n_650),
.C(n_651),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_5206),
.B(n_5216),
.Y(n_5227)
);

NAND4xp25_ASAP7_75t_L g5228 ( 
.A(n_5211),
.B(n_651),
.C(n_652),
.D(n_653),
.Y(n_5228)
);

NOR2x1_ASAP7_75t_L g5229 ( 
.A(n_5208),
.B(n_4573),
.Y(n_5229)
);

OR2x2_ASAP7_75t_L g5230 ( 
.A(n_5214),
.B(n_4541),
.Y(n_5230)
);

OR2x2_ASAP7_75t_L g5231 ( 
.A(n_5205),
.B(n_5212),
.Y(n_5231)
);

NOR3xp33_ASAP7_75t_L g5232 ( 
.A(n_5222),
.B(n_652),
.C(n_654),
.Y(n_5232)
);

O2A1O1Ixp5_ASAP7_75t_SL g5233 ( 
.A1(n_5209),
.A2(n_654),
.B(n_655),
.C(n_656),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_5210),
.B(n_4603),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_5224),
.B(n_5217),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5228),
.Y(n_5236)
);

OR2x2_ASAP7_75t_L g5237 ( 
.A(n_5234),
.B(n_5219),
.Y(n_5237)
);

NOR2x1_ASAP7_75t_L g5238 ( 
.A(n_5227),
.B(n_5221),
.Y(n_5238)
);

NOR2x1_ASAP7_75t_L g5239 ( 
.A(n_5231),
.B(n_5218),
.Y(n_5239)
);

AND2x2_ASAP7_75t_L g5240 ( 
.A(n_5225),
.B(n_4492),
.Y(n_5240)
);

OAI22xp5_ASAP7_75t_L g5241 ( 
.A1(n_5226),
.A2(n_4492),
.B1(n_4488),
.B2(n_4485),
.Y(n_5241)
);

NAND4xp25_ASAP7_75t_L g5242 ( 
.A(n_5239),
.B(n_5232),
.C(n_5223),
.D(n_5233),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_5240),
.B(n_5229),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_5236),
.B(n_5230),
.Y(n_5244)
);

INVx3_ASAP7_75t_SL g5245 ( 
.A(n_5237),
.Y(n_5245)
);

AO22x2_ASAP7_75t_L g5246 ( 
.A1(n_5243),
.A2(n_5235),
.B1(n_5238),
.B2(n_5241),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5245),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5247),
.Y(n_5248)
);

INVx3_ASAP7_75t_SL g5249 ( 
.A(n_5248),
.Y(n_5249)
);

OAI22xp5_ASAP7_75t_L g5250 ( 
.A1(n_5249),
.A2(n_5246),
.B1(n_5244),
.B2(n_5242),
.Y(n_5250)
);

OAI22xp5_ASAP7_75t_L g5251 ( 
.A1(n_5250),
.A2(n_4485),
.B1(n_4603),
.B2(n_4606),
.Y(n_5251)
);

HB1xp67_ASAP7_75t_L g5252 ( 
.A(n_5251),
.Y(n_5252)
);

NOR2xp67_ASAP7_75t_L g5253 ( 
.A(n_5252),
.B(n_655),
.Y(n_5253)
);

AOI22xp33_ASAP7_75t_L g5254 ( 
.A1(n_5253),
.A2(n_4603),
.B1(n_4606),
.B2(n_658),
.Y(n_5254)
);

HB1xp67_ASAP7_75t_L g5255 ( 
.A(n_5254),
.Y(n_5255)
);

NAND2xp67_ASAP7_75t_SL g5256 ( 
.A(n_5255),
.B(n_656),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_5256),
.Y(n_5257)
);

OR2x6_ASAP7_75t_L g5258 ( 
.A(n_5257),
.B(n_657),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_5257),
.B(n_657),
.Y(n_5259)
);

OAI221xp5_ASAP7_75t_L g5260 ( 
.A1(n_5258),
.A2(n_658),
.B1(n_659),
.B2(n_660),
.C(n_661),
.Y(n_5260)
);

AOI22xp33_ASAP7_75t_L g5261 ( 
.A1(n_5260),
.A2(n_5259),
.B1(n_661),
.B2(n_662),
.Y(n_5261)
);

AOI211xp5_ASAP7_75t_L g5262 ( 
.A1(n_5261),
.A2(n_659),
.B(n_662),
.C(n_663),
.Y(n_5262)
);


endmodule