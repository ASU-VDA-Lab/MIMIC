module fake_jpeg_6420_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_42),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_8),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_17),
.B1(n_24),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_32),
.B1(n_39),
.B2(n_34),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_18),
.B1(n_22),
.B2(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_54),
.B1(n_60),
.B2(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_53),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_18),
.B1(n_22),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_24),
.B1(n_31),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_63),
.B1(n_32),
.B2(n_27),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_22),
.B1(n_23),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_62),
.B1(n_30),
.B2(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_38),
.B1(n_36),
.B2(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_23),
.B1(n_30),
.B2(n_25),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_21),
.B1(n_32),
.B2(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_82),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_38),
.B1(n_39),
.B2(n_25),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_84),
.B1(n_95),
.B2(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_77),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_36),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_67),
.B(n_41),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_61),
.B1(n_59),
.B2(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_36),
.B1(n_27),
.B2(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_100),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_40),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_103),
.Y(n_146)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_105),
.A2(n_40),
.B(n_35),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_49),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_94),
.B(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_67),
.B1(n_55),
.B2(n_72),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_96),
.B1(n_81),
.B2(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_51),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_118),
.Y(n_132)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_28),
.Y(n_118)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_40),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_81),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_142),
.B1(n_152),
.B2(n_109),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_98),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_106),
.B(n_104),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_134),
.B(n_140),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_123),
.B1(n_129),
.B2(n_125),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_81),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_73),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_112),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_153),
.B(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_144),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_96),
.B1(n_76),
.B2(n_88),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_83),
.B(n_80),
.C(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_85),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_35),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_95),
.B1(n_99),
.B2(n_64),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_73),
.B(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_40),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_140),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_171),
.B1(n_173),
.B2(n_187),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_164),
.B(n_177),
.CI(n_132),
.CON(n_216),
.SN(n_216)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_106),
.B1(n_112),
.B2(n_114),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_174),
.B1(n_188),
.B2(n_152),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_179),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_73),
.B1(n_121),
.B2(n_107),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_121),
.B1(n_107),
.B2(n_119),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_119),
.B1(n_64),
.B2(n_65),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_182),
.C(n_177),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_28),
.B(n_40),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_35),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_33),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_136),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_192),
.B(n_156),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_119),
.B1(n_117),
.B2(n_101),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_130),
.A2(n_64),
.B1(n_68),
.B2(n_40),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_189),
.B(n_160),
.Y(n_202)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_56),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_144),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_56),
.B(n_33),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_205),
.C(n_208),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_188),
.B1(n_162),
.B2(n_171),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_195),
.A2(n_199),
.B(n_207),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_150),
.B(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_103),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_206),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_214),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_131),
.C(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_147),
.C(n_153),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_213),
.C(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_154),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_160),
.B(n_134),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_217),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_144),
.B1(n_158),
.B2(n_136),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_191),
.B1(n_161),
.B2(n_172),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_178),
.C(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_218),
.B(n_161),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_164),
.A2(n_132),
.B(n_133),
.Y(n_217)
);

XOR2x1_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_33),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_167),
.C(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_180),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_162),
.B1(n_165),
.B2(n_163),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_243),
.B1(n_0),
.B2(n_1),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_192),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_233),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_195),
.B(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_240),
.B1(n_211),
.B2(n_199),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_166),
.C(n_185),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_213),
.C(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_241),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_56),
.A3(n_26),
.B1(n_34),
.B2(n_33),
.C1(n_145),
.C2(n_103),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_26),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_128),
.B1(n_93),
.B2(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_209),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_237),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_220),
.B1(n_194),
.B2(n_208),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_222),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_256),
.C(n_262),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_261),
.B1(n_243),
.B2(n_228),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_264),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_216),
.B1(n_196),
.B2(n_128),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_196),
.C(n_128),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_227),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_236),
.B(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_238),
.B(n_120),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_266),
.B(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_226),
.A2(n_26),
.B1(n_34),
.B2(n_93),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_120),
.C(n_33),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_9),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_26),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_244),
.B1(n_222),
.B2(n_246),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_234),
.C(n_229),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_0),
.C(n_2),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_277),
.B(n_252),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_224),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_273),
.B(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_245),
.B(n_239),
.C(n_240),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_275),
.B(n_259),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_223),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_223),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.C(n_256),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_246),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_285),
.A2(n_286),
.B(n_290),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_278),
.B1(n_275),
.B2(n_282),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_294),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_250),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_295),
.B(n_9),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_267),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_297),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_2),
.C(n_3),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_269),
.A2(n_251),
.B1(n_266),
.B2(n_262),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_250),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_276),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_299),
.B(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.C(n_308),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_2),
.C(n_3),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_9),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_12),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_2),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_3),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_13),
.B(n_16),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_287),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_312),
.A3(n_7),
.B1(n_11),
.B2(n_13),
.C1(n_15),
.C2(n_4),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_294),
.C(n_289),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_317),
.C(n_13),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_7),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_285),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_10),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_303),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_284),
.B(n_10),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_6),
.B(n_7),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_306),
.A3(n_302),
.B1(n_309),
.B2(n_301),
.C1(n_8),
.C2(n_10),
.Y(n_319)
);

AOI332xp33_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_324),
.A3(n_4),
.B1(n_5),
.B2(n_311),
.B3(n_312),
.C1(n_231),
.C2(n_111),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_4),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_11),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_319),
.B1(n_322),
.B2(n_328),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_327),
.Y(n_331)
);


endmodule