module fake_jpeg_14522_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_12),
.B1(n_9),
.B2(n_18),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_16),
.B1(n_18),
.B2(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_16),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_28),
.B1(n_8),
.B2(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_3),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_0),
.B(n_7),
.Y(n_27)
);

XNOR2x1_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_23),
.B1(n_28),
.B2(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_36),
.B(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_17),
.B1(n_11),
.B2(n_15),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_24),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_44),
.B1(n_31),
.B2(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_41),
.B(n_45),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B(n_50),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_34),
.B(n_40),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_56),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_42),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_47),
.Y(n_57)
);

AOI321xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_38),
.A3(n_40),
.B1(n_20),
.B2(n_15),
.C(n_29),
.Y(n_58)
);

AOI21x1_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_22),
.B(n_7),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_17),
.B1(n_59),
.B2(n_44),
.Y(n_61)
);


endmodule