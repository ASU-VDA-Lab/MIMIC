module fake_jpeg_10965_n_440 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_440);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_44),
.B(n_48),
.Y(n_128)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_7),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_60),
.Y(n_112)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_53),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_86),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_66),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_29),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

CKINVDCx9p33_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_13),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_83),
.Y(n_111)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_91),
.Y(n_109)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_55),
.B1(n_53),
.B2(n_73),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_16),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_97),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_99),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_49),
.A2(n_51),
.B1(n_88),
.B2(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_138),
.B1(n_150),
.B2(n_76),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_27),
.C(n_39),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_139),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_23),
.B1(n_27),
.B2(n_31),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_137),
.B1(n_62),
.B2(n_32),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_50),
.A2(n_23),
.B1(n_39),
.B2(n_37),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_30),
.B1(n_77),
.B2(n_78),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_82),
.B(n_35),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_143),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_54),
.A2(n_31),
.B1(n_41),
.B2(n_34),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_59),
.A2(n_79),
.B1(n_68),
.B2(n_72),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_37),
.C(n_34),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_54),
.B(n_25),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_46),
.B(n_25),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_8),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_65),
.A2(n_31),
.B1(n_30),
.B2(n_41),
.Y(n_150)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_85),
.B1(n_96),
.B2(n_97),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_159),
.B1(n_166),
.B2(n_180),
.Y(n_196)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_162),
.A2(n_165),
.B(n_168),
.Y(n_215)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_177),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_101),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_R g168 ( 
.A(n_112),
.B(n_8),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_181),
.B1(n_186),
.B2(n_187),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_9),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g208 ( 
.A(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_3),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_195),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_182),
.Y(n_203)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_119),
.B(n_111),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_194),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_103),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_193),
.Y(n_216)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_10),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_106),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_98),
.A2(n_10),
.B1(n_12),
.B2(n_0),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_137),
.B1(n_103),
.B2(n_130),
.Y(n_206)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_107),
.B(n_12),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_120),
.B1(n_152),
.B2(n_108),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_187),
.B1(n_105),
.B2(n_106),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_111),
.B(n_120),
.C(n_109),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_110),
.C(n_141),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_190),
.C(n_158),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_206),
.A2(n_210),
.B1(n_212),
.B2(n_225),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_140),
.B1(n_152),
.B2(n_116),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_161),
.B1(n_162),
.B2(n_124),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_130),
.A3(n_104),
.B1(n_124),
.B2(n_132),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_186),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_108),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_162),
.A2(n_132),
.B1(n_133),
.B2(n_148),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_228),
.B(n_241),
.Y(n_273)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_133),
.B1(n_148),
.B2(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_207),
.C(n_215),
.Y(n_274)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_154),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_240),
.Y(n_267)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_199),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_153),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_199),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_157),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_174),
.B1(n_188),
.B2(n_181),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_216),
.B1(n_215),
.B2(n_202),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_252),
.B(n_168),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_178),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_254),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_212),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_263),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_245),
.B1(n_228),
.B2(n_230),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_215),
.B1(n_222),
.B2(n_225),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_275),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_231),
.C(n_235),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_254),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_238),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_201),
.B1(n_203),
.B2(n_200),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_203),
.B(n_219),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_284),
.C(n_287),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_238),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_264),
.B1(n_273),
.B2(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_231),
.C(n_236),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_241),
.C(n_244),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_260),
.C(n_268),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_256),
.A2(n_253),
.B1(n_272),
.B2(n_248),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_290),
.A2(n_297),
.B1(n_299),
.B2(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_258),
.B(n_252),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_291),
.B(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_256),
.A2(n_247),
.B1(n_234),
.B2(n_240),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_266),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_298),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_269),
.B(n_267),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_301),
.A2(n_268),
.B(n_262),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_263),
.A2(n_239),
.B1(n_250),
.B2(n_246),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_263),
.A2(n_264),
.B1(n_270),
.B2(n_275),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_271),
.B1(n_263),
.B2(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_309),
.B(n_325),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_293),
.B(n_289),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_321),
.B(n_280),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_281),
.A2(n_263),
.B1(n_265),
.B2(n_273),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_317),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_315),
.B(n_323),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_277),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_322),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_289),
.B1(n_317),
.B2(n_280),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_284),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_291),
.B(n_276),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_295),
.C(n_300),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_293),
.A2(n_271),
.B(n_262),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_333),
.C(n_337),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_313),
.B(n_325),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_233),
.B1(n_251),
.B2(n_229),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_303),
.C(n_297),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_281),
.C(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_296),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_341),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_292),
.C(n_217),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_311),
.C(n_320),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_261),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_261),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_350),
.Y(n_361)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_345),
.Y(n_353)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_348),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_310),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_232),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_364),
.B(n_173),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_360),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_344),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_321),
.C(n_318),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_342),
.A2(n_319),
.B1(n_314),
.B2(n_312),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_362),
.A2(n_365),
.B1(n_336),
.B2(n_333),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_329),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_208),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_342),
.A2(n_319),
.B(n_312),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_337),
.A2(n_251),
.B1(n_242),
.B2(n_243),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_217),
.C(n_242),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_370),
.C(n_344),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_219),
.B1(n_198),
.B2(n_213),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_198),
.C(n_200),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_372),
.A2(n_376),
.B1(n_360),
.B2(n_354),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_352),
.A2(n_332),
.B1(n_330),
.B2(n_350),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_381),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_356),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_374),
.B(n_382),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_375),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_362),
.A2(n_343),
.B1(n_341),
.B2(n_339),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_367),
.Y(n_378)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_379),
.A2(n_361),
.B1(n_214),
.B2(n_221),
.Y(n_402)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_380),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_213),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_386),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_357),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_384),
.Y(n_389)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_221),
.C(n_163),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_385),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_366),
.Y(n_390)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_351),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_397),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_377),
.A2(n_368),
.B1(n_359),
.B2(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_401),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_351),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_375),
.A2(n_353),
.B1(n_364),
.B2(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_402),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_387),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_403),
.B(n_405),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_399),
.Y(n_405)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_400),
.A2(n_381),
.B(n_361),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_391),
.B(n_390),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_214),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_414),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_208),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_402),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_155),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_416),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_406),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_420),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_410),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_392),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_392),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_404),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_427),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_423),
.A2(n_404),
.B(n_397),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_429),
.C(n_227),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_422),
.B(n_105),
.Y(n_429)
);

A2O1A1O1Ixp25_ASAP7_75t_L g430 ( 
.A1(n_424),
.A2(n_415),
.B(n_419),
.C(n_417),
.D(n_227),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_432),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_425),
.A2(n_417),
.B(n_227),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_431),
.A2(n_433),
.B(n_426),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_434),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_433),
.Y(n_436)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_436),
.B(n_435),
.C(n_208),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_126),
.B(n_0),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_0),
.Y(n_440)
);


endmodule