module fake_netlist_1_3012_n_48 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_48);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_48;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
BUFx6f_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_12), .B(n_10), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_11), .B(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_7), .B(n_4), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_1), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_2), .B(n_9), .Y(n_22) );
AND2x6_ASAP7_75t_L g23 ( .A(n_0), .B(n_5), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_18), .B(n_1), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_22), .B(n_3), .Y(n_26) );
OR2x6_ASAP7_75t_L g27 ( .A(n_22), .B(n_8), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_16), .Y(n_28) );
OA21x2_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_20), .B(n_19), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_25), .Y(n_30) );
AO21x2_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_17), .B(n_23), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
INVx5_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_30), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_33), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
OAI21xp5_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_33), .B(n_29), .Y(n_39) );
OAI221xp5_ASAP7_75t_L g40 ( .A1(n_36), .A2(n_24), .B1(n_27), .B2(n_29), .C(n_16), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
OR2x2_ASAP7_75t_L g42 ( .A(n_41), .B(n_40), .Y(n_42) );
AND2x2_ASAP7_75t_L g43 ( .A(n_39), .B(n_27), .Y(n_43) );
CKINVDCx5p33_ASAP7_75t_R g44 ( .A(n_41), .Y(n_44) );
NOR2xp33_ASAP7_75t_L g45 ( .A(n_44), .B(n_31), .Y(n_45) );
AO22x2_ASAP7_75t_L g46 ( .A1(n_42), .A2(n_23), .B1(n_15), .B2(n_13), .Y(n_46) );
CKINVDCx20_ASAP7_75t_R g47 ( .A(n_45), .Y(n_47) );
AOI22xp5_ASAP7_75t_L g48 ( .A1(n_47), .A2(n_46), .B1(n_43), .B2(n_23), .Y(n_48) );
endmodule