module fake_ariane_775_n_1850 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1850);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1850;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_93),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_99),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_68),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_34),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_63),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_83),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_23),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_62),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_120),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_79),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_32),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_17),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_24),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_78),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_21),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_65),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_37),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_87),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_114),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_157),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_64),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_17),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_86),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_2),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_113),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_117),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_25),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_96),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_26),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_123),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_160),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_30),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_50),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_45),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_104),
.Y(n_252)
);

BUFx2_ASAP7_75t_SL g253 ( 
.A(n_43),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_41),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_18),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_61),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_25),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_35),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_115),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_67),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_107),
.Y(n_262)
);

INVxp33_ASAP7_75t_R g263 ( 
.A(n_50),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_175),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_30),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_44),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_106),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_58),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_69),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_77),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_48),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_135),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_178),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_20),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_40),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_35),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_148),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_34),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_26),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_49),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_100),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_75),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_176),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_85),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_172),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_45),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_47),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_163),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_112),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_37),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_151),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_56),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_47),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_149),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_18),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_13),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_137),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_16),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_82),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_146),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_2),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_46),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_42),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_109),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_110),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_36),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_10),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_132),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_153),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_105),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_28),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_126),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_31),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_169),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_9),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_24),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_170),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_20),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_7),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_84),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_128),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_1),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_11),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_31),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_10),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_74),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_91),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_119),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_179),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_1),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_141),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_70),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_111),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_138),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_101),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_40),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_0),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_33),
.Y(n_347)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_15),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_136),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_81),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_59),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_14),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_7),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_6),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_88),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_95),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_150),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_43),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_41),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_250),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_250),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_318),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_206),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_276),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_236),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_214),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_233),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_254),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_259),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_318),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_283),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_236),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_278),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_278),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_352),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_352),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_290),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_209),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_318),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_277),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_282),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_180),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_180),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_295),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_291),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_253),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_181),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_181),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_266),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_186),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_266),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_325),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_207),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_182),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_182),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_189),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_184),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_206),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_187),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_192),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_217),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_189),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_193),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_194),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_198),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_197),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_200),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_184),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_201),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_198),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_183),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_331),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_215),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_222),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_185),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_225),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_226),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_217),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_237),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_239),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_202),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_247),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_268),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_331),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_333),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_411),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_447),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_269),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_411),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_270),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_365),
.A2(n_272),
.B(n_271),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_437),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_367),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_415),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_415),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_368),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_369),
.B(n_245),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_370),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_406),
.B(n_363),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_431),
.A2(n_302),
.B1(n_315),
.B2(n_332),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_369),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_371),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_373),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_429),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_429),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_427),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_451),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_385),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_275),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_425),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_394),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_375),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_398),
.B(n_284),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_364),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_245),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_248),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_285),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_439),
.B(n_248),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_440),
.B(n_256),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_387),
.B(n_333),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_388),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_398),
.B(n_400),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_443),
.B(n_202),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_400),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_392),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_289),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_360),
.B(n_334),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_445),
.B(n_446),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_448),
.B(n_256),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_361),
.B(n_334),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_449),
.B(n_296),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_377),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_378),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_379),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_380),
.A2(n_320),
.B(n_316),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_362),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_322),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_381),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_383),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_412),
.B(n_416),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_472),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_501),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_513),
.B(n_366),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_477),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_472),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_418),
.B1(n_450),
.B2(n_438),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_521),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_469),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_469),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_500),
.B(n_216),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_474),
.B(n_493),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_513),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_474),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_477),
.B(n_351),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_470),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_500),
.B(n_501),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_475),
.A2(n_393),
.B1(n_382),
.B2(n_366),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_529),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_529),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_477),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_510),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_478),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_478),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_500),
.B(n_382),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_512),
.B(n_408),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_498),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_478),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_477),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_473),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_478),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_473),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_480),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_491),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_476),
.B(n_409),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_521),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_521),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_493),
.B(n_409),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_480),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_480),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_480),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_491),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_516),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_482),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_527),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_501),
.B(n_393),
.Y(n_589)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_463),
.A2(n_257),
.B(n_216),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_475),
.A2(n_404),
.B1(n_441),
.B2(n_419),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_453),
.A2(n_441),
.B1(n_434),
.B2(n_422),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_518),
.B(n_501),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_482),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_476),
.B(n_419),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_476),
.B(n_495),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_455),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_457),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_482),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_482),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_487),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_514),
.B(n_420),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_525),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_476),
.B(n_420),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_487),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_422),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_487),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_518),
.B(n_414),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_487),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_487),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_515),
.A2(n_434),
.B1(n_436),
.B2(n_421),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_488),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_488),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_506),
.B(n_417),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_488),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_525),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_490),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_522),
.B(n_389),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_471),
.B(n_390),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_494),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_471),
.B(n_391),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_488),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_488),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_453),
.B(n_395),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_460),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_492),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_496),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_492),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_492),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_515),
.B(n_353),
.C(n_346),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_496),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_492),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_471),
.B(n_396),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_497),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_519),
.B(n_185),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_471),
.B(n_399),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_519),
.B(n_188),
.Y(n_644)
);

AND3x2_ASAP7_75t_L g645 ( 
.A(n_458),
.B(n_263),
.C(n_403),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_503),
.B(n_188),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_503),
.B(n_190),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_525),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_486),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_511),
.B(n_351),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

AO21x2_ASAP7_75t_L g653 ( 
.A1(n_489),
.A2(n_336),
.B(n_329),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_486),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_522),
.B(n_405),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_484),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_497),
.B(n_288),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_503),
.B(n_190),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_483),
.A2(n_450),
.B1(n_346),
.B2(n_353),
.Y(n_660)
);

CKINVDCx6p67_ASAP7_75t_R g661 ( 
.A(n_454),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_503),
.B(n_191),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_504),
.Y(n_663)
);

NOR2x1p5_ASAP7_75t_L g664 ( 
.A(n_516),
.B(n_354),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_504),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_483),
.A2(n_238),
.B1(n_359),
.B2(n_273),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_467),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_484),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_484),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_485),
.A2(n_354),
.B1(n_251),
.B2(n_305),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_508),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_468),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_499),
.B(n_340),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_508),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_524),
.A2(n_293),
.B1(n_335),
.B2(n_350),
.Y(n_675)
);

INVx11_ASAP7_75t_L g676 ( 
.A(n_511),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_484),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_508),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_505),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_505),
.B(n_191),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_522),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_551),
.A2(n_520),
.B1(n_489),
.B2(n_502),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_593),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_531),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_546),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_603),
.B(n_485),
.Y(n_686)
);

AO22x1_ASAP7_75t_L g687 ( 
.A1(n_534),
.A2(n_479),
.B1(n_481),
.B2(n_530),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_608),
.B(n_522),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_631),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_583),
.B(n_505),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_534),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_563),
.B(n_507),
.Y(n_692)
);

BUFx5_ASAP7_75t_L g693 ( 
.A(n_534),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_546),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_534),
.B(n_505),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_573),
.Y(n_696)
);

BUFx6f_ASAP7_75t_SL g697 ( 
.A(n_610),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_537),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_597),
.B(n_527),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_582),
.B(n_458),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_547),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_507),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_545),
.B(n_517),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_561),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_534),
.B(n_517),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_545),
.B(n_517),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_604),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_534),
.B(n_517),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_554),
.B(n_527),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_544),
.A2(n_524),
.B1(n_511),
.B2(n_463),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_592),
.B(n_526),
.C(n_219),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_561),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_589),
.B(n_527),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_562),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_621),
.B(n_527),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_544),
.A2(n_524),
.B1(n_511),
.B2(n_463),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_549),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_550),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_562),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_549),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_655),
.B(n_528),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_553),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_655),
.B(n_528),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_553),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_617),
.B(n_528),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_544),
.A2(n_511),
.B1(n_463),
.B2(n_528),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_679),
.B(n_528),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_679),
.B(n_528),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_557),
.B(n_558),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_631),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_572),
.B(n_502),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_550),
.Y(n_733)
);

AO22x2_ASAP7_75t_L g734 ( 
.A1(n_539),
.A2(n_520),
.B1(n_509),
.B2(n_523),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_572),
.B(n_195),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_535),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_566),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_560),
.B(n_459),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_572),
.B(n_195),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_568),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_574),
.B(n_462),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_566),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_568),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_569),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_569),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_544),
.A2(n_511),
.B1(n_509),
.B2(n_462),
.Y(n_746)
);

AND2x6_ASAP7_75t_SL g747 ( 
.A(n_610),
.B(n_364),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_604),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_595),
.B(n_509),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_593),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_533),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_584),
.B(n_511),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_572),
.B(n_196),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_650),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_560),
.B(n_213),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_557),
.B(n_372),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_571),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_572),
.B(n_196),
.Y(n_758)
);

NOR2xp67_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_199),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_620),
.B(n_511),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_571),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_588),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_624),
.B(n_199),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_630),
.B(n_203),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_558),
.B(n_203),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_650),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_598),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_560),
.B(n_221),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_593),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_598),
.Y(n_770)
);

BUFx6f_ASAP7_75t_SL g771 ( 
.A(n_610),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_633),
.B(n_204),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_578),
.B(n_231),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_599),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_578),
.A2(n_204),
.B1(n_357),
.B2(n_330),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_667),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_637),
.B(n_208),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_641),
.B(n_208),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_596),
.B(n_328),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_565),
.Y(n_780)
);

INVxp33_ASAP7_75t_L g781 ( 
.A(n_628),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_593),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_596),
.B(n_328),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_652),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_610),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_657),
.B(n_330),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_SL g787 ( 
.A1(n_672),
.A2(n_372),
.B1(n_401),
.B2(n_397),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_544),
.B(n_337),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_544),
.B(n_337),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_606),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_654),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_596),
.B(n_343),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_596),
.B(n_343),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_636),
.B(n_242),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_643),
.B(n_344),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_643),
.B(n_606),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_643),
.B(n_344),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_673),
.A2(n_341),
.B(n_342),
.C(n_355),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_619),
.B(n_349),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_619),
.B(n_349),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_656),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_653),
.A2(n_335),
.B1(n_350),
.B2(n_257),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_653),
.A2(n_356),
.B1(n_246),
.B2(n_255),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_656),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_654),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_666),
.B(n_258),
.C(n_294),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_642),
.B(n_265),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_267),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_649),
.B(n_357),
.Y(n_810)
);

BUFx5_ASAP7_75t_L g811 ( 
.A(n_542),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_596),
.B(n_351),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_659),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_668),
.A2(n_464),
.B(n_461),
.C(n_452),
.Y(n_814)
);

NOR2xp67_ASAP7_75t_L g815 ( 
.A(n_564),
.B(n_672),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_661),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_635),
.B(n_351),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_668),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_669),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_677),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_635),
.B(n_351),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_681),
.B(n_280),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_622),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_661),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_681),
.B(n_281),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_591),
.A2(n_680),
.B1(n_647),
.B2(n_648),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_658),
.A2(n_662),
.B1(n_605),
.B2(n_639),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_625),
.B(n_286),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_536),
.B(n_297),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_540),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_575),
.B(n_301),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_576),
.B(n_304),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_664),
.A2(n_210),
.B1(n_211),
.B2(n_218),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_676),
.Y(n_835)
);

INVx8_ASAP7_75t_L g836 ( 
.A(n_559),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_653),
.B(n_308),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_532),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_663),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_536),
.B(n_587),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_738),
.B(n_663),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_693),
.B(n_635),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_698),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_698),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_691),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_691),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_762),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_767),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_770),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_738),
.B(n_665),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_700),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_689),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_SL g853 ( 
.A1(n_787),
.A2(n_401),
.B1(n_397),
.B2(n_731),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_750),
.B(n_645),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_782),
.B(n_670),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_766),
.Y(n_856)
);

BUFx4f_ASAP7_75t_L g857 ( 
.A(n_719),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_816),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_785),
.B(n_586),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_693),
.B(n_635),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_781),
.B(n_556),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_688),
.B(n_665),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_733),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_835),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_774),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_734),
.A2(n_675),
.B1(n_678),
.B2(n_674),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_781),
.B(n_646),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_SL g868 ( 
.A1(n_688),
.A2(n_581),
.B(n_548),
.C(n_567),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_717),
.B(n_660),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_835),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_686),
.B(n_671),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_683),
.B(n_586),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_780),
.Y(n_873)
);

BUFx4f_ASAP7_75t_L g874 ( 
.A(n_756),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_776),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_686),
.B(n_671),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_766),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_773),
.A2(n_587),
.B1(n_600),
.B2(n_602),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_790),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_685),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_711),
.B(n_323),
.C(n_313),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_836),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_692),
.B(n_682),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_693),
.B(n_532),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_682),
.B(n_678),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_683),
.B(n_587),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_734),
.A2(n_651),
.B1(n_601),
.B2(n_640),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_773),
.A2(n_324),
.B1(n_327),
.B2(n_651),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_736),
.B(n_824),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_703),
.B(n_600),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_838),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_694),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_701),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_SL g894 ( 
.A(n_755),
.B(n_260),
.C(n_252),
.Y(n_894)
);

NOR2x2_ASAP7_75t_L g895 ( 
.A(n_697),
.B(n_585),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_769),
.B(n_600),
.Y(n_896)
);

AND2x6_ASAP7_75t_SL g897 ( 
.A(n_755),
.B(n_607),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_706),
.B(n_696),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_769),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_741),
.B(n_602),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_751),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_684),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_718),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_827),
.B(n_536),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_702),
.B(n_602),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_836),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_796),
.B(n_548),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_690),
.B(n_548),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_721),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_723),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_693),
.B(n_532),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_693),
.B(n_532),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_768),
.B(n_786),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_693),
.B(n_532),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_838),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_730),
.B(n_567),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_825),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_805),
.B(n_542),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_828),
.B(n_577),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_695),
.B(n_705),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_699),
.A2(n_581),
.B(n_577),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_740),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_836),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_805),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_708),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_687),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_754),
.Y(n_928)
);

NOR2x1p5_ASAP7_75t_L g929 ( 
.A(n_795),
.B(n_797),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_743),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_757),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_761),
.B(n_726),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_SL g933 ( 
.A1(n_803),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_801),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_734),
.B(n_581),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_811),
.B(n_559),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_803),
.A2(n_585),
.B1(n_640),
.B2(n_638),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_830),
.B(n_829),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_707),
.B(n_559),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_838),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_830),
.B(n_607),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_804),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_794),
.B(n_570),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_715),
.B(n_611),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_811),
.B(n_559),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_798),
.A2(n_612),
.B(n_611),
.C(n_615),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_697),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_784),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_838),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_791),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_722),
.B(n_615),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_818),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_771),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_819),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_707),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_771),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_748),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_815),
.B(n_594),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_811),
.B(n_559),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_724),
.B(n_618),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_802),
.A2(n_601),
.B1(n_638),
.B2(n_634),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_806),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_820),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_794),
.A2(n_618),
.B1(n_580),
.B2(n_579),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_821),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_813),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_747),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_765),
.B(n_594),
.Y(n_968)
);

INVxp33_ASAP7_75t_L g969 ( 
.A(n_808),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_749),
.B(n_609),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_831),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_704),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_699),
.A2(n_538),
.B(n_555),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_712),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_759),
.B(n_609),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_748),
.B(n_613),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_714),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_713),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_807),
.B(n_613),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_720),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_728),
.B(n_616),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_832),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_811),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_802),
.A2(n_837),
.B1(n_839),
.B2(n_746),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_737),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_811),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_742),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_799),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_808),
.B(n_538),
.Y(n_989)
);

INVx5_ASAP7_75t_L g990 ( 
.A(n_744),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_809),
.A2(n_626),
.B1(n_634),
.B2(n_632),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_745),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_729),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_840),
.A2(n_676),
.B1(n_632),
.B2(n_629),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_833),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_709),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_752),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_760),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_809),
.A2(n_627),
.B1(n_626),
.B2(n_623),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_732),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_732),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_823),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_746),
.B(n_623),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_812),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_834),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_775),
.B(n_627),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_840),
.B(n_629),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_763),
.B(n_541),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_727),
.B(n_541),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_L g1010 ( 
.A(n_764),
.B(n_590),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_772),
.B(n_543),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_777),
.B(n_543),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_826),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_812),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_778),
.B(n_555),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_817),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_862),
.A2(n_735),
.B(n_758),
.Y(n_1017)
);

OR2x2_ASAP7_75t_SL g1018 ( 
.A(n_869),
.B(n_800),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_851),
.B(n_798),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_914),
.B(n_810),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_883),
.A2(n_814),
.B(n_822),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_857),
.Y(n_1022)
);

CKINVDCx8_ASAP7_75t_R g1023 ( 
.A(n_897),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_947),
.Y(n_1024)
);

OR2x6_ASAP7_75t_SL g1025 ( 
.A(n_1005),
.B(n_788),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_941),
.A2(n_753),
.B(n_735),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_932),
.A2(n_739),
.B(n_793),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_914),
.A2(n_792),
.B(n_779),
.C(n_783),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_SL g1029 ( 
.A(n_852),
.B(n_779),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_857),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_969),
.B(n_789),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_875),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_938),
.A2(n_792),
.B(n_783),
.C(n_793),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_863),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_1010),
.A2(n_973),
.B(n_885),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_847),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_876),
.B(n_889),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_841),
.A2(n_739),
.B(n_822),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_845),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_873),
.Y(n_1040)
);

BUFx12f_ASAP7_75t_L g1041 ( 
.A(n_918),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_973),
.A2(n_817),
.B(n_590),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_845),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_898),
.B(n_710),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_874),
.B(n_969),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_874),
.B(n_727),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_904),
.A2(n_716),
.B1(n_710),
.B2(n_274),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_858),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_889),
.B(n_716),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_SL g1050 ( 
.A(n_894),
.B(n_311),
.C(n_223),
.Y(n_1050)
);

OAI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_867),
.A2(n_317),
.B1(n_224),
.B2(n_220),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_858),
.B(n_552),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_988),
.B(n_552),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_867),
.B(n_3),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_894),
.B(n_227),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_850),
.A2(n_279),
.B(n_229),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_854),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_904),
.A2(n_849),
.B1(n_865),
.B2(n_848),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_906),
.B(n_230),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_906),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_933),
.A2(n_292),
.B1(n_235),
.B2(n_240),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_868),
.A2(n_466),
.B(n_464),
.C(n_461),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_861),
.B(n_232),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_R g1064 ( 
.A(n_899),
.B(n_234),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_871),
.B(n_3),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_879),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_921),
.A2(n_466),
.B(n_461),
.C(n_452),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_853),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1002),
.B(n_4),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_861),
.B(n_249),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_880),
.Y(n_1071)
);

BUFx12f_ASAP7_75t_L g1072 ( 
.A(n_854),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1013),
.B(n_4),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_996),
.B(n_5),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_845),
.B(n_183),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_900),
.A2(n_298),
.B(n_312),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_970),
.A2(n_287),
.B(n_307),
.Y(n_1077)
);

BUFx4f_ASAP7_75t_SL g1078 ( 
.A(n_958),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_978),
.A2(n_264),
.B(n_306),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_921),
.A2(n_262),
.B(n_261),
.C(n_303),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_901),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_892),
.B(n_9),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_978),
.A2(n_456),
.B(n_300),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_982),
.B(n_995),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_906),
.B(n_351),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_855),
.B(n_12),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_886),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_924),
.B(n_351),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_893),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_903),
.B(n_909),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_910),
.B(n_13),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_946),
.A2(n_456),
.B(n_351),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_913),
.B(n_14),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_923),
.B(n_15),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_927),
.B(n_73),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_855),
.B(n_16),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_920),
.A2(n_205),
.B(n_183),
.C(n_456),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_888),
.A2(n_205),
.B1(n_183),
.B2(n_456),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_845),
.B(n_183),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_843),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_930),
.B(n_19),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_888),
.A2(n_205),
.B1(n_456),
.B2(n_27),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_886),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_953),
.B(n_19),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_920),
.A2(n_22),
.B(n_27),
.C(n_28),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_931),
.B(n_926),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_944),
.A2(n_76),
.B(n_156),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_926),
.B(n_22),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_881),
.B(n_29),
.C(n_32),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_971),
.B(n_33),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_844),
.Y(n_1111)
);

OR2x6_ASAP7_75t_SL g1112 ( 
.A(n_895),
.B(n_36),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_855),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_924),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_891),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_881),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.C(n_49),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_872),
.B(n_38),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_934),
.A2(n_965),
.B1(n_952),
.B2(n_954),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_929),
.A2(n_39),
.B(n_52),
.C(n_53),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_924),
.B(n_872),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_955),
.B(n_54),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_942),
.A2(n_55),
.B1(n_60),
.B2(n_66),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_SL g1123 ( 
.A(n_963),
.B(n_90),
.C(n_92),
.Y(n_1123)
);

INVx6_ASAP7_75t_L g1124 ( 
.A(n_924),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_846),
.B(n_919),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_953),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_984),
.A2(n_98),
.B1(n_102),
.B2(n_116),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_974),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_890),
.B(n_124),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_856),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_989),
.A2(n_134),
.B(n_140),
.C(n_145),
.Y(n_1131)
);

AO32x1_ASAP7_75t_L g1132 ( 
.A1(n_1000),
.A2(n_152),
.A3(n_174),
.B1(n_1001),
.B2(n_994),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_956),
.B(n_967),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_957),
.B(n_925),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_877),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_993),
.B(n_989),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_882),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_846),
.B(n_919),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_917),
.A2(n_905),
.B(n_868),
.C(n_946),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_985),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_SL g1141 ( 
.A(n_864),
.B(n_870),
.Y(n_1141)
);

OR2x6_ASAP7_75t_SL g1142 ( 
.A(n_895),
.B(n_935),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_902),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_956),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_922),
.A2(n_884),
.B(n_912),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_951),
.A2(n_960),
.B(n_1007),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_943),
.A2(n_878),
.B(n_1006),
.C(n_964),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_SL g1148 ( 
.A(n_896),
.B(n_983),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_987),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_975),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_943),
.B(n_925),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_896),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_891),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_891),
.Y(n_1154)
);

BUFx4f_ASAP7_75t_L g1155 ( 
.A(n_1006),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_972),
.B(n_977),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_957),
.B(n_980),
.Y(n_1157)
);

OR2x6_ASAP7_75t_SL g1158 ( 
.A(n_968),
.B(n_907),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_908),
.A2(n_1011),
.B(n_1015),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_928),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_859),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1008),
.A2(n_1012),
.B(n_922),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1036),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1041),
.Y(n_1164)
);

AOI211x1_ASAP7_75t_L g1165 ( 
.A1(n_1058),
.A2(n_1003),
.B(n_997),
.C(n_998),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1032),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1063),
.A2(n_859),
.B1(n_984),
.B2(n_979),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1159),
.A2(n_1146),
.B(n_1162),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1020),
.A2(n_986),
.B(n_983),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1070),
.A2(n_842),
.B(n_860),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1114),
.Y(n_1172)
);

AO32x2_ASAP7_75t_L g1173 ( 
.A1(n_1058),
.A2(n_986),
.A3(n_887),
.B1(n_866),
.B2(n_1009),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1037),
.B(n_949),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_1117),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1084),
.B(n_980),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1139),
.A2(n_1003),
.B(n_991),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_SL g1178 ( 
.A1(n_1080),
.A2(n_945),
.B(n_936),
.C(n_959),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1087),
.B(n_950),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1028),
.A2(n_842),
.B(n_860),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1127),
.A2(n_916),
.B(n_979),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1155),
.B(n_891),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1092),
.A2(n_1009),
.B(n_884),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1024),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1147),
.A2(n_1016),
.A3(n_1014),
.B(n_1004),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1105),
.A2(n_911),
.B(n_915),
.C(n_981),
.Y(n_1186)
);

AO22x2_ASAP7_75t_L g1187 ( 
.A1(n_1127),
.A2(n_962),
.B1(n_948),
.B2(n_966),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1040),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_R g1189 ( 
.A(n_1068),
.B(n_976),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1038),
.A2(n_911),
.B(n_887),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1026),
.A2(n_916),
.B(n_949),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1086),
.A2(n_937),
.B1(n_976),
.B2(n_999),
.Y(n_1192)
);

CKINVDCx6p67_ASAP7_75t_R g1193 ( 
.A(n_1048),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1126),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1017),
.A2(n_937),
.B(n_981),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1075),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1097),
.A2(n_866),
.A3(n_961),
.B(n_992),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1061),
.A2(n_990),
.B1(n_940),
.B2(n_949),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1027),
.A2(n_990),
.B(n_961),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1156),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1087),
.B(n_990),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1150),
.Y(n_1202)
);

O2A1O1Ixp5_ASAP7_75t_L g1203 ( 
.A1(n_1083),
.A2(n_940),
.B(n_939),
.C(n_990),
.Y(n_1203)
);

AO21x2_ASAP7_75t_L g1204 ( 
.A1(n_1062),
.A2(n_992),
.B(n_940),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1151),
.A2(n_992),
.B(n_1033),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_SL g1206 ( 
.A(n_1155),
.B(n_992),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1054),
.B(n_1019),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1021),
.A2(n_1065),
.B(n_1083),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1107),
.A2(n_1129),
.B(n_1088),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1061),
.A2(n_1098),
.B1(n_1049),
.B2(n_1090),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1098),
.A2(n_1067),
.B(n_1074),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1136),
.A2(n_1047),
.B(n_1075),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1085),
.A2(n_1118),
.B(n_1152),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1044),
.A2(n_1057),
.B1(n_1046),
.B2(n_1102),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1148),
.A2(n_1132),
.B(n_1075),
.Y(n_1215)
);

OR2x6_ASAP7_75t_L g1216 ( 
.A(n_1099),
.B(n_1161),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1031),
.A2(n_1069),
.B(n_1073),
.C(n_1119),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1118),
.A2(n_1152),
.B(n_1122),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1122),
.A2(n_1137),
.B(n_1106),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1103),
.B(n_1034),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1109),
.A2(n_1050),
.B(n_1116),
.C(n_1108),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1137),
.A2(n_1120),
.B(n_1081),
.Y(n_1222)
);

O2A1O1Ixp5_ASAP7_75t_SL g1223 ( 
.A1(n_1128),
.A2(n_1149),
.B(n_1140),
.C(n_1071),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1082),
.A2(n_1091),
.B(n_1093),
.Y(n_1224)
);

AND2x2_ASAP7_75t_SL g1225 ( 
.A(n_1096),
.B(n_1113),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_L g1226 ( 
.A(n_1114),
.B(n_1153),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1103),
.B(n_1034),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1157),
.A2(n_1110),
.B(n_1101),
.C(n_1094),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1125),
.A2(n_1138),
.B(n_1066),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1089),
.A2(n_1100),
.B(n_1135),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1111),
.A2(n_1130),
.B(n_1134),
.Y(n_1231)
);

NOR4xp25_ASAP7_75t_L g1232 ( 
.A(n_1131),
.B(n_1023),
.C(n_1045),
.D(n_1144),
.Y(n_1232)
);

AND2x6_ASAP7_75t_L g1233 ( 
.A(n_1039),
.B(n_1043),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1148),
.A2(n_1132),
.B(n_1099),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1143),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1059),
.A2(n_1076),
.B(n_1077),
.Y(n_1236)
);

O2A1O1Ixp5_ASAP7_75t_L g1237 ( 
.A1(n_1029),
.A2(n_1141),
.B(n_1154),
.C(n_1056),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1132),
.A2(n_1099),
.B(n_1079),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1160),
.A2(n_1053),
.B(n_1121),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1018),
.B(n_1133),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_1052),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1123),
.A2(n_1022),
.B(n_1030),
.C(n_1158),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1142),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1051),
.B(n_1112),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1115),
.A2(n_1060),
.B(n_1043),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1115),
.B(n_1055),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1115),
.A2(n_1025),
.B(n_1095),
.C(n_1078),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1064),
.A2(n_1104),
.B(n_1124),
.C(n_1060),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1072),
.B(n_1104),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_883),
.B(n_914),
.C(n_1063),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1037),
.B(n_733),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1041),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1054),
.B(n_781),
.Y(n_1253)
);

NOR2x1_ASAP7_75t_SL g1254 ( 
.A(n_1114),
.B(n_1075),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1037),
.B(n_969),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1037),
.B(n_686),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1063),
.A2(n_914),
.B(n_883),
.C(n_1070),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1041),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1116),
.A2(n_883),
.B1(n_1105),
.B2(n_682),
.C(n_1058),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1037),
.B(n_686),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1087),
.B(n_1103),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1087),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1037),
.B(n_686),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1037),
.B(n_686),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1036),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1063),
.A2(n_914),
.B(n_883),
.C(n_1070),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1037),
.B(n_883),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1041),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1037),
.B(n_686),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1063),
.A2(n_883),
.B1(n_686),
.B2(n_1070),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1054),
.B(n_781),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1036),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1037),
.B(n_686),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1037),
.B(n_686),
.Y(n_1282)
);

NOR2x1_ASAP7_75t_R g1283 ( 
.A(n_1041),
.B(n_689),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1063),
.A2(n_883),
.B1(n_686),
.B2(n_1070),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1041),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1020),
.A2(n_883),
.B1(n_914),
.B2(n_686),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1063),
.A2(n_591),
.B1(n_660),
.B2(n_686),
.C(n_773),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1036),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1037),
.B(n_686),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1159),
.A2(n_883),
.B(n_938),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_SL g1294 ( 
.A(n_1041),
.B(n_689),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1114),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1063),
.A2(n_914),
.B(n_883),
.C(n_1070),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1063),
.A2(n_883),
.B1(n_686),
.B2(n_1070),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1037),
.B(n_883),
.Y(n_1298)
);

O2A1O1Ixp5_ASAP7_75t_L g1299 ( 
.A1(n_1063),
.A2(n_883),
.B(n_914),
.C(n_1070),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1139),
.A2(n_883),
.B(n_978),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1301)
);

O2A1O1Ixp5_ASAP7_75t_SL g1302 ( 
.A1(n_1058),
.A2(n_447),
.B(n_1127),
.C(n_457),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1037),
.B(n_686),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1037),
.B(n_686),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1020),
.A2(n_883),
.B(n_914),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1035),
.A2(n_1145),
.B(n_1042),
.Y(n_1307)
);

O2A1O1Ixp5_ASAP7_75t_L g1308 ( 
.A1(n_1257),
.A2(n_1270),
.B(n_1296),
.C(n_1299),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1277),
.A2(n_1297),
.B1(n_1284),
.B2(n_1288),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1172),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1188),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1207),
.B(n_1253),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1169),
.A2(n_1272),
.B(n_1260),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1281),
.A2(n_1292),
.B(n_1291),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1163),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1284),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1287),
.B(n_1256),
.Y(n_1317)
);

CKINVDCx6p67_ASAP7_75t_R g1318 ( 
.A(n_1164),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1278),
.B(n_1255),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1301),
.A2(n_1307),
.B(n_1306),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1208),
.A2(n_1177),
.B(n_1190),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1244),
.A2(n_1189),
.B1(n_1261),
.B2(n_1241),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1199),
.A2(n_1211),
.B(n_1195),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1263),
.B(n_1245),
.Y(n_1325)
);

AOI21xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1184),
.A2(n_1286),
.B(n_1290),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1262),
.B(n_1267),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1191),
.A2(n_1205),
.B(n_1209),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1269),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1279),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1172),
.Y(n_1331)
);

CKINVDCx6p67_ASAP7_75t_R g1332 ( 
.A(n_1258),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1180),
.A2(n_1239),
.B(n_1285),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1251),
.B(n_1240),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1293),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1250),
.A2(n_1221),
.B(n_1217),
.C(n_1305),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1231),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1185),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1220),
.B(n_1227),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1208),
.A2(n_1177),
.B(n_1219),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1261),
.A2(n_1211),
.B(n_1224),
.C(n_1210),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1289),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1224),
.A2(n_1167),
.B(n_1300),
.C(n_1273),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1266),
.A2(n_1274),
.B(n_1213),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1218),
.A2(n_1170),
.B(n_1203),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1302),
.A2(n_1186),
.B(n_1300),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1236),
.A2(n_1171),
.B(n_1181),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1228),
.A2(n_1198),
.A3(n_1187),
.B(n_1235),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1265),
.B(n_1166),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1223),
.A2(n_1222),
.B(n_1229),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1194),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1268),
.A2(n_1304),
.B(n_1276),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1237),
.A2(n_1174),
.B(n_1212),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1200),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1185),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_SL g1356 ( 
.A1(n_1242),
.A2(n_1271),
.B(n_1298),
.C(n_1303),
.Y(n_1356)
);

BUFx4_ASAP7_75t_SL g1357 ( 
.A(n_1202),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1280),
.B(n_1282),
.Y(n_1358)
);

BUFx4_ASAP7_75t_R g1359 ( 
.A(n_1254),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1232),
.A2(n_1167),
.B(n_1178),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1214),
.A2(n_1187),
.B1(n_1225),
.B2(n_1192),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1175),
.B(n_1182),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1232),
.A2(n_1248),
.B(n_1247),
.C(n_1243),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1246),
.A2(n_1201),
.B(n_1226),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1179),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1175),
.A2(n_1294),
.B1(n_1249),
.B2(n_1206),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1263),
.A2(n_1265),
.B1(n_1183),
.B2(n_1176),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1185),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1173),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1173),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1165),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1196),
.B(n_1216),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1165),
.Y(n_1373)
);

AOI22x1_ASAP7_75t_L g1374 ( 
.A1(n_1172),
.A2(n_1295),
.B1(n_1275),
.B2(n_1252),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1193),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1216),
.Y(n_1376)
);

INVx5_ASAP7_75t_L g1377 ( 
.A(n_1196),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1173),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1197),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1295),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1204),
.A2(n_1197),
.B(n_1233),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1197),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1295),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1283),
.A2(n_1284),
.B(n_1277),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1277),
.A2(n_1297),
.B1(n_1284),
.B2(n_1288),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1202),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1277),
.A2(n_1297),
.B1(n_1284),
.B2(n_1270),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1284),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1284),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1257),
.A2(n_1296),
.B(n_1270),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1288),
.B(n_1284),
.C(n_1277),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1256),
.B(n_1262),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1202),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1188),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1168),
.A2(n_1260),
.B(n_1169),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1207),
.B(n_1253),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1169),
.A2(n_1272),
.B(n_1260),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1207),
.B(n_1253),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1230),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1251),
.B(n_1240),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1210),
.A2(n_415),
.B1(n_429),
.B2(n_411),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1188),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1284),
.Y(n_1407)
);

BUFx4_ASAP7_75t_SL g1408 ( 
.A(n_1202),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1163),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1163),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1168),
.A2(n_1260),
.B(n_1169),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1168),
.A2(n_1260),
.B(n_1169),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1169),
.A2(n_1272),
.B(n_1260),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1202),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1174),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1224),
.A2(n_1284),
.B(n_1277),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1163),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1168),
.A2(n_1260),
.B(n_1169),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1169),
.A2(n_1272),
.B(n_1260),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1163),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1215),
.A2(n_1234),
.B(n_1238),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1284),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1163),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1168),
.A2(n_1260),
.B(n_1169),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1163),
.Y(n_1426)
);

NAND2x1p5_ASAP7_75t_L g1427 ( 
.A(n_1196),
.B(n_1114),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1163),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1277),
.B(n_1284),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1163),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1169),
.A2(n_1272),
.B(n_1260),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1393),
.A2(n_1387),
.B1(n_1407),
.B2(n_1316),
.C(n_1389),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_SL g1433 ( 
.A1(n_1429),
.A2(n_1391),
.B(n_1423),
.C(n_1384),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1315),
.Y(n_1434)
);

O2A1O1Ixp5_ASAP7_75t_L g1435 ( 
.A1(n_1429),
.A2(n_1392),
.B(n_1308),
.C(n_1341),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1335),
.A2(n_1344),
.B(n_1328),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1317),
.B(n_1358),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1343),
.A2(n_1308),
.B(n_1341),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1402),
.B(n_1319),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1349),
.B(n_1339),
.Y(n_1440)
);

BUFx8_ASAP7_75t_L g1441 ( 
.A(n_1398),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1343),
.A2(n_1317),
.B(n_1309),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1360),
.B(n_1325),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1397),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1334),
.B(n_1404),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1358),
.B(n_1327),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1323),
.B(n_1406),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1357),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1394),
.B(n_1385),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1363),
.A2(n_1336),
.B(n_1352),
.Y(n_1450)
);

O2A1O1Ixp5_ASAP7_75t_L g1451 ( 
.A1(n_1415),
.A2(n_1371),
.B(n_1373),
.C(n_1362),
.Y(n_1451)
);

AND2x4_ASAP7_75t_SL g1452 ( 
.A(n_1414),
.B(n_1318),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1365),
.B(n_1329),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1417),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1330),
.B(n_1342),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1350),
.A2(n_1333),
.B(n_1347),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1409),
.B(n_1410),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1325),
.B(n_1372),
.Y(n_1458)
);

INVx3_ASAP7_75t_SL g1459 ( 
.A(n_1414),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1340),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1311),
.B(n_1418),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1311),
.B(n_1421),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1424),
.B(n_1426),
.Y(n_1463)
);

OAI22x1_ASAP7_75t_L g1464 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_1374),
.B2(n_1386),
.Y(n_1464)
);

O2A1O1Ixp5_ASAP7_75t_L g1465 ( 
.A1(n_1368),
.A2(n_1355),
.B(n_1338),
.C(n_1378),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1313),
.A2(n_1314),
.B(n_1413),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1361),
.A2(n_1405),
.B(n_1346),
.C(n_1369),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1354),
.B(n_1367),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1356),
.B(n_1405),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1397),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1325),
.B(n_1372),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1416),
.B(n_1383),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1356),
.B(n_1383),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1340),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1357),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1361),
.B(n_1310),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1346),
.A2(n_1431),
.B(n_1320),
.Y(n_1477)
);

O2A1O1Ixp5_ASAP7_75t_L g1478 ( 
.A1(n_1338),
.A2(n_1355),
.B(n_1370),
.C(n_1369),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1367),
.B(n_1376),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1370),
.A2(n_1353),
.B(n_1382),
.C(n_1381),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1401),
.A2(n_1420),
.B(n_1345),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1380),
.B(n_1331),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1348),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1380),
.B(n_1364),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1380),
.B(n_1322),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1375),
.A2(n_1332),
.B1(n_1322),
.B2(n_1351),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1322),
.B(n_1324),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1324),
.A2(n_1321),
.B(n_1422),
.C(n_1396),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1408),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1375),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1351),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1353),
.A2(n_1337),
.B(n_1403),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1321),
.B(n_1396),
.Y(n_1493)
);

O2A1O1Ixp5_ASAP7_75t_L g1494 ( 
.A1(n_1379),
.A2(n_1395),
.B(n_1422),
.C(n_1390),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1388),
.B(n_1395),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1390),
.A2(n_1427),
.B(n_1425),
.C(n_1419),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1359),
.A2(n_1377),
.B(n_1399),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1412),
.B(n_1419),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1425),
.A2(n_1385),
.B1(n_1309),
.B2(n_1284),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1429),
.A2(n_1284),
.B(n_1297),
.C(n_1277),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1315),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1340),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1317),
.B(n_1358),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1309),
.A2(n_1385),
.B1(n_1284),
.B2(n_1297),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1393),
.A2(n_1270),
.B(n_1257),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1315),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1429),
.A2(n_1284),
.B(n_1297),
.C(n_1277),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1317),
.B(n_1358),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1339),
.B(n_1334),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1387),
.A2(n_1257),
.B(n_1296),
.C(n_1270),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1309),
.A2(n_1385),
.B1(n_1284),
.B2(n_1297),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1312),
.B(n_1400),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1340),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_1326),
.B(n_1366),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1312),
.B(n_1400),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1317),
.B(n_1358),
.Y(n_1517)
);

O2A1O1Ixp5_ASAP7_75t_L g1518 ( 
.A1(n_1316),
.A2(n_1391),
.B(n_1407),
.C(n_1389),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1315),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1340),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1434),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1442),
.B(n_1432),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1460),
.B(n_1474),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1501),
.B(n_1508),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1432),
.B(n_1458),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1502),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1487),
.B(n_1485),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1493),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1507),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1519),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1503),
.B(n_1514),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1494),
.A2(n_1438),
.B(n_1480),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1503),
.B(n_1514),
.Y(n_1533)
);

AO21x2_ASAP7_75t_L g1534 ( 
.A1(n_1488),
.A2(n_1480),
.B(n_1495),
.Y(n_1534)
);

AOI211xp5_ASAP7_75t_L g1535 ( 
.A1(n_1450),
.A2(n_1506),
.B(n_1505),
.C(n_1512),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1467),
.A2(n_1508),
.B(n_1501),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_SL g1537 ( 
.A(n_1511),
.B(n_1442),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1478),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1457),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1478),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1437),
.B(n_1504),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1520),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1492),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1463),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1455),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1509),
.B(n_1517),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1499),
.B(n_1456),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1444),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1456),
.B(n_1477),
.Y(n_1550)
);

AO21x2_ASAP7_75t_L g1551 ( 
.A1(n_1483),
.A2(n_1496),
.B(n_1500),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1456),
.B(n_1477),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1440),
.B(n_1479),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1453),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1465),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1465),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1496),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1451),
.A2(n_1435),
.B(n_1518),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1461),
.B(n_1462),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1497),
.B(n_1443),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1466),
.B(n_1436),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1441),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1484),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1472),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1433),
.B(n_1449),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1433),
.B(n_1454),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1481),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1481),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1541),
.B(n_1454),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1522),
.A2(n_1469),
.B1(n_1476),
.B2(n_1447),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1521),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1542),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1567),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1548),
.B(n_1443),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1548),
.B(n_1471),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1543),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1522),
.A2(n_1515),
.B1(n_1439),
.B2(n_1443),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1446),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1547),
.B(n_1435),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1542),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1516),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1539),
.B(n_1511),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1550),
.B(n_1552),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1550),
.B(n_1513),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1528),
.B(n_1518),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1528),
.B(n_1523),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1527),
.B(n_1510),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1527),
.B(n_1445),
.Y(n_1588)
);

OR2x2_ASAP7_75t_SL g1589 ( 
.A(n_1532),
.B(n_1473),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1552),
.B(n_1468),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1486),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1563),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1482),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1526),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1582),
.B(n_1546),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1577),
.A2(n_1535),
.B1(n_1524),
.B2(n_1565),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1585),
.A2(n_1536),
.B1(n_1537),
.B2(n_1524),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1575),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1588),
.B(n_1553),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1577),
.A2(n_1535),
.B1(n_1565),
.B2(n_1525),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1570),
.A2(n_1536),
.B1(n_1537),
.B2(n_1525),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1571),
.Y(n_1604)
);

OAI33xp33_ASAP7_75t_L g1605 ( 
.A1(n_1582),
.A2(n_1546),
.A3(n_1545),
.B1(n_1566),
.B2(n_1554),
.B3(n_1544),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1586),
.B(n_1559),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1572),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1585),
.A2(n_1566),
.B(n_1525),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1594),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1585),
.A2(n_1536),
.B1(n_1525),
.B2(n_1557),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1575),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1573),
.A2(n_1557),
.B(n_1556),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1579),
.B(n_1544),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1570),
.A2(n_1556),
.B1(n_1555),
.B2(n_1563),
.C(n_1554),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1594),
.Y(n_1616)
);

OAI33xp33_ASAP7_75t_L g1617 ( 
.A1(n_1569),
.A2(n_1545),
.A3(n_1564),
.B1(n_1526),
.B2(n_1529),
.B3(n_1530),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1594),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1575),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1587),
.A2(n_1560),
.B1(n_1536),
.B2(n_1464),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1571),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1575),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1588),
.B(n_1587),
.Y(n_1623)
);

AOI322xp5_ASAP7_75t_L g1624 ( 
.A1(n_1590),
.A2(n_1555),
.A3(n_1536),
.B1(n_1540),
.B2(n_1538),
.C1(n_1533),
.C2(n_1531),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_R g1625 ( 
.A(n_1569),
.B(n_1549),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1575),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1593),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1590),
.A2(n_1534),
.B1(n_1551),
.B2(n_1532),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_1532),
.C(n_1558),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1579),
.B(n_1459),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1531),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1580),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1586),
.B(n_1564),
.Y(n_1634)
);

AOI33xp33_ASAP7_75t_L g1635 ( 
.A1(n_1591),
.A2(n_1531),
.A3(n_1533),
.B1(n_1529),
.B2(n_1530),
.B3(n_1475),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1596),
.B(n_1584),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1604),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1609),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1616),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1618),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1612),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1603),
.B(n_1574),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1598),
.B(n_1558),
.C(n_1532),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1625),
.Y(n_1644)
);

AOI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1610),
.A2(n_1534),
.B(n_1532),
.Y(n_1645)
);

INVxp33_ASAP7_75t_L g1646 ( 
.A(n_1625),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1621),
.Y(n_1647)
);

OA21x2_ASAP7_75t_L g1648 ( 
.A1(n_1629),
.A2(n_1568),
.B(n_1573),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1623),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1600),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1608),
.A2(n_1568),
.B(n_1576),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1614),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1635),
.B(n_1595),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1578),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1633),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1634),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1620),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1612),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1634),
.Y(n_1660)
);

AO21x2_ASAP7_75t_L g1661 ( 
.A1(n_1615),
.A2(n_1534),
.B(n_1538),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1605),
.A2(n_1591),
.B(n_1578),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1627),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1606),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1597),
.B(n_1549),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1660),
.B(n_1603),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1637),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1603),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1637),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1641),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1662),
.B(n_1624),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1638),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1638),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1648),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1648),
.B(n_1636),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1648),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1642),
.B(n_1611),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1649),
.B(n_1631),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1643),
.B(n_1628),
.C(n_1602),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1663),
.B(n_1619),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1653),
.B(n_1590),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1644),
.B(n_1626),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1644),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1666),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1643),
.B(n_1602),
.C(n_1601),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1657),
.B(n_1606),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1641),
.B(n_1599),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1654),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1639),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1655),
.B(n_1590),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1663),
.B(n_1622),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1639),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1640),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.B(n_1622),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1661),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1652),
.B(n_1592),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1640),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1652),
.B(n_1583),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1665),
.B(n_1607),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1649),
.B(n_1589),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1691),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1690),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_R g1707 ( 
.A(n_1684),
.B(n_1549),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1685),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1668),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1668),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1683),
.B(n_1650),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1690),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1683),
.B(n_1650),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1686),
.B(n_1645),
.C(n_1651),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1687),
.B(n_1654),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1670),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1686),
.A2(n_1658),
.B1(n_1589),
.B2(n_1664),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1672),
.B(n_1656),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1670),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1693),
.B(n_1656),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1673),
.Y(n_1722)
);

OAI21xp33_ASAP7_75t_L g1723 ( 
.A1(n_1672),
.A2(n_1591),
.B(n_1665),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.B(n_1664),
.Y(n_1724)
);

NAND2x1p5_ASAP7_75t_L g1725 ( 
.A(n_1671),
.B(n_1562),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1687),
.B(n_1661),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1673),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1703),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1701),
.B(n_1584),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1690),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1682),
.B(n_1661),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1674),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1682),
.B(n_1647),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1674),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1699),
.B(n_1647),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1680),
.A2(n_1651),
.B1(n_1617),
.B2(n_1630),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1701),
.B(n_1581),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1680),
.A2(n_1591),
.B(n_1659),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1692),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1709),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1708),
.B(n_1701),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1708),
.B(n_1703),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1699),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1732),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1725),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1715),
.B(n_1675),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1725),
.B(n_1712),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1714),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1714),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1712),
.B(n_1704),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1710),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_R g1754 ( 
.A(n_1714),
.B(n_1651),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1723),
.B(n_1704),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1728),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1736),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1706),
.Y(n_1758)
);

NAND2x1_ASAP7_75t_L g1759 ( 
.A(n_1728),
.B(n_1675),
.Y(n_1759)
);

OR2x6_ASAP7_75t_L g1760 ( 
.A(n_1713),
.B(n_1671),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1738),
.B(n_1667),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1738),
.B(n_1667),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1705),
.B(n_1676),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1711),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1716),
.B(n_1676),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1736),
.B(n_1459),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1717),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1741),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1747),
.B(n_1739),
.C(n_1718),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1754),
.A2(n_1737),
.B1(n_1731),
.B2(n_1677),
.Y(n_1770)
);

OAI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1747),
.A2(n_1742),
.B(n_1743),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1757),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1759),
.A2(n_1707),
.B(n_1677),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1745),
.B(n_1688),
.C(n_1671),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1742),
.B(n_1716),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1757),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1748),
.Y(n_1777)
);

OAI32xp33_ASAP7_75t_L g1778 ( 
.A1(n_1755),
.A2(n_1726),
.A3(n_1677),
.B1(n_1675),
.B2(n_1676),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1743),
.B(n_1729),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1757),
.Y(n_1780)
);

AO22x1_ASAP7_75t_L g1781 ( 
.A1(n_1746),
.A2(n_1562),
.B1(n_1689),
.B2(n_1688),
.Y(n_1781)
);

INVxp67_ASAP7_75t_SL g1782 ( 
.A(n_1757),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1744),
.A2(n_1721),
.B1(n_1734),
.B2(n_1589),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1753),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1744),
.B(n_1720),
.Y(n_1785)
);

OAI32xp33_ASAP7_75t_L g1786 ( 
.A1(n_1763),
.A2(n_1721),
.A3(n_1659),
.B1(n_1669),
.B2(n_1698),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1756),
.B(n_1729),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1765),
.A2(n_1669),
.B(n_1678),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1750),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1782),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1772),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1776),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1777),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1775),
.B(n_1752),
.Y(n_1794)
);

NAND2xp33_ASAP7_75t_SL g1795 ( 
.A(n_1768),
.B(n_1748),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1787),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1771),
.B(n_1751),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1769),
.B(n_1751),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1770),
.A2(n_1698),
.B1(n_1749),
.B2(n_1758),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1781),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1785),
.B(n_1751),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1795),
.A2(n_1778),
.B(n_1759),
.Y(n_1802)
);

OAI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1798),
.A2(n_1766),
.B(n_1788),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1796),
.B(n_1785),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1797),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1793),
.B(n_1751),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1800),
.B(n_1773),
.Y(n_1807)
);

NAND4xp25_ASAP7_75t_L g1808 ( 
.A(n_1789),
.B(n_1774),
.C(n_1780),
.D(n_1784),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1799),
.A2(n_1783),
.B1(n_1760),
.B2(n_1688),
.C(n_1698),
.Y(n_1809)
);

AOI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1797),
.A2(n_1786),
.B(n_1783),
.C(n_1765),
.Y(n_1810)
);

OAI222xp33_ASAP7_75t_L g1811 ( 
.A1(n_1799),
.A2(n_1760),
.B1(n_1749),
.B2(n_1758),
.C1(n_1659),
.C2(n_1767),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1790),
.A2(n_1767),
.B1(n_1764),
.B2(n_1753),
.C(n_1749),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1802),
.A2(n_1792),
.B(n_1791),
.C(n_1764),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1811),
.A2(n_1760),
.B(n_1801),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1807),
.A2(n_1758),
.B1(n_1730),
.B2(n_1713),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1804),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1809),
.A2(n_1730),
.B1(n_1760),
.B2(n_1651),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1810),
.B(n_1794),
.Y(n_1818)
);

AOI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1812),
.A2(n_1722),
.B1(n_1727),
.B2(n_1733),
.C(n_1735),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1803),
.A2(n_1760),
.B1(n_1761),
.B2(n_1762),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1820),
.B(n_1816),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1818),
.A2(n_1805),
.B(n_1808),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1815),
.Y(n_1823)
);

NOR3x1_ASAP7_75t_L g1824 ( 
.A(n_1813),
.B(n_1806),
.C(n_1491),
.Y(n_1824)
);

AOI221x1_ASAP7_75t_L g1825 ( 
.A1(n_1814),
.A2(n_1740),
.B1(n_1761),
.B2(n_1762),
.C(n_1689),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1819),
.B(n_1470),
.Y(n_1826)
);

AOI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1817),
.A2(n_1669),
.B(n_1689),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1822),
.B(n_1724),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1821),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1823),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1826),
.B(n_1689),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1827),
.A2(n_1700),
.B1(n_1692),
.B2(n_1695),
.C(n_1696),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1824),
.B(n_1678),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1829),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1828),
.B(n_1825),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1830),
.B(n_1695),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_SL g1837 ( 
.A(n_1834),
.B(n_1832),
.C(n_1833),
.Y(n_1837)
);

NOR3xp33_ASAP7_75t_L g1838 ( 
.A(n_1837),
.B(n_1835),
.C(n_1836),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1838),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1838),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1840),
.B1(n_1831),
.B2(n_1448),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1839),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1842),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1841),
.A2(n_1724),
.B1(n_1490),
.B2(n_1489),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1843),
.A2(n_1562),
.B1(n_1452),
.B2(n_1700),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1845),
.A2(n_1844),
.B1(n_1696),
.B2(n_1694),
.Y(n_1846)
);

AO21x2_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1694),
.B(n_1697),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1847),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1848),
.A2(n_1679),
.B1(n_1702),
.B2(n_1697),
.Y(n_1849)
);

AOI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1441),
.B(n_1681),
.C(n_1697),
.Y(n_1850)
);


endmodule