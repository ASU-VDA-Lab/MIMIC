module fake_jpeg_16871_n_352 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_45),
.B(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_53),
.Y(n_112)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_63),
.Y(n_73)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_24),
.Y(n_61)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_8),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_33),
.B1(n_37),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_66),
.A2(n_87),
.B1(n_79),
.B2(n_113),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_93),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_37),
.B1(n_24),
.B2(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_72),
.A2(n_90),
.B1(n_103),
.B2(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_24),
.B(n_1),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_72),
.B(n_21),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_91),
.Y(n_136)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_39),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_15),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_97),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_62),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_104),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_20),
.B1(n_32),
.B2(n_22),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_22),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_29),
.Y(n_111)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_52),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_29),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_125),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_120),
.B(n_126),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_133),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_70),
.A2(n_85),
.B1(n_78),
.B2(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_122),
.A2(n_132),
.B1(n_141),
.B2(n_156),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_123),
.A2(n_99),
.B1(n_69),
.B2(n_75),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_34),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_146),
.B1(n_84),
.B2(n_67),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_21),
.B1(n_26),
.B2(n_23),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_150),
.B1(n_74),
.B2(n_109),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_34),
.C(n_26),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_144),
.C(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_21),
.A3(n_34),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_9),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_134),
.A2(n_152),
.B1(n_157),
.B2(n_163),
.Y(n_194)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_74),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_9),
.B(n_1),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_9),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_92),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_3),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_73),
.A2(n_5),
.B(n_11),
.C(n_12),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_154),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_83),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_104),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_92),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_71),
.B(n_13),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_83),
.A2(n_0),
.B1(n_12),
.B2(n_101),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_97),
.B(n_12),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_0),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_71),
.B(n_0),
.Y(n_163)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_0),
.C(n_88),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_171),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_172),
.A2(n_156),
.B(n_163),
.C(n_165),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_191),
.Y(n_224)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_182),
.B(n_183),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_131),
.B(n_125),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_190),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_135),
.B1(n_137),
.B2(n_127),
.Y(n_231)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_84),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_89),
.B1(n_67),
.B2(n_98),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_196),
.B1(n_203),
.B2(n_197),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_86),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_196),
.A2(n_209),
.B1(n_199),
.B2(n_198),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_102),
.C(n_86),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_205),
.C(n_170),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_121),
.A2(n_89),
.B1(n_82),
.B2(n_98),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_206),
.B1(n_215),
.B2(n_142),
.Y(n_220)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_69),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_209),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_210),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_102),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_75),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_140),
.B(n_99),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_211),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_134),
.Y(n_223)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_168),
.B1(n_158),
.B2(n_151),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_124),
.A2(n_132),
.B1(n_168),
.B2(n_161),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_218),
.A2(n_231),
.B1(n_235),
.B2(n_248),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_136),
.B(n_152),
.C(n_165),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_SL g286 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_163),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_223),
.B(n_234),
.C(n_224),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_157),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_157),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_232),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_127),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_149),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_149),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_242),
.Y(n_263)
);

OR2x4_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_188),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_180),
.B(n_185),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_203),
.B1(n_187),
.B2(n_188),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_244),
.B1(n_239),
.B2(n_235),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_207),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_184),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_194),
.A2(n_170),
.B1(n_189),
.B2(n_213),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_174),
.A2(n_179),
.B1(n_200),
.B2(n_176),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_193),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_217),
.Y(n_278)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_192),
.B(n_186),
.C(n_178),
.D(n_201),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_257),
.B(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_269),
.B1(n_271),
.B2(n_225),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_275),
.C(n_216),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_255),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_226),
.B(n_219),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_282),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_222),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_284),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_226),
.A2(n_220),
.B1(n_238),
.B2(n_246),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_285),
.A2(n_287),
.B1(n_256),
.B2(n_262),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_217),
.A2(n_229),
.B1(n_242),
.B2(n_232),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_294),
.C(n_296),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_265),
.B(n_228),
.CI(n_227),
.CON(n_292),
.SN(n_292)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_292),
.B(n_308),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_216),
.C(n_252),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_226),
.B1(n_280),
.B2(n_286),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_301),
.B1(n_306),
.B2(n_293),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_226),
.C(n_269),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_263),
.C(n_287),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_286),
.B1(n_285),
.B2(n_277),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_260),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_256),
.C(n_278),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_272),
.A2(n_259),
.B(n_283),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_306),
.A2(n_288),
.B(n_305),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_268),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_303),
.C(n_292),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_301),
.B(n_295),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_296),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_320),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_299),
.B1(n_294),
.B2(n_308),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_310),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_309),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_298),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_313),
.C(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_302),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_330),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_298),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_334),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_314),
.C(n_322),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_335),
.C(n_336),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_320),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_326),
.C(n_312),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_319),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_321),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.C(n_329),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_332),
.C(n_339),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_331),
.A2(n_333),
.B1(n_334),
.B2(n_330),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_342),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_344),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_346),
.B(n_342),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_347),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_340),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_339),
.C(n_343),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_341),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_341),
.Y(n_352)
);


endmodule