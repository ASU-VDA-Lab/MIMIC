module fake_jpeg_3586_n_73 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx9p33_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_10),
.B1(n_19),
.B2(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_23),
.B(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_29),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_32),
.B(n_23),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_43),
.B1(n_34),
.B2(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_58),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_13),
.C(n_17),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_59),
.C(n_51),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_12),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_62),
.C(n_57),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_48),
.C(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_60),
.B2(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_61),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_67),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_56),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_6),
.C(n_9),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_16),
.B(n_20),
.Y(n_73)
);


endmodule