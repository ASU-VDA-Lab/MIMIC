module fake_jpeg_22823_n_48 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_48);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_48;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_11),
.B1(n_19),
.B2(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_23),
.B1(n_1),
.B2(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_23),
.B1(n_24),
.B2(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_4),
.B2(n_6),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_38),
.B1(n_32),
.B2(n_34),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_41),
.B(n_22),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_43),
.C(n_8),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_7),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_9),
.B(n_10),
.Y(n_47)
);

OAI321xp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C(n_17),
.Y(n_48)
);


endmodule