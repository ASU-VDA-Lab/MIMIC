module fake_netlist_5_2299_n_1385 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1385);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1385;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1043;
wire n_486;
wire n_614;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_700;
wire n_1237;
wire n_573;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1184;
wire n_1011;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_252),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_311),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_357),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_168),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_258),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_92),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_118),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_135),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_352),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_361),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_150),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_1),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_94),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_189),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_369),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_124),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_31),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_362),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_128),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_33),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_77),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_20),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_363),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_200),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_148),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_44),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_183),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_315),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_164),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_125),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_109),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_228),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_226),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_91),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_121),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_99),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_222),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_37),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_55),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_197),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_264),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_251),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_54),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_146),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_173),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_131),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_195),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_106),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_271),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_249),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_265),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_72),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_219),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_266),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_38),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_140),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_184),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_160),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_13),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_40),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_203),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_290),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_263),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_333),
.B(n_49),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_136),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_289),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_229),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_245),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_67),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_167),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_321),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_151),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_114),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_256),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_86),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_364),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_126),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_270),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_192),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_161),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_247),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_38),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_172),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_181),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_346),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_304),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_141),
.B(n_239),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_77),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_227),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_314),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_13),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_24),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_207),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_158),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_72),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_351),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_302),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_113),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_157),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_62),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_205),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_138),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g479 ( 
.A(n_83),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_312),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_257),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_325),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_74),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_66),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_293),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_331),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_253),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_277),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_82),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_287),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_186),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_0),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_95),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_89),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_65),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_210),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_342),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_370),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_108),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_246),
.B(n_334),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_137),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_50),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_238),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_56),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_117),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_116),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_358),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_3),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_340),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_154),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_100),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_102),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_335),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_185),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_82),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_115),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_323),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_230),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_215),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_345),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_63),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_43),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_310),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_243),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_176),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_188),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_103),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_144),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_46),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_259),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_159),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_61),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_182),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_142),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_44),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_371),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_244),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_42),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_119),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_234),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_139),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_286),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_224),
.Y(n_543)
);

BUFx5_ASAP7_75t_L g544 ( 
.A(n_187),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_255),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_177),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_11),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_317),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_278),
.Y(n_549)
);

AOI22x1_ASAP7_75t_SL g550 ( 
.A1(n_476),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_419),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_372),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_475),
.B(n_4),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_479),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_375),
.A2(n_5),
.B(n_6),
.Y(n_556)
);

BUFx12f_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_479),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_453),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_414),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_437),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_450),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_469),
.Y(n_566)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_531),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_479),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_479),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_515),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_544),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_499),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_391),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_433),
.A2(n_85),
.B(n_84),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_483),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_395),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_508),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_396),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_398),
.B(n_8),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_447),
.A2(n_88),
.B(n_87),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_401),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_413),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_428),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_544),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_544),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_373),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_407),
.B(n_9),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_464),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_540),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_492),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_409),
.B(n_10),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_509),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_544),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_504),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_427),
.B(n_11),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_439),
.B(n_12),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_509),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_12),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_374),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_526),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_535),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_526),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_376),
.Y(n_607)
);

INVx6_ASAP7_75t_L g608 ( 
.A(n_526),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_452),
.B(n_14),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_542),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_440),
.B(n_14),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_542),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_544),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_542),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_485),
.B(n_15),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_377),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_378),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_379),
.Y(n_618)
);

AOI22x1_ASAP7_75t_SL g619 ( 
.A1(n_435),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_444),
.B(n_16),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_385),
.B(n_17),
.Y(n_621)
);

NOR2x1_ASAP7_75t_L g622 ( 
.A(n_463),
.B(n_18),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_454),
.B(n_18),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_384),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_386),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_389),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_390),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_510),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_553),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_566),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_SL g632 ( 
.A(n_611),
.B(n_436),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_599),
.B(n_512),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_577),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_587),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_602),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_573),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_R g638 ( 
.A(n_592),
.B(n_556),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_583),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_557),
.Y(n_640)
);

INVxp33_ASAP7_75t_SL g641 ( 
.A(n_580),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_607),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_590),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_563),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_608),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_551),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_564),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_567),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_567),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_560),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_618),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_611),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_560),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_608),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_570),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_570),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_572),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_R g658 ( 
.A(n_624),
.B(n_380),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_578),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_578),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_589),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_559),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_626),
.B(n_405),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_589),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_597),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_597),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_621),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_616),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_576),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_R g670 ( 
.A(n_627),
.B(n_423),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_R g671 ( 
.A(n_556),
.B(n_445),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_617),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_625),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_565),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_629),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_642),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_659),
.B(n_661),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_641),
.A2(n_580),
.B1(n_620),
.B2(n_593),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_630),
.B(n_588),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_635),
.B(n_588),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_651),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_656),
.B(n_615),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_646),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_662),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_658),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_636),
.B(n_593),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_650),
.B(n_598),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_653),
.B(n_598),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_674),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_643),
.B(n_430),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_669),
.Y(n_692)
);

AO221x1_ASAP7_75t_L g693 ( 
.A1(n_671),
.A2(n_561),
.B1(n_406),
.B2(n_408),
.C(n_402),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_638),
.B(n_620),
.C(n_609),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_645),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_654),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_632),
.B(n_609),
.C(n_601),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_633),
.B(n_612),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_633),
.B(n_612),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_664),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_668),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_657),
.B(n_614),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_672),
.B(n_601),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_673),
.Y(n_704)
);

AO221x1_ASAP7_75t_L g705 ( 
.A1(n_671),
.A2(n_561),
.B1(n_412),
.B2(n_416),
.C(n_411),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_SL g706 ( 
.A(n_648),
.B(n_565),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_649),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_631),
.B(n_455),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_663),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_652),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_647),
.B(n_615),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_670),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_634),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_667),
.B(n_554),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_655),
.B(n_628),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_660),
.B(n_552),
.C(n_622),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_640),
.B(n_554),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_637),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_665),
.B(n_562),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_639),
.B(n_623),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_666),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_642),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_641),
.B(n_623),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_629),
.B(n_628),
.Y(n_725)
);

BUFx6f_ASAP7_75t_SL g726 ( 
.A(n_642),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_629),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_658),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_642),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_629),
.B(n_565),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_659),
.B(n_562),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_658),
.Y(n_732)
);

AO221x1_ASAP7_75t_L g733 ( 
.A1(n_671),
.A2(n_418),
.B1(n_421),
.B2(n_417),
.C(n_397),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_659),
.B(n_596),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_708),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_730),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_681),
.B(n_687),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_703),
.B(n_422),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_680),
.B(n_459),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_675),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_724),
.B(n_424),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_688),
.B(n_496),
.Y(n_742)
);

XNOR2xp5_ASAP7_75t_L g743 ( 
.A(n_709),
.B(n_501),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_727),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_720),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_514),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_712),
.B(n_441),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_694),
.B(n_443),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_684),
.Y(n_749)
);

BUFx6f_ASAP7_75t_SL g750 ( 
.A(n_719),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_685),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_713),
.B(n_520),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_694),
.B(n_451),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_679),
.A2(n_584),
.B(n_591),
.C(n_582),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_697),
.A2(n_575),
.B1(n_400),
.B2(n_410),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_722),
.B(n_731),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_SL g757 ( 
.A(n_717),
.B(n_467),
.C(n_458),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_733),
.A2(n_456),
.B1(n_381),
.B2(n_383),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_710),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_683),
.A2(n_581),
.B(n_574),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_728),
.B(n_604),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_710),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_710),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_711),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_678),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_693),
.A2(n_524),
.B1(n_525),
.B2(n_523),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_686),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_732),
.B(n_605),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_700),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_676),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_702),
.B(n_472),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_692),
.B(n_575),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_716),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_715),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_701),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_695),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_704),
.B(n_468),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_473),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_682),
.B(n_471),
.Y(n_779)
);

AND2x2_ASAP7_75t_SL g780 ( 
.A(n_691),
.B(n_478),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_696),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_676),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_723),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_690),
.B(n_382),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_729),
.B(n_481),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_725),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_721),
.B(n_484),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_718),
.Y(n_788)
);

OAI21xp33_ASAP7_75t_L g789 ( 
.A1(n_706),
.A2(n_495),
.B(n_489),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_705),
.A2(n_517),
.B1(n_530),
.B2(n_518),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_698),
.A2(n_534),
.B1(n_541),
.B2(n_539),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_726),
.A2(n_388),
.B1(n_392),
.B2(n_387),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_707),
.B(n_393),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_726),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_699),
.A2(n_403),
.B1(n_404),
.B2(n_399),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_714),
.B(n_522),
.C(n_521),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_698),
.A2(n_558),
.B(n_555),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_675),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_730),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_710),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_SL g801 ( 
.A1(n_717),
.A2(n_538),
.B1(n_547),
.B2(n_532),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_681),
.B(n_546),
.Y(n_802)
);

BUFx4f_ASAP7_75t_L g803 ( 
.A(n_710),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_681),
.B(n_548),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_681),
.B(n_415),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_734),
.B(n_420),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_717),
.A2(n_550),
.B1(n_619),
.B2(n_426),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_681),
.B(n_425),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_677),
.B(n_500),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_676),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_730),
.Y(n_811)
);

OR2x6_ASAP7_75t_SL g812 ( 
.A(n_717),
.B(n_429),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_720),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_710),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_730),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_710),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_681),
.B(n_432),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_434),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_720),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_675),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_730),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_720),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_681),
.B(n_438),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_676),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_737),
.B(n_442),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_739),
.A2(n_448),
.B1(n_457),
.B2(n_446),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_746),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_827)
);

OAI22x1_ASAP7_75t_L g828 ( 
.A1(n_743),
.A2(n_466),
.B1(n_470),
.B2(n_465),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_768),
.B(n_474),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_748),
.A2(n_569),
.B(n_571),
.C(n_568),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_753),
.A2(n_585),
.B(n_586),
.C(n_579),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_802),
.B(n_477),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_804),
.B(n_480),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_744),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_R g835 ( 
.A(n_757),
.B(n_482),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_738),
.A2(n_487),
.B1(n_488),
.B2(n_486),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_742),
.B(n_490),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_755),
.A2(n_613),
.B(n_595),
.C(n_493),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_798),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_786),
.A2(n_600),
.B(n_594),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_805),
.A2(n_808),
.B(n_823),
.C(n_817),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_741),
.B(n_491),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_752),
.A2(n_497),
.B1(n_498),
.B2(n_494),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_800),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_781),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_773),
.B(n_767),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_803),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_745),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_800),
.B(n_90),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_736),
.B(n_503),
.Y(n_851)
);

O2A1O1Ixp5_ASAP7_75t_L g852 ( 
.A1(n_760),
.A2(n_506),
.B(n_507),
.C(n_505),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_819),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_759),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_754),
.A2(n_513),
.B(n_516),
.C(n_511),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_774),
.A2(n_528),
.B1(n_533),
.B2(n_527),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_766),
.A2(n_537),
.B1(n_543),
.B2(n_536),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_787),
.A2(n_549),
.B(n_545),
.C(n_603),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_803),
.B(n_606),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_763),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_816),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_777),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_756),
.B(n_19),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_747),
.A2(n_610),
.B(n_606),
.C(n_21),
.Y(n_864)
);

OR2x6_ASAP7_75t_SL g865 ( 
.A(n_772),
.B(n_19),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_751),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_750),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_783),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_765),
.B(n_20),
.C(n_21),
.Y(n_869)
);

CKINVDCx8_ASAP7_75t_R g870 ( 
.A(n_735),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_799),
.B(n_22),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_790),
.A2(n_96),
.B1(n_97),
.B2(n_93),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_811),
.B(n_22),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_815),
.B(n_23),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_821),
.B(n_23),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_814),
.B(n_98),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_SL g877 ( 
.A(n_807),
.B(n_24),
.C(n_25),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_813),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_749),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_814),
.B(n_25),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_769),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_780),
.B(n_101),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_778),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_775),
.B(n_104),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_764),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_R g886 ( 
.A(n_750),
.B(n_105),
.Y(n_886)
);

OA22x2_ASAP7_75t_L g887 ( 
.A1(n_801),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_770),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_788),
.B(n_29),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_806),
.B(n_29),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_761),
.B(n_107),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_794),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_812),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_818),
.B(n_32),
.Y(n_895)
);

AND2x6_ASAP7_75t_L g896 ( 
.A(n_758),
.B(n_110),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_818),
.B(n_33),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_776),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_771),
.B(n_34),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_797),
.A2(n_112),
.B(n_111),
.Y(n_900)
);

BUFx2_ASAP7_75t_SL g901 ( 
.A(n_810),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_779),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_785),
.A2(n_39),
.B(n_36),
.C(n_37),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_782),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_810),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_809),
.B(n_824),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_SL g907 ( 
.A1(n_784),
.A2(n_41),
.B(n_42),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_793),
.A2(n_46),
.B(n_43),
.C(n_45),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_810),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_809),
.B(n_824),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_789),
.A2(n_48),
.B(n_45),
.C(n_47),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_796),
.B(n_47),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_792),
.B(n_48),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_795),
.B(n_50),
.Y(n_914)
);

INVx3_ASAP7_75t_SL g915 ( 
.A(n_791),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_739),
.B(n_51),
.Y(n_916)
);

CKINVDCx14_ASAP7_75t_R g917 ( 
.A(n_743),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_740),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_762),
.B(n_120),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_737),
.B(n_52),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_770),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_768),
.B(n_52),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_740),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_739),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_800),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_748),
.A2(n_123),
.B(n_122),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_745),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_737),
.B(n_53),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_740),
.Y(n_929)
);

BUFx8_ASAP7_75t_L g930 ( 
.A(n_750),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_748),
.A2(n_129),
.B(n_127),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_800),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_803),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_737),
.B(n_56),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_759),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_737),
.B(n_57),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_739),
.B(n_58),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_739),
.A2(n_132),
.B1(n_133),
.B2(n_130),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_737),
.B(n_59),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_737),
.B(n_60),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_768),
.B(n_60),
.Y(n_941)
);

NOR2x1_ASAP7_75t_L g942 ( 
.A(n_800),
.B(n_134),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_756),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_822),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_745),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_737),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_800),
.B(n_143),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_737),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_737),
.A2(n_68),
.B(n_64),
.C(n_67),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_745),
.B(n_68),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_739),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_762),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_SL g953 ( 
.A(n_762),
.B(n_69),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_759),
.Y(n_954)
);

BUFx8_ASAP7_75t_L g955 ( 
.A(n_750),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_768),
.B(n_70),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_737),
.A2(n_74),
.B(n_71),
.C(n_73),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_739),
.A2(n_147),
.B1(n_149),
.B2(n_145),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_762),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_957),
.B(n_73),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_935),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_841),
.A2(n_153),
.B(n_152),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_881),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_829),
.B(n_75),
.Y(n_965)
);

CKINVDCx6p67_ASAP7_75t_R g966 ( 
.A(n_954),
.Y(n_966)
);

AO21x2_ASAP7_75t_L g967 ( 
.A1(n_926),
.A2(n_156),
.B(n_155),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_860),
.B(n_861),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_839),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_847),
.B(n_922),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_852),
.A2(n_163),
.B(n_162),
.Y(n_971)
);

AOI22x1_ASAP7_75t_L g972 ( 
.A1(n_931),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_860),
.B(n_861),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_846),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_868),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_927),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_845),
.B(n_925),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_861),
.B(n_165),
.Y(n_978)
);

AO21x1_ASAP7_75t_L g979 ( 
.A1(n_916),
.A2(n_76),
.B(n_78),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_854),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_848),
.B(n_842),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_918),
.Y(n_982)
);

AO21x2_ASAP7_75t_L g983 ( 
.A1(n_900),
.A2(n_169),
.B(n_166),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_929),
.Y(n_984)
);

BUFx2_ASAP7_75t_SL g985 ( 
.A(n_842),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_945),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_890),
.B(n_79),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_932),
.B(n_170),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_955),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_952),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_930),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_941),
.B(n_956),
.Y(n_992)
);

NOR2x1_ASAP7_75t_L g993 ( 
.A(n_952),
.B(n_171),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_898),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_937),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_930),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_906),
.B(n_174),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_952),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_885),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_920),
.B(n_80),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_928),
.B(n_81),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_878),
.Y(n_1002)
);

BUFx8_ASAP7_75t_L g1003 ( 
.A(n_894),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_960),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_934),
.A2(n_175),
.B(n_178),
.Y(n_1005)
);

BUFx2_ASAP7_75t_SL g1006 ( 
.A(n_960),
.Y(n_1006)
);

BUFx2_ASAP7_75t_SL g1007 ( 
.A(n_850),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_867),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_862),
.B(n_179),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_853),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_905),
.B(n_180),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_943),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_936),
.B(n_368),
.Y(n_1013)
);

INVx8_ASAP7_75t_L g1014 ( 
.A(n_888),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_849),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_866),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_870),
.Y(n_1017)
);

INVx3_ASAP7_75t_SL g1018 ( 
.A(n_933),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_888),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_834),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_850),
.Y(n_1021)
);

AOI22x1_ASAP7_75t_L g1022 ( 
.A1(n_923),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_913),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_871),
.A2(n_194),
.B(n_196),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_863),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_939),
.A2(n_198),
.B(n_199),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_940),
.A2(n_201),
.B(n_202),
.Y(n_1027)
);

AO21x2_ASAP7_75t_L g1028 ( 
.A1(n_858),
.A2(n_204),
.B(n_206),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_950),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_944),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_910),
.A2(n_208),
.B(n_209),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_899),
.A2(n_211),
.B(n_212),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_876),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_896),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_947),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_904),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_909),
.Y(n_1037)
);

BUFx4f_ASAP7_75t_SL g1038 ( 
.A(n_884),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_947),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_879),
.Y(n_1040)
);

INVx6_ASAP7_75t_L g1041 ( 
.A(n_895),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_R g1042 ( 
.A(n_901),
.B(n_217),
.Y(n_1042)
);

AO21x2_ASAP7_75t_L g1043 ( 
.A1(n_882),
.A2(n_218),
.B(n_220),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_832),
.A2(n_221),
.B(n_223),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_915),
.B(n_225),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_SL g1046 ( 
.A(n_896),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_893),
.Y(n_1047)
);

AO21x2_ASAP7_75t_L g1048 ( 
.A1(n_833),
.A2(n_231),
.B(n_232),
.Y(n_1048)
);

AO21x2_ASAP7_75t_L g1049 ( 
.A1(n_843),
.A2(n_233),
.B(n_235),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_838),
.A2(n_236),
.B(n_237),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_825),
.B(n_240),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_830),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_831),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_873),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_897),
.Y(n_1055)
);

BUFx5_ASAP7_75t_L g1056 ( 
.A(n_896),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_917),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_921),
.B(n_241),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_874),
.B(n_242),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_875),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_835),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_887),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_953),
.B(n_942),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_828),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_919),
.B(n_248),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_908),
.B(n_250),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_911),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_865),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_891),
.B(n_254),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_886),
.Y(n_1071)
);

OA21x2_ASAP7_75t_L g1072 ( 
.A1(n_851),
.A2(n_260),
.B(n_261),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_914),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_864),
.Y(n_1074)
);

BUFx2_ASAP7_75t_R g1075 ( 
.A(n_859),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_880),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_907),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_946),
.Y(n_1078)
);

BUFx2_ASAP7_75t_R g1079 ( 
.A(n_877),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_912),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_892),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_837),
.B(n_262),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_840),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_924),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_856),
.Y(n_1085)
);

CKINVDCx8_ASAP7_75t_R g1086 ( 
.A(n_958),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_949),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_855),
.A2(n_267),
.B(n_268),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_872),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_869),
.Y(n_1090)
);

BUFx5_ASAP7_75t_L g1091 ( 
.A(n_938),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1016),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_974),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1052),
.A2(n_1053),
.B(n_1013),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1021),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_SL g1096 ( 
.A1(n_1023),
.A2(n_959),
.B1(n_826),
.B2(n_827),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_975),
.Y(n_1097)
);

INVx6_ASAP7_75t_L g1098 ( 
.A(n_998),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_964),
.Y(n_1099)
);

OAI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1080),
.A2(n_844),
.B1(n_836),
.B2(n_948),
.Y(n_1100)
);

OA21x2_ASAP7_75t_L g1101 ( 
.A1(n_963),
.A2(n_902),
.B(n_951),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1054),
.A2(n_857),
.B(n_903),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_999),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_998),
.B(n_883),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1021),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_986),
.Y(n_1106)
);

OAI21xp33_ASAP7_75t_SL g1107 ( 
.A1(n_1082),
.A2(n_269),
.B(n_272),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_962),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_1036),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1084),
.A2(n_1023),
.B1(n_987),
.B2(n_1091),
.Y(n_1110)
);

CKINVDCx11_ASAP7_75t_R g1111 ( 
.A(n_989),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_970),
.B(n_992),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_1057),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1040),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_976),
.B(n_273),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1055),
.B(n_274),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_968),
.Y(n_1117)
);

INVx6_ASAP7_75t_L g1118 ( 
.A(n_973),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1081),
.A2(n_275),
.B1(n_276),
.B2(n_279),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1033),
.B(n_367),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1020),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1054),
.B(n_280),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1076),
.B(n_281),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_969),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_982),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_1030),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1010),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_984),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1084),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_994),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_1010),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1062),
.B(n_285),
.Y(n_1132)
);

BUFx8_ASAP7_75t_SL g1133 ( 
.A(n_991),
.Y(n_1133)
);

CKINVDCx14_ASAP7_75t_R g1134 ( 
.A(n_996),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1091),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1091),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1047),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1008),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_980),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1037),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1069),
.B(n_365),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_SL g1142 ( 
.A1(n_1046),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1073),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1074),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_981),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1074),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1091),
.A2(n_301),
.B1(n_303),
.B2(n_305),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_990),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1038),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1067),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_961),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1035),
.B(n_309),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1007),
.A2(n_1060),
.B1(n_1089),
.B2(n_1085),
.Y(n_1153)
);

AO22x1_ASAP7_75t_L g1154 ( 
.A1(n_1050),
.A2(n_313),
.B1(n_316),
.B2(n_318),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1083),
.Y(n_1155)
);

NOR2xp67_ASAP7_75t_SL g1156 ( 
.A(n_1071),
.B(n_322),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1015),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_SL g1158 ( 
.A1(n_965),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1078),
.Y(n_1159)
);

BUFx2_ASAP7_75t_R g1160 ( 
.A(n_1018),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1060),
.B(n_328),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1045),
.B(n_329),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_1014),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1002),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1014),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1071),
.B(n_330),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_977),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_SL g1168 ( 
.A1(n_1005),
.A2(n_332),
.B(n_336),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1053),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1068),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1087),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_1017),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1077),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1058),
.Y(n_1174)
);

BUFx2_ASAP7_75t_R g1175 ( 
.A(n_1061),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1000),
.B(n_347),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1087),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1001),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_997),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1025),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_990),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_997),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_978),
.B(n_353),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_972),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_966),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1019),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1003),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1019),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1015),
.B(n_359),
.Y(n_1189)
);

CKINVDCx11_ASAP7_75t_R g1190 ( 
.A(n_1029),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1098),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1112),
.B(n_1064),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_R g1193 ( 
.A(n_1113),
.B(n_1071),
.Y(n_1193)
);

AO32x2_ASAP7_75t_L g1194 ( 
.A1(n_1153),
.A2(n_979),
.A3(n_972),
.B1(n_995),
.B2(n_1086),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1127),
.B(n_1051),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1102),
.A2(n_1026),
.B(n_1027),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1178),
.B(n_1012),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1099),
.Y(n_1198)
);

AND2x4_ASAP7_75t_SL g1199 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1100),
.A2(n_971),
.B(n_1066),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1151),
.B(n_978),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1096),
.B(n_1034),
.C(n_1063),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1143),
.B(n_1059),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1137),
.B(n_1189),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_R g1205 ( 
.A(n_1172),
.B(n_1039),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1157),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1111),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1110),
.B(n_1009),
.C(n_1031),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1184),
.B(n_1066),
.C(n_1022),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1109),
.B(n_1131),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1126),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1183),
.B(n_1041),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1159),
.B(n_1059),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1123),
.B(n_1041),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1133),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1092),
.B(n_1171),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1101),
.A2(n_1090),
.B1(n_1056),
.B2(n_967),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1174),
.B(n_1090),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_SL g1219 ( 
.A(n_1119),
.B(n_1070),
.C(n_1011),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1116),
.B(n_1079),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1093),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1103),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1160),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1132),
.B(n_1006),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1139),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1140),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1121),
.B(n_985),
.Y(n_1227)
);

NOR3xp33_ASAP7_75t_SL g1228 ( 
.A(n_1141),
.B(n_1003),
.C(n_1075),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1163),
.B(n_1004),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_1164),
.B(n_1004),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1180),
.B(n_1173),
.C(n_1158),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1162),
.A2(n_1056),
.B1(n_1043),
.B2(n_983),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1097),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1138),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1108),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1117),
.B(n_1056),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_1122),
.A2(n_1042),
.B(n_1065),
.C(n_993),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1106),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_1187),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1134),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_R g1241 ( 
.A(n_1185),
.B(n_1004),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1179),
.A2(n_1182),
.B1(n_1144),
.B2(n_1146),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1177),
.A2(n_1114),
.B1(n_1104),
.B2(n_1145),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1118),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1169),
.B(n_988),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1190),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1175),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1124),
.B(n_1125),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1165),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1128),
.B(n_1044),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_R g1251 ( 
.A(n_1148),
.B(n_1181),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_SL g1252 ( 
.A(n_1166),
.B(n_1024),
.C(n_1049),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1170),
.A2(n_1028),
.B1(n_1088),
.B2(n_1072),
.Y(n_1253)
);

CKINVDCx16_ASAP7_75t_R g1254 ( 
.A(n_1115),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_1120),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1130),
.B(n_1048),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1152),
.B(n_1032),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1233),
.B(n_1155),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1210),
.B(n_1150),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1221),
.B(n_1094),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1226),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1250),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1238),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1206),
.B(n_1176),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1223),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1248),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1231),
.A2(n_1168),
.B1(n_1149),
.B2(n_1136),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1198),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1257),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1204),
.B(n_1161),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1216),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1256),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1242),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1236),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1213),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1202),
.A2(n_1135),
.B1(n_1147),
.B2(n_1142),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1191),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1227),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1200),
.B(n_1186),
.Y(n_1279)
);

CKINVDCx6p67_ASAP7_75t_R g1280 ( 
.A(n_1239),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1195),
.B(n_1243),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1194),
.B(n_1105),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1201),
.B(n_1255),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1194),
.B(n_1095),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1197),
.B(n_1152),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1254),
.B(n_1167),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1222),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1203),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1191),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1217),
.B(n_1188),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1196),
.B(n_1154),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1291),
.B(n_1245),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1291),
.B(n_1209),
.C(n_1154),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1269),
.B(n_1192),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1275),
.B(n_1225),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1263),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1262),
.B(n_1211),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1260),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1258),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1275),
.B(n_1218),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1269),
.B(n_1278),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1281),
.B(n_1208),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1271),
.B(n_1224),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1261),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1287),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1272),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1262),
.B(n_1252),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1259),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1265),
.B(n_1207),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1288),
.B(n_1232),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1259),
.Y(n_1311)
);

OAI211xp5_ASAP7_75t_L g1312 ( 
.A1(n_1267),
.A2(n_1107),
.B(n_1129),
.C(n_1253),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1266),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1292),
.B(n_1281),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1299),
.B(n_1282),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1298),
.Y(n_1316)
);

NOR2xp67_ASAP7_75t_L g1317 ( 
.A(n_1304),
.B(n_1268),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1298),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1303),
.B(n_1287),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1301),
.B(n_1280),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1294),
.B(n_1280),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1296),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1295),
.B(n_1274),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1302),
.B(n_1306),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1296),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1302),
.B(n_1274),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1300),
.B(n_1292),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1293),
.B(n_1288),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1328),
.A2(n_1312),
.B1(n_1276),
.B2(n_1310),
.Y(n_1329)
);

OAI221xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1324),
.A2(n_1264),
.B1(n_1285),
.B2(n_1297),
.C(n_1270),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1326),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1316),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1322),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1316),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1328),
.A2(n_1286),
.B1(n_1273),
.B2(n_1283),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1327),
.B(n_1313),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1319),
.B(n_1308),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1317),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1318),
.Y(n_1339)
);

NAND4xp25_ASAP7_75t_L g1340 ( 
.A(n_1314),
.B(n_1220),
.C(n_1309),
.D(n_1310),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1314),
.B(n_1311),
.Y(n_1341)
);

OAI321xp33_ASAP7_75t_L g1342 ( 
.A1(n_1323),
.A2(n_1307),
.A3(n_1279),
.B1(n_1219),
.B2(n_1284),
.C(n_1290),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1318),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1331),
.B(n_1315),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1341),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1332),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1329),
.A2(n_1320),
.B(n_1321),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1335),
.B(n_1305),
.C(n_1307),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1334),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1333),
.B(n_1325),
.Y(n_1350)
);

OAI31xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1340),
.A2(n_1338),
.A3(n_1342),
.B(n_1330),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1345),
.B(n_1336),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1346),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1344),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1350),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1348),
.B(n_1337),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1355),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1352),
.B(n_1351),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1356),
.B(n_1351),
.C(n_1340),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_SL g1360 ( 
.A(n_1354),
.B(n_1347),
.C(n_1193),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1353),
.B(n_1246),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1352),
.B(n_1215),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1359),
.B(n_1263),
.Y(n_1363)
);

AOI211xp5_ASAP7_75t_L g1364 ( 
.A1(n_1358),
.A2(n_1247),
.B(n_1237),
.C(n_1349),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1357),
.Y(n_1365)
);

NAND4xp25_ASAP7_75t_SL g1366 ( 
.A(n_1363),
.B(n_1364),
.C(n_1365),
.D(n_1360),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1363),
.A2(n_1362),
.B(n_1361),
.Y(n_1367)
);

NOR3xp33_ASAP7_75t_L g1368 ( 
.A(n_1366),
.B(n_1240),
.C(n_1265),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1368),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1369),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1369),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1370),
.A2(n_1234),
.B1(n_1235),
.B2(n_1249),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1371),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1373),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1372),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1374),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_L g1377 ( 
.A1(n_1375),
.A2(n_1367),
.B(n_1191),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1376),
.A2(n_1277),
.B1(n_1289),
.B2(n_1305),
.Y(n_1378)
);

OAI22x1_ASAP7_75t_SL g1379 ( 
.A1(n_1377),
.A2(n_1205),
.B1(n_1241),
.B2(n_1228),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1378),
.B(n_1339),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_SL g1381 ( 
.A(n_1379),
.B(n_1277),
.Y(n_1381)
);

AOI222xp33_ASAP7_75t_L g1382 ( 
.A1(n_1380),
.A2(n_1156),
.B1(n_1289),
.B2(n_1343),
.C1(n_1229),
.C2(n_1214),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1381),
.A2(n_1199),
.B1(n_1230),
.B2(n_1244),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1383),
.B(n_1212),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1384),
.A2(n_1382),
.B1(n_1230),
.B2(n_1251),
.Y(n_1385)
);


endmodule