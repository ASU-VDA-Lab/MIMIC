module real_jpeg_30749_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_703, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_703;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_372;
wire n_219;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_635;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_0),
.Y(n_133)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_0),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_0),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_164),
.B1(n_165),
.B2(n_170),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_2),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_2),
.A2(n_164),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_2),
.A2(n_164),
.B1(n_296),
.B2(n_300),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_2),
.A2(n_164),
.B1(n_407),
.B2(n_410),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_3),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_3),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_3),
.A2(n_190),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_3),
.A2(n_190),
.B1(n_376),
.B2(n_379),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_3),
.A2(n_190),
.B1(n_467),
.B2(n_470),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_117),
.B1(n_124),
.B2(n_125),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_124),
.B1(n_150),
.B2(n_155),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_4),
.A2(n_124),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

AO22x1_ASAP7_75t_L g632 ( 
.A1(n_4),
.A2(n_124),
.B1(n_633),
.B2(n_635),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_243),
.B1(n_244),
.B2(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_5),
.A2(n_243),
.B1(n_345),
.B2(n_349),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_5),
.A2(n_243),
.B1(n_438),
.B2(n_441),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_5),
.A2(n_243),
.B1(n_538),
.B2(n_540),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_6),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_6),
.A2(n_81),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_6),
.A2(n_81),
.B1(n_641),
.B2(n_642),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_6),
.A2(n_81),
.B1(n_679),
.B2(n_681),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_7),
.B(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_7),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_7),
.B(n_174),
.Y(n_412)
);

OAI32xp33_ASAP7_75t_L g445 ( 
.A1(n_7),
.A2(n_446),
.A3(n_449),
.B1(n_451),
.B2(n_456),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_7),
.A2(n_372),
.B1(n_488),
.B2(n_491),
.Y(n_487)
);

OAI21xp33_ASAP7_75t_L g519 ( 
.A1(n_7),
.A2(n_224),
.B(n_520),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_20),
.B(n_23),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_10),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_11),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_12),
.A2(n_112),
.B1(n_210),
.B2(n_213),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_12),
.A2(n_112),
.B1(n_333),
.B2(n_336),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_12),
.A2(n_112),
.B1(n_321),
.B2(n_610),
.Y(n_609)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_16),
.A2(n_275),
.B1(n_276),
.B2(n_282),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_16),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_16),
.A2(n_275),
.B1(n_387),
.B2(n_393),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_16),
.A2(n_275),
.B1(n_494),
.B2(n_496),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_16),
.A2(n_275),
.B1(n_508),
.B2(n_512),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_17),
.Y(n_111)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_18),
.A2(n_64),
.B1(n_219),
.B2(n_222),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_18),
.A2(n_64),
.B1(n_619),
.B2(n_622),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_18),
.A2(n_64),
.B1(n_660),
.B2(n_663),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_596),
.B(n_687),
.C(n_697),
.D(n_700),
.Y(n_25)
);

NAND2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_426),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_351),
.B(n_422),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_29),
.B(n_593),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_250),
.B(n_301),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g424 ( 
.A(n_30),
.B(n_250),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_30),
.B(n_250),
.Y(n_425)
);

XOR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_206),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_128),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_32),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_87),
.B(n_127),
.Y(n_32)
);

NAND2x1_ASAP7_75t_L g127 ( 
.A(n_33),
.B(n_87),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_62),
.B1(n_75),
.B2(n_85),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_34),
.A2(n_375),
.B1(n_381),
.B2(n_382),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_34),
.B(n_570),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_34),
.A2(n_85),
.B1(n_375),
.B2(n_580),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g615 ( 
.A1(n_34),
.A2(n_75),
.B(n_85),
.Y(n_615)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_35),
.A2(n_63),
.B1(n_149),
.B2(n_158),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_35),
.A2(n_149),
.B1(n_158),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_35),
.A2(n_158),
.B1(n_209),
.B2(n_295),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_SL g436 ( 
.A1(n_35),
.A2(n_437),
.B(n_443),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_35),
.A2(n_158),
.B1(n_437),
.B2(n_493),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_50),
.Y(n_35)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

OAI22x1_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_44),
.B2(n_47),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_38),
.Y(n_514)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_43),
.Y(n_555)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_45),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_47),
.Y(n_471)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_49),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_49),
.Y(n_469)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_49),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_50)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_51),
.Y(n_450)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_52),
.Y(n_380)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_58),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_58),
.Y(n_442)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_69),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g495 ( 
.A(n_68),
.Y(n_495)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_73),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_74),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g561 ( 
.A(n_74),
.Y(n_561)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_80),
.Y(n_212)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_80),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_80),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_85),
.B(n_375),
.Y(n_443)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_86),
.B(n_372),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_106),
.B1(n_115),
.B2(n_116),
.Y(n_87)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_88),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_88),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_88),
.B(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_88),
.A2(n_116),
.B1(n_385),
.B2(n_618),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_88),
.A2(n_115),
.B1(n_618),
.B2(n_640),
.Y(n_639)
);

OAI21xp33_ASAP7_75t_SL g657 ( 
.A1(n_88),
.A2(n_115),
.B(n_640),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_92),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_97),
.B1(n_101),
.B2(n_105),
.Y(n_96)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_97),
.Y(n_349)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_99),
.Y(n_622)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_106),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_109),
.Y(n_265)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_110),
.Y(n_235)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

BUFx4f_ASAP7_75t_L g313 ( 
.A(n_113),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_114),
.Y(n_232)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_114),
.Y(n_348)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_114),
.Y(n_621)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_115),
.Y(n_236)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_115),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_115),
.B(n_263),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_115),
.B(n_386),
.Y(n_415)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_122),
.Y(n_394)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_122),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_123),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_123),
.Y(n_392)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_127),
.B(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_127),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_128),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_159),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_129),
.A2(n_203),
.B(n_604),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_148),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_130),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B(n_141),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_131),
.Y(n_464)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_134),
.A2(n_141),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_134),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_134),
.A2(n_227),
.B1(n_287),
.B2(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_134),
.B(n_466),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_134),
.A2(n_292),
.B1(n_535),
.B2(n_536),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_137),
.Y(n_289)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_137),
.Y(n_531)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_140),
.Y(n_517)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_141),
.Y(n_225)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_146),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_147),
.Y(n_335)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_147),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_147),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_148),
.A2(n_202),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_148),
.Y(n_257)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx4f_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_158),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_202),
.B2(n_203),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_161),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_187),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g607 ( 
.A1(n_163),
.A2(n_608),
.B1(n_609),
.B2(n_612),
.Y(n_607)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_171),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_169),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_169),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_174),
.B(n_188),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g273 ( 
.A1(n_174),
.A2(n_194),
.B1(n_242),
.B2(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_174),
.B(n_274),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_174),
.Y(n_612)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_178),
.Y(n_328)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_180),
.Y(n_490)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_184),
.Y(n_325)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_186),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_186),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_187),
.B(n_341),
.Y(n_340)
);

NAND2x1_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_193),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_194),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_194),
.B(n_367),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_194),
.Y(n_608)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_197),
.Y(n_315)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_205),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_205),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_R g599 ( 
.A(n_206),
.B(n_600),
.C(n_601),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_228),
.C(n_238),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_217),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_208),
.B(n_217),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_212),
.Y(n_300)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_218),
.A2(n_224),
.B1(n_286),
.B2(n_291),
.Y(n_285)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_221),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22x1_ASAP7_75t_L g401 ( 
.A1(n_224),
.A2(n_332),
.B1(n_402),
.B2(n_406),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_224),
.A2(n_520),
.B(n_537),
.Y(n_577)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_238),
.B1(n_239),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_237),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_230),
.B1(n_262),
.B2(n_271),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_229),
.A2(n_344),
.B(n_350),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_229),
.A2(n_350),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_240),
.B(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_247),
.Y(n_680)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_258),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_259),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_272),
.C(n_284),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_273),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_262),
.Y(n_418)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_267),
.Y(n_458)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_271),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_271),
.B(n_372),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_279),
.Y(n_636)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_279),
.Y(n_685)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_285),
.B(n_294),
.Y(n_362)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_293),
.Y(n_528)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_295),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_302),
.B(n_304),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.C(n_309),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_339),
.C(n_342),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_SL g358 ( 
.A(n_310),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_329),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_311),
.A2(n_312),
.B1(n_329),
.B2(n_330),
.Y(n_419)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI32xp33_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.A3(n_316),
.B1(n_320),
.B2(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_319),
.Y(n_634)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_319),
.Y(n_662)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_337),
.Y(n_542)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_340),
.B1(n_343),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_357),
.C(n_395),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_353),
.A2(n_594),
.B(n_595),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_357),
.Y(n_594)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.C(n_363),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_358),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_364),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_374),
.C(n_383),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_365),
.B(n_398),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_372),
.B(n_373),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_372),
.B(n_452),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_372),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_372),
.B(n_558),
.Y(n_557)
);

OAI21xp33_ASAP7_75t_SL g570 ( 
.A1(n_372),
.A2(n_557),
.B(n_571),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_383),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_378),
.Y(n_500)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_420),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_396),
.B(n_420),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.C(n_419),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_397),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_400),
.A2(n_419),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_412),
.B1(n_413),
.B2(n_416),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_412),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_412),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_401),
.A2(n_412),
.B1(n_413),
.B2(n_416),
.Y(n_476)
);

INVx3_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_406),
.A2(n_464),
.B(n_465),
.Y(n_463)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_417),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B(n_425),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_592),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_477),
.B(n_590),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_472),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_430),
.B(n_591),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_435),
.C(n_444),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_432),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_435),
.A2(n_436),
.B1(n_444),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_443),
.B(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_463),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_445),
.B(n_463),
.Y(n_484)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_465),
.A2(n_507),
.B(n_515),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_466),
.B(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_501),
.B(n_589),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_479),
.B(n_482),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.C(n_492),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_484),
.B(n_575),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_486),
.B(n_492),
.Y(n_575)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_493),
.Y(n_580)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

OAI321xp33_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_573),
.A3(n_582),
.B1(n_587),
.B2(n_588),
.C(n_703),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_533),
.B(n_572),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_504),
.A2(n_518),
.B(n_532),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_505),
.B(n_506),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_507),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx2_ASAP7_75t_SL g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_519),
.B(n_526),
.Y(n_518)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_529),
.Y(n_526)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_543),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_534),
.B(n_543),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_568),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_544),
.B(n_568),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_545),
.A2(n_556),
.B1(n_562),
.B2(n_567),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_550),
.Y(n_545)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_546),
.Y(n_567)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_565),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_564),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_574),
.B(n_576),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_576),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_577),
.B(n_578),
.C(n_581),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_585),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_578),
.A2(n_579),
.B1(n_581),
.B2(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_581),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_584),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_583),
.B(n_584),
.Y(n_587)
);

NOR3x1_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_651),
.C(n_671),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_598),
.B(n_624),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_602),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_599),
.B(n_602),
.Y(n_696)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_605),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_603),
.B(n_649),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_603),
.B(n_649),
.Y(n_650)
);

INVxp33_ASAP7_75t_L g647 ( 
.A(n_606),
.Y(n_647)
);

XNOR2x1_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_613),
.Y(n_606)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_607),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_607),
.B(n_626),
.C(n_670),
.Y(n_669)
);

AO22x1_ASAP7_75t_SL g631 ( 
.A1(n_608),
.A2(n_609),
.B1(n_612),
.B2(n_632),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_608),
.A2(n_612),
.B1(n_632),
.B2(n_659),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_608),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_608),
.A2(n_612),
.B(n_678),
.Y(n_699)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_612),
.Y(n_676)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_614),
.A2(n_616),
.B(n_623),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_614),
.A2(n_615),
.B1(n_638),
.B2(n_639),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_614),
.B(n_638),
.C(n_655),
.Y(n_654)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_615),
.B(n_617),
.Y(n_623)
);

MAJx2_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_616),
.C(n_627),
.Y(n_626)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_620),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_621),
.Y(n_620)
);

INVx3_ASAP7_75t_SL g641 ( 
.A(n_622),
.Y(n_641)
);

NAND4xp25_ASAP7_75t_L g695 ( 
.A(n_624),
.B(n_652),
.C(n_672),
.D(n_696),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_625),
.B(n_646),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_625),
.B(n_646),
.Y(n_692)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_626),
.B(n_628),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_627),
.B(n_629),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_629),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_637),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_631),
.Y(n_655)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_647),
.A2(n_648),
.B(n_650),
.Y(n_646)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

AOI31xp33_ASAP7_75t_L g691 ( 
.A1(n_652),
.A2(n_672),
.A3(n_692),
.B(n_693),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_653),
.B(n_669),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_653),
.B(n_669),
.Y(n_690)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_654),
.B(n_656),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_654),
.B(n_658),
.C(n_667),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_657),
.A2(n_658),
.B1(n_667),
.B2(n_668),
.Y(n_656)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_657),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_658),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_659),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_662),
.Y(n_661)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_662),
.Y(n_666)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_665),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_672),
.B(n_689),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_673),
.B(n_686),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_673),
.B(n_686),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_673),
.B(n_698),
.Y(n_697)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_673),
.Y(n_701)
);

OA22x2_ASAP7_75t_L g673 ( 
.A1(n_674),
.A2(n_675),
.B1(n_676),
.B2(n_677),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_678),
.Y(n_677)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_680),
.Y(n_679)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_682),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_683),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_684),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_685),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_SL g687 ( 
.A(n_688),
.B(n_691),
.C(n_695),
.Y(n_687)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_690),
.Y(n_689)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_694),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_699),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_699),
.B(n_701),
.Y(n_700)
);


endmodule