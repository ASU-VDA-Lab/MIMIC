module fake_jpeg_30899_n_528 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_58),
.Y(n_124)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_52),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_78),
.Y(n_127)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_17),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_17),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_79),
.B(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g152 ( 
.A(n_93),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_1),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_2),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_41),
.Y(n_136)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_49),
.Y(n_126)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_37),
.B1(n_42),
.B2(n_19),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_119),
.A2(n_134),
.B1(n_56),
.B2(n_57),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_60),
.A2(n_37),
.B1(n_49),
.B2(n_46),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_125),
.A2(n_157),
.B1(n_65),
.B2(n_82),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_138),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_19),
.B1(n_42),
.B2(n_51),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_136),
.B(n_16),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_81),
.B(n_51),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_141),
.B(n_72),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_55),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_70),
.A2(n_50),
.B1(n_20),
.B2(n_21),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_50),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_170),
.B(n_204),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_190),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_127),
.A2(n_31),
.B(n_22),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_173),
.A2(n_222),
.B(n_227),
.C(n_11),
.Y(n_252)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_183),
.A2(n_184),
.B1(n_189),
.B2(n_194),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_59),
.C(n_102),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_186),
.B(n_201),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_31),
.B(n_21),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_187),
.A2(n_219),
.B(n_225),
.Y(n_237)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_140),
.A2(n_103),
.B1(n_91),
.B2(n_90),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_25),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_192),
.A2(n_210),
.B1(n_218),
.B2(n_220),
.Y(n_234)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_77),
.B1(n_76),
.B2(n_22),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_196),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_34),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_202),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_112),
.A2(n_33),
.B1(n_73),
.B2(n_99),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_199),
.A2(n_208),
.B1(n_221),
.B2(n_219),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_211),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_87),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_124),
.B(n_42),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_203),
.B(n_214),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_115),
.B(n_130),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_205),
.Y(n_265)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_161),
.B1(n_163),
.B2(n_135),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_42),
.B1(n_41),
.B2(n_4),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_128),
.A2(n_42),
.B1(n_41),
.B2(n_5),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_150),
.A2(n_41),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_114),
.Y(n_215)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_116),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_216),
.Y(n_269)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_137),
.A2(n_2),
.B(n_3),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_129),
.A2(n_41),
.B1(n_3),
.B2(n_5),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_118),
.A2(n_16),
.B1(n_3),
.B2(n_5),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_151),
.A2(n_2),
.B(n_6),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_146),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_143),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_154),
.A2(n_8),
.B(n_11),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_171),
.B(n_168),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_228),
.B(n_235),
.Y(n_300)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_134),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_232),
.B(n_252),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_170),
.B(n_142),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_233),
.B(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_187),
.B(n_139),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_236),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_133),
.B1(n_117),
.B2(n_166),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_238),
.A2(n_253),
.B1(n_256),
.B2(n_264),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_241),
.A2(n_273),
.B1(n_218),
.B2(n_178),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_204),
.B(n_162),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_201),
.B(n_163),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_258),
.Y(n_276)
);

NAND2x1_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_116),
.Y(n_251)
);

XOR2x1_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_250),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_182),
.A2(n_161),
.B1(n_158),
.B2(n_148),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_217),
.A2(n_153),
.B1(n_14),
.B2(n_16),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_16),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_13),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_268),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_226),
.A2(n_13),
.B1(n_14),
.B2(n_212),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_186),
.B(n_14),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_213),
.A2(n_14),
.B1(n_211),
.B2(n_180),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_271),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_173),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_251),
.B1(n_255),
.B2(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_231),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_278),
.B(n_281),
.Y(n_345)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_240),
.A2(n_221),
.B1(n_188),
.B2(n_193),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_280),
.A2(n_283),
.B1(n_284),
.B2(n_241),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

AOI32xp33_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_196),
.A3(n_185),
.B1(n_174),
.B2(n_198),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_303),
.B(n_234),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_255),
.A2(n_215),
.B1(n_206),
.B2(n_209),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_260),
.A3(n_258),
.B1(n_273),
.B2(n_235),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_177),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_292),
.Y(n_320)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_228),
.B(n_181),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_293),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_191),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_304),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_175),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_302),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_229),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_237),
.A2(n_175),
.B(n_176),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_243),
.B(n_179),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_305),
.B(n_242),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_247),
.B(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_270),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_243),
.B(n_261),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_310),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_267),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_261),
.B(n_252),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_262),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_314),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_229),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_321),
.C(n_341),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_316),
.A2(n_324),
.B(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_344),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_251),
.C(n_270),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_265),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_323),
.B(n_332),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_301),
.A2(n_263),
.B1(n_249),
.B2(n_230),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_232),
.B(n_230),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_257),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_329),
.B(n_334),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_265),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_259),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_249),
.B1(n_246),
.B2(n_263),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_336),
.A2(n_278),
.B1(n_296),
.B2(n_309),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_259),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_340),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_285),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_276),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_284),
.A2(n_249),
.B1(n_254),
.B2(n_262),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_275),
.B(n_292),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_345),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_347),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_348),
.A2(n_361),
.B1(n_344),
.B2(n_328),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_318),
.A2(n_311),
.B1(n_298),
.B2(n_274),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_364),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_378),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_286),
.B(n_303),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_351),
.A2(n_340),
.B(n_322),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_363),
.C(n_365),
.Y(n_386)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_311),
.B1(n_286),
.B2(n_280),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_276),
.C(n_305),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_318),
.A2(n_277),
.B(n_282),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_294),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_316),
.A2(n_303),
.B(n_327),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_366),
.A2(n_322),
.B(n_320),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_300),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_367),
.B(n_369),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_298),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_368),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_326),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_310),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_373),
.C(n_333),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_325),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_371),
.B(n_376),
.Y(n_381)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_330),
.Y(n_372)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_307),
.C(n_299),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_330),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_375),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_346),
.B(n_287),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_335),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_377),
.Y(n_389)
);

XOR2x2_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_317),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_320),
.Y(n_379)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_379),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_352),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_382),
.B(n_384),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_360),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_372),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_387),
.B(n_392),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_333),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_393),
.Y(n_431)
);

AND2x4_ASAP7_75t_SL g391 ( 
.A(n_366),
.B(n_317),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_338),
.C(n_334),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_395),
.C(n_397),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_329),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_335),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_319),
.C(n_328),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_403),
.C(n_378),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_348),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_400),
.B(n_405),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_350),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_374),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_314),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_375),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_406),
.A2(n_355),
.B1(n_368),
.B2(n_364),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_408),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_413),
.B(n_426),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_358),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_415),
.Y(n_441)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_416),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_417),
.B(n_419),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_425),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_420),
.A2(n_349),
.B1(n_361),
.B2(n_362),
.Y(n_456)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_423),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_356),
.C(n_370),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_429),
.C(n_394),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_379),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_358),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_432),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_388),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_428),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_356),
.C(n_368),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_325),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_430),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_383),
.B(n_404),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_380),
.Y(n_448)
);

AOI211xp5_ASAP7_75t_SL g435 ( 
.A1(n_412),
.A2(n_391),
.B(n_398),
.C(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_386),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_417),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_412),
.A2(n_406),
.B1(n_407),
.B2(n_403),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_437),
.A2(n_450),
.B1(n_420),
.B2(n_414),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_429),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_390),
.C(n_393),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_443),
.C(n_445),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_397),
.C(n_401),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_395),
.C(n_402),
.Y(n_445)
);

FAx1_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_391),
.CI(n_407),
.CON(n_446),
.SN(n_446)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_433),
.Y(n_460)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_409),
.A2(n_351),
.B(n_354),
.Y(n_449)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_409),
.A2(n_362),
.B1(n_354),
.B2(n_364),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_456),
.A2(n_402),
.B1(n_427),
.B2(n_421),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_441),
.B(n_411),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_457),
.B(n_463),
.Y(n_488)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_458),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_460),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_439),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_464),
.A2(n_466),
.B1(n_471),
.B2(n_472),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_465),
.A2(n_437),
.B1(n_450),
.B2(n_442),
.Y(n_474)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_470),
.C(n_438),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_455),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_419),
.C(n_424),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_453),
.B(n_434),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_454),
.A2(n_430),
.B1(n_423),
.B2(n_422),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_451),
.B1(n_444),
.B2(n_416),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_475),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_480),
.C(n_483),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_461),
.A2(n_442),
.B1(n_447),
.B2(n_435),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_383),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_459),
.B1(n_465),
.B2(n_466),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_436),
.C(n_443),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_449),
.B1(n_452),
.B2(n_456),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_445),
.C(n_455),
.Y(n_483)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_484),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_432),
.C(n_446),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_279),
.C(n_290),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_460),
.A2(n_468),
.B(n_463),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_293),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_485),
.A2(n_470),
.B(n_451),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_490),
.A2(n_495),
.B(n_487),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_446),
.B(n_458),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_496),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_481),
.Y(n_493)
);

INVx6_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_494),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_357),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_469),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_342),
.C(n_337),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_499),
.C(n_501),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_291),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_479),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_495),
.A2(n_476),
.B1(n_484),
.B2(n_486),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_504),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_493),
.A2(n_476),
.B1(n_486),
.B2(n_478),
.Y(n_504)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_505),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_507),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_483),
.Y(n_507)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_510),
.Y(n_511)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_511),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_489),
.C(n_492),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_515),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_501),
.Y(n_515)
);

OAI321xp33_ASAP7_75t_L g519 ( 
.A1(n_513),
.A2(n_502),
.A3(n_505),
.B1(n_498),
.B2(n_508),
.C(n_474),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_519),
.A2(n_514),
.B(n_511),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_516),
.A2(n_509),
.B(n_492),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_512),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_522),
.B(n_518),
.C(n_517),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_523),
.A2(n_496),
.B(n_297),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_246),
.Y(n_525)
);

OAI21xp33_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_245),
.B(n_242),
.Y(n_526)
);

MAJx2_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_242),
.C(n_245),
.Y(n_527)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_527),
.Y(n_528)
);


endmodule