module real_aes_17609_n_376 (n_76, n_113, n_1999, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_1999;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1994;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_1632;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1973;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1985;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1691;
wire n_640;
wire n_1931;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1889;
wire n_1533;
wire n_1679;
wire n_460;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_0), .A2(n_119), .B1(n_644), .B2(n_684), .C(n_687), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_0), .A2(n_248), .B1(n_724), .B2(n_726), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1720 ( .A1(n_1), .A2(n_96), .B1(n_1677), .B2(n_1680), .Y(n_1720) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_2), .A2(n_297), .B1(n_872), .B2(n_1460), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1478 ( .A1(n_2), .A2(n_260), .B1(n_557), .B2(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g786 ( .A(n_3), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_4), .A2(n_127), .B1(n_534), .B2(n_613), .Y(n_1318) );
OAI22xp33_ASAP7_75t_L g1352 ( .A1(n_4), .A2(n_202), .B1(n_464), .B2(n_467), .Y(n_1352) );
AND2x2_ASAP7_75t_L g484 ( .A(n_5), .B(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_5), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g529 ( .A(n_5), .Y(n_529) );
AND2x2_ASAP7_75t_L g537 ( .A(n_5), .B(n_267), .Y(n_537) );
INVx1_ASAP7_75t_L g587 ( .A(n_6), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_6), .A2(n_14), .B1(n_616), .B2(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g1091 ( .A(n_7), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_7), .A2(n_87), .B1(n_401), .B2(n_1102), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1972 ( .A1(n_8), .A2(n_287), .B1(n_1973), .B2(n_1974), .Y(n_1972) );
OAI22xp33_ASAP7_75t_L g1985 ( .A1(n_8), .A2(n_287), .B1(n_1986), .B2(n_1988), .Y(n_1985) );
OAI22xp33_ASAP7_75t_L g1890 ( .A1(n_9), .A2(n_307), .B1(n_1891), .B2(n_1892), .Y(n_1890) );
OAI22xp33_ASAP7_75t_L g1903 ( .A1(n_9), .A2(n_307), .B1(n_1904), .B2(n_1905), .Y(n_1903) );
INVx1_ASAP7_75t_L g462 ( .A(n_10), .Y(n_462) );
INVx1_ASAP7_75t_L g916 ( .A(n_11), .Y(n_916) );
INVx1_ASAP7_75t_L g661 ( .A(n_12), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_12), .A2(n_102), .B1(n_738), .B2(n_742), .Y(n_737) );
INVx1_ASAP7_75t_L g1078 ( .A(n_13), .Y(n_1078) );
INVx1_ASAP7_75t_L g603 ( .A(n_14), .Y(n_603) );
INVxp67_ASAP7_75t_SL g903 ( .A(n_15), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_15), .A2(n_134), .B1(n_424), .B2(n_814), .Y(n_937) );
INVx1_ASAP7_75t_L g898 ( .A(n_16), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_16), .A2(n_182), .B1(n_727), .B2(n_808), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g1462 ( .A1(n_17), .A2(n_221), .B1(n_720), .B2(n_1463), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_17), .A2(n_131), .B1(n_650), .B2(n_758), .C(n_1477), .Y(n_1476) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_18), .A2(n_365), .B1(n_401), .B2(n_406), .C(n_412), .Y(n_1128) );
OAI21xp33_ASAP7_75t_SL g1155 ( .A1(n_18), .A2(n_545), .B(n_1068), .Y(n_1155) );
INVx1_ASAP7_75t_L g1969 ( .A(n_19), .Y(n_1969) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_20), .A2(n_101), .B1(n_644), .B2(n_646), .C(n_649), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_20), .A2(n_214), .B1(n_424), .B2(n_721), .Y(n_736) );
INVx2_ASAP7_75t_L g397 ( .A(n_21), .Y(n_397) );
INVx1_ASAP7_75t_L g785 ( .A(n_22), .Y(n_785) );
OAI322xp33_ASAP7_75t_L g789 ( .A1(n_22), .A2(n_790), .A3(n_796), .B1(n_798), .B2(n_805), .C1(n_815), .C2(n_818), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_23), .A2(n_182), .B1(n_557), .B2(n_653), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_23), .A2(n_333), .B1(n_727), .B2(n_940), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g1253 ( .A(n_24), .Y(n_1253) );
INVx1_ASAP7_75t_L g1944 ( .A(n_25), .Y(n_1944) );
AOI221xp5_ASAP7_75t_L g775 ( .A1(n_26), .A2(n_247), .B1(n_649), .B2(n_776), .C(n_777), .Y(n_775) );
INVx1_ASAP7_75t_L g803 ( .A(n_26), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g1139 ( .A1(n_27), .A2(n_311), .B1(n_464), .B2(n_467), .Y(n_1139) );
INVx1_ASAP7_75t_L g1154 ( .A(n_27), .Y(n_1154) );
OAI211xp5_ASAP7_75t_L g1967 ( .A1(n_28), .A2(n_520), .B(n_1562), .C(n_1968), .Y(n_1967) );
INVx1_ASAP7_75t_L g1984 ( .A(n_28), .Y(n_1984) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_29), .A2(n_364), .B1(n_432), .B2(n_731), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_29), .A2(n_179), .B1(n_630), .B2(n_632), .Y(n_1439) );
INVx1_ASAP7_75t_L g1924 ( .A(n_30), .Y(n_1924) );
XOR2x1_ASAP7_75t_L g1362 ( .A(n_31), .B(n_1363), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_32), .A2(n_340), .B1(n_464), .B2(n_467), .Y(n_463) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_32), .Y(n_475) );
INVx1_ASAP7_75t_L g1202 ( .A(n_33), .Y(n_1202) );
AOI221xp5_ASAP7_75t_L g1217 ( .A1(n_33), .A2(n_160), .B1(n_1017), .B2(n_1218), .C(n_1220), .Y(n_1217) );
INVx1_ASAP7_75t_L g1049 ( .A(n_34), .Y(n_1049) );
AOI221x1_ASAP7_75t_SL g1054 ( .A1(n_34), .A2(n_213), .B1(n_557), .B2(n_848), .C(n_1055), .Y(n_1054) );
OA22x2_ASAP7_75t_L g1489 ( .A1(n_35), .A2(n_1490), .B1(n_1590), .B2(n_1591), .Y(n_1489) );
INVxp67_ASAP7_75t_L g1591 ( .A(n_35), .Y(n_1591) );
HB1xp67_ASAP7_75t_L g1656 ( .A(n_36), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_36), .B(n_1654), .Y(n_1671) );
INVx1_ASAP7_75t_L g1952 ( .A(n_37), .Y(n_1952) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_38), .A2(n_319), .B1(n_764), .B2(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_L g794 ( .A(n_38), .Y(n_794) );
INVx1_ASAP7_75t_L g1042 ( .A(n_39), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_39), .A2(n_196), .B1(n_618), .B2(n_764), .Y(n_1062) );
INVx1_ASAP7_75t_L g1531 ( .A(n_40), .Y(n_1531) );
INVx1_ASAP7_75t_L g750 ( .A(n_41), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_42), .A2(n_278), .B1(n_455), .B2(n_574), .Y(n_1369) );
INVxp33_ASAP7_75t_L g1412 ( .A(n_42), .Y(n_1412) );
INVx1_ASAP7_75t_L g443 ( .A(n_43), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_44), .A2(n_318), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_44), .A2(n_247), .B1(n_424), .B2(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g1209 ( .A(n_45), .Y(n_1209) );
OAI22xp33_ASAP7_75t_L g1215 ( .A1(n_45), .A2(n_56), .B1(n_401), .B2(n_406), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1719 ( .A1(n_46), .A2(n_74), .B1(n_1670), .B2(n_1674), .Y(n_1719) );
AOI22xp33_ASAP7_75t_L g1459 ( .A1(n_47), .A2(n_260), .B1(n_872), .B2(n_1460), .Y(n_1459) );
AOI221xp5_ASAP7_75t_L g1473 ( .A1(n_47), .A2(n_297), .B1(n_645), .B2(n_648), .C(n_975), .Y(n_1473) );
OAI22xp33_ASAP7_75t_L g1880 ( .A1(n_48), .A2(n_189), .B1(n_1881), .B2(n_1883), .Y(n_1880) );
OAI22xp33_ASAP7_75t_L g1907 ( .A1(n_48), .A2(n_189), .B1(n_1582), .B2(n_1908), .Y(n_1907) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_49), .A2(n_949), .B1(n_950), .B2(n_951), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_49), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_50), .Y(n_1040) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_51), .Y(n_905) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_51), .A2(n_98), .B1(n_424), .B2(n_814), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_52), .A2(n_574), .B1(n_1239), .B2(n_1242), .Y(n_1238) );
INVx1_ASAP7_75t_L g1259 ( .A(n_52), .Y(n_1259) );
CKINVDCx5p33_ASAP7_75t_R g1454 ( .A(n_53), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_54), .A2(n_208), .B1(n_557), .B2(n_621), .Y(n_976) );
INVx1_ASAP7_75t_L g1006 ( .A(n_54), .Y(n_1006) );
AOI221xp5_ASAP7_75t_L g1325 ( .A1(n_55), .A2(n_71), .B1(n_1266), .B2(n_1326), .C(n_1328), .Y(n_1325) );
AOI221xp5_ASAP7_75t_L g1349 ( .A1(n_55), .A2(n_151), .B1(n_424), .B2(n_1344), .C(n_1350), .Y(n_1349) );
OAI221xp5_ASAP7_75t_L g1205 ( .A1(n_56), .A2(n_327), .B1(n_532), .B2(n_541), .C(n_545), .Y(n_1205) );
INVx1_ASAP7_75t_L g386 ( .A(n_57), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g1430 ( .A1(n_58), .A2(n_143), .B1(n_721), .B2(n_859), .Y(n_1430) );
INVxp67_ASAP7_75t_SL g1445 ( .A(n_58), .Y(n_1445) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_59), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_60), .A2(n_424), .B(n_426), .Y(n_423) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_60), .Y(n_505) );
INVx1_ASAP7_75t_L g1467 ( .A(n_61), .Y(n_1467) );
INVx1_ASAP7_75t_L g585 ( .A(n_62), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_62), .A2(n_203), .B1(n_616), .B2(n_625), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_63), .A2(n_124), .B1(n_1670), .B2(n_1674), .Y(n_1695) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_64), .Y(n_1197) );
AOI22xp5_ASAP7_75t_L g1685 ( .A1(n_65), .A2(n_274), .B1(n_1670), .B2(n_1674), .Y(n_1685) );
INVx1_ASAP7_75t_L g1246 ( .A(n_66), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_66), .A2(n_68), .B1(n_621), .B2(n_641), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_67), .A2(n_230), .B1(n_653), .B2(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g1000 ( .A(n_67), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_68), .A2(n_358), .B1(n_451), .B2(n_727), .C(n_1234), .Y(n_1233) );
OAI222xp33_ASAP7_75t_L g829 ( .A1(n_69), .A2(n_88), .B1(n_666), .B2(n_830), .C1(n_838), .C2(n_844), .Y(n_829) );
INVx1_ASAP7_75t_L g864 ( .A(n_69), .Y(n_864) );
INVxp67_ASAP7_75t_SL g1207 ( .A(n_70), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_70), .A2(n_574), .B1(n_1222), .B2(n_1223), .Y(n_1221) );
INVx1_ASAP7_75t_L g1346 ( .A(n_71), .Y(n_1346) );
AOI22xp33_ASAP7_75t_SL g1291 ( .A1(n_72), .A2(n_188), .B1(n_726), .B2(n_1282), .Y(n_1291) );
AOI221xp5_ASAP7_75t_L g1305 ( .A1(n_72), .A2(n_141), .B1(n_617), .B2(n_1306), .C(n_1309), .Y(n_1305) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_73), .A2(n_270), .B1(n_401), .B2(n_406), .C(n_412), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_73), .A2(n_340), .B1(n_532), .B2(n_541), .C(n_545), .Y(n_531) );
INVx1_ASAP7_75t_L g1295 ( .A(n_75), .Y(n_1295) );
AOI21xp33_ASAP7_75t_L g1140 ( .A1(n_76), .A2(n_1141), .B(n_1144), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_76), .A2(n_120), .B1(n_644), .B2(n_1169), .C(n_1170), .Y(n_1168) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_77), .Y(n_821) );
INVx1_ASAP7_75t_L g771 ( .A(n_78), .Y(n_771) );
OAI211xp5_ASAP7_75t_L g822 ( .A1(n_78), .A2(n_738), .B(n_746), .C(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g1707 ( .A1(n_79), .A2(n_253), .B1(n_1670), .B2(n_1674), .Y(n_1707) );
INVx1_ASAP7_75t_L g1211 ( .A(n_80), .Y(n_1211) );
OAI222xp33_ASAP7_75t_L g1214 ( .A1(n_80), .A2(n_316), .B1(n_327), .B2(n_459), .C1(n_804), .C2(n_1037), .Y(n_1214) );
INVxp67_ASAP7_75t_SL g1337 ( .A(n_81), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_81), .A2(n_121), .B1(n_455), .B2(n_574), .Y(n_1341) );
INVx1_ASAP7_75t_L g1925 ( .A(n_82), .Y(n_1925) );
INVx1_ASAP7_75t_L g1296 ( .A(n_83), .Y(n_1296) );
INVx1_ASAP7_75t_L g1422 ( .A(n_84), .Y(n_1422) );
XOR2x2_ASAP7_75t_L g1123 ( .A(n_85), .B(n_1124), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g1689 ( .A1(n_85), .A2(n_265), .B1(n_1677), .B2(n_1680), .Y(n_1689) );
AOI22xp33_ASAP7_75t_L g1616 ( .A1(n_86), .A2(n_338), .B1(n_1289), .B2(n_1617), .Y(n_1616) );
AOI221xp5_ASAP7_75t_L g1628 ( .A1(n_86), .A2(n_355), .B1(n_616), .B2(n_650), .C(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1083 ( .A(n_87), .Y(n_1083) );
INVx1_ASAP7_75t_L g865 ( .A(n_88), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g1520 ( .A1(n_89), .A2(n_204), .B1(n_1521), .B2(n_1523), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1573 ( .A1(n_89), .A2(n_204), .B1(n_1574), .B2(n_1578), .Y(n_1573) );
AOI22xp5_ASAP7_75t_L g1690 ( .A1(n_90), .A2(n_111), .B1(n_1670), .B2(n_1691), .Y(n_1690) );
XNOR2xp5_ASAP7_75t_L g1414 ( .A(n_91), .B(n_1415), .Y(n_1414) );
AO22x1_ASAP7_75t_L g1713 ( .A1(n_91), .A2(n_275), .B1(n_1677), .B2(n_1680), .Y(n_1713) );
NAND2xp33_ASAP7_75t_SL g1324 ( .A(n_92), .B(n_900), .Y(n_1324) );
INVx1_ASAP7_75t_L g1351 ( .A(n_92), .Y(n_1351) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_93), .A2(n_142), .B1(n_955), .B2(n_956), .C(n_959), .Y(n_954) );
INVx1_ASAP7_75t_L g984 ( .A(n_93), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_94), .Y(n_928) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_95), .A2(n_215), .B1(n_464), .B2(n_467), .Y(n_1382) );
INVxp67_ASAP7_75t_SL g1396 ( .A(n_95), .Y(n_1396) );
XOR2xp5_ASAP7_75t_L g1450 ( .A(n_96), .B(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1548 ( .A(n_97), .Y(n_1548) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_98), .A2(n_134), .B1(n_616), .B2(n_850), .C(n_911), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_99), .A2(n_216), .B1(n_699), .B2(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g961 ( .A(n_100), .Y(n_961) );
OAI221xp5_ASAP7_75t_SL g989 ( .A1(n_100), .A2(n_137), .B1(n_404), .B2(n_712), .C(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_101), .A2(n_295), .B1(n_717), .B2(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g658 ( .A(n_102), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_103), .A2(n_224), .B1(n_455), .B2(n_574), .Y(n_1129) );
INVxp67_ASAP7_75t_SL g1167 ( .A(n_103), .Y(n_1167) );
INVx1_ASAP7_75t_L g1274 ( .A(n_104), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_105), .B(n_874), .Y(n_1381) );
AOI221xp5_ASAP7_75t_L g1410 ( .A1(n_105), .A2(n_233), .B1(n_630), .B2(n_632), .C(n_1266), .Y(n_1410) );
INVx1_ASAP7_75t_L g1482 ( .A(n_106), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_107), .A2(n_335), .B1(n_720), .B2(n_874), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_107), .A2(n_156), .B1(n_1301), .B2(n_1304), .Y(n_1303) );
AOI222xp33_ASAP7_75t_L g1145 ( .A1(n_108), .A2(n_169), .B1(n_353), .B2(n_432), .C1(n_452), .C2(n_593), .Y(n_1145) );
INVx1_ASAP7_75t_L g1172 ( .A(n_108), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_109), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_110), .B(n_1377), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_110), .A2(n_192), .B1(n_625), .B2(n_644), .Y(n_1409) );
INVx1_ASAP7_75t_L g1279 ( .A(n_112), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_113), .A2(n_211), .B1(n_1289), .B2(n_1426), .Y(n_1425) );
INVxp67_ASAP7_75t_SL g1444 ( .A(n_113), .Y(n_1444) );
OAI22xp33_ASAP7_75t_L g1254 ( .A1(n_114), .A2(n_164), .B1(n_401), .B2(n_406), .Y(n_1254) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_114), .A2(n_315), .B1(n_532), .B2(n_541), .Y(n_1269) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_115), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_115), .A2(n_302), .B1(n_424), .B2(n_721), .Y(n_870) );
INVx1_ASAP7_75t_L g1549 ( .A(n_116), .Y(n_1549) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_117), .Y(n_1203) );
OAI221xp5_ASAP7_75t_L g1599 ( .A1(n_118), .A2(n_243), .B1(n_881), .B2(n_1600), .C(n_1601), .Y(n_1599) );
OAI211xp5_ASAP7_75t_L g1624 ( .A1(n_118), .A2(n_1442), .B(n_1625), .C(n_1630), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_119), .A2(n_298), .B1(n_729), .B2(n_731), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_120), .A2(n_236), .B1(n_1132), .B2(n_1134), .C(n_1136), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g1354 ( .A(n_121), .Y(n_1354) );
INVx1_ASAP7_75t_L g1654 ( .A(n_122), .Y(n_1654) );
INVx1_ASAP7_75t_L g1241 ( .A(n_123), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_123), .A2(n_358), .B1(n_557), .B2(n_621), .Y(n_1265) );
XOR2x2_ASAP7_75t_L g1877 ( .A(n_124), .B(n_1878), .Y(n_1877) );
AOI22xp5_ASAP7_75t_L g1935 ( .A1(n_124), .A2(n_1936), .B1(n_1991), .B2(n_1994), .Y(n_1935) );
INVx1_ASAP7_75t_L g1208 ( .A(n_125), .Y(n_1208) );
AO221x2_ASAP7_75t_L g1780 ( .A1(n_126), .A2(n_354), .B1(n_1677), .B2(n_1680), .C(n_1781), .Y(n_1780) );
OAI221xp5_ASAP7_75t_L g1340 ( .A1(n_127), .A2(n_149), .B1(n_401), .B2(n_406), .C(n_412), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_128), .A2(n_171), .B1(n_776), .B2(n_848), .C(n_850), .Y(n_977) );
INVx1_ASAP7_75t_L g995 ( .A(n_128), .Y(n_995) );
INVx1_ASAP7_75t_L g1127 ( .A(n_129), .Y(n_1127) );
OAI21xp33_ASAP7_75t_L g1151 ( .A1(n_129), .A2(n_1067), .B(n_1152), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1622 ( .A1(n_130), .A2(n_283), .B1(n_699), .B2(n_701), .Y(n_1622) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_131), .A2(n_266), .B1(n_1284), .B2(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1947 ( .A(n_132), .Y(n_1947) );
INVx1_ASAP7_75t_L g601 ( .A(n_133), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_133), .A2(n_181), .B1(n_557), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g1281 ( .A1(n_135), .A2(n_141), .B1(n_1282), .B2(n_1284), .Y(n_1281) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_135), .A2(n_326), .B1(n_644), .B2(n_650), .C(n_758), .Y(n_1298) );
INVx1_ASAP7_75t_L g1331 ( .A(n_136), .Y(n_1331) );
INVx1_ASAP7_75t_L g970 ( .A(n_137), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_138), .Y(n_581) );
INVx1_ASAP7_75t_L g854 ( .A(n_139), .Y(n_854) );
INVx1_ASAP7_75t_L g1021 ( .A(n_140), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_140), .A2(n_263), .B1(n_532), .B2(n_541), .Y(n_1063) );
INVx1_ASAP7_75t_L g982 ( .A(n_142), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g1435 ( .A1(n_143), .A2(n_211), .B1(n_650), .B2(n_1306), .C(n_1436), .Y(n_1435) );
OAI21xp5_ASAP7_75t_SL g1312 ( .A1(n_144), .A2(n_699), .B(n_1313), .Y(n_1312) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_145), .A2(n_308), .B1(n_455), .B2(n_574), .C(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g633 ( .A(n_145), .Y(n_633) );
INVx1_ASAP7_75t_L g1921 ( .A(n_146), .Y(n_1921) );
INVx1_ASAP7_75t_L g967 ( .A(n_147), .Y(n_967) );
OAI21xp33_ASAP7_75t_L g987 ( .A1(n_147), .A2(n_694), .B(n_988), .Y(n_987) );
CKINVDCx5p33_ASAP7_75t_R g1236 ( .A(n_148), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1336 ( .A(n_149), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_150), .A2(n_334), .B1(n_401), .B2(n_406), .C(n_412), .Y(n_1368) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_150), .B(n_561), .Y(n_1400) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_151), .A2(n_157), .B1(n_623), .B2(n_1328), .C(n_1333), .Y(n_1332) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_152), .A2(n_276), .B1(n_653), .B2(n_1088), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_152), .A2(n_352), .B1(n_424), .B2(n_426), .C(n_1108), .Y(n_1109) );
OAI22xp33_ASAP7_75t_L g1975 ( .A1(n_153), .A2(n_339), .B1(n_1976), .B2(n_1977), .Y(n_1975) );
OAI22xp5_ASAP7_75t_L g1979 ( .A1(n_153), .A2(n_339), .B1(n_1501), .B2(n_1980), .Y(n_1979) );
INVx1_ASAP7_75t_L g768 ( .A(n_154), .Y(n_768) );
OAI211xp5_ASAP7_75t_SL g908 ( .A1(n_155), .A2(n_639), .B(n_909), .C(n_914), .Y(n_908) );
INVx1_ASAP7_75t_L g935 ( .A(n_155), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_156), .A2(n_326), .B1(n_1284), .B2(n_1289), .C(n_1290), .Y(n_1288) );
INVx1_ASAP7_75t_L g1348 ( .A(n_157), .Y(n_1348) );
AO22x1_ASAP7_75t_L g1676 ( .A1(n_158), .A2(n_359), .B1(n_1677), .B2(n_1680), .Y(n_1676) );
OAI222xp33_ASAP7_75t_L g893 ( .A1(n_159), .A2(n_289), .B1(n_671), .B2(n_894), .C1(n_895), .C2(n_902), .Y(n_893) );
INVx1_ASAP7_75t_L g931 ( .A(n_159), .Y(n_931) );
INVx1_ASAP7_75t_L g1185 ( .A(n_160), .Y(n_1185) );
INVx1_ASAP7_75t_L g1608 ( .A(n_161), .Y(n_1608) );
INVx1_ASAP7_75t_L g836 ( .A(n_162), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_162), .A2(n_220), .B1(n_872), .B2(n_874), .Y(n_871) );
XNOR2x1_ASAP7_75t_L g889 ( .A(n_163), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g1260 ( .A(n_164), .Y(n_1260) );
AOI221xp5_ASAP7_75t_SL g974 ( .A1(n_165), .A2(n_332), .B1(n_776), .B2(n_848), .C(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g1003 ( .A(n_165), .Y(n_1003) );
INVx1_ASAP7_75t_L g1889 ( .A(n_166), .Y(n_1889) );
OAI211xp5_ASAP7_75t_L g1895 ( .A1(n_166), .A2(n_1896), .B(n_1897), .C(n_1898), .Y(n_1895) );
OAI222xp33_ASAP7_75t_L g1431 ( .A1(n_167), .A2(n_261), .B1(n_272), .B2(n_693), .C1(n_699), .C2(n_701), .Y(n_1431) );
OAI211xp5_ASAP7_75t_L g1433 ( .A1(n_167), .A2(n_639), .B(n_1434), .C(n_1440), .Y(n_1433) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_168), .Y(n_972) );
INVx1_ASAP7_75t_L g1163 ( .A(n_169), .Y(n_1163) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_170), .A2(n_223), .B1(n_758), .B2(n_759), .C(n_762), .Y(n_757) );
INVxp67_ASAP7_75t_L g791 ( .A(n_170), .Y(n_791) );
INVx1_ASAP7_75t_L g1007 ( .A(n_171), .Y(n_1007) );
XOR2xp5_ASAP7_75t_L g1937 ( .A(n_172), .B(n_1938), .Y(n_1937) );
INVx1_ASAP7_75t_L g1919 ( .A(n_173), .Y(n_1919) );
INVxp67_ASAP7_75t_SL g1604 ( .A(n_174), .Y(n_1604) );
AOI221xp5_ASAP7_75t_L g1638 ( .A1(n_174), .A2(n_273), .B1(n_645), .B2(n_975), .C(n_1629), .Y(n_1638) );
INVx1_ASAP7_75t_L g577 ( .A(n_175), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_175), .A2(n_349), .B1(n_534), .B2(n_613), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_176), .Y(n_1033) );
AO22x1_ASAP7_75t_L g1711 ( .A1(n_177), .A2(n_360), .B1(n_1670), .B2(n_1712), .Y(n_1711) );
CKINVDCx16_ASAP7_75t_R g1782 ( .A(n_178), .Y(n_1782) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_179), .A2(n_363), .B1(n_729), .B2(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g1922 ( .A(n_180), .Y(n_1922) );
INVx1_ASAP7_75t_L g591 ( .A(n_181), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_183), .A2(n_367), .B1(n_451), .B2(n_452), .Y(n_450) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_183), .Y(n_525) );
INVx1_ASAP7_75t_L g1453 ( .A(n_184), .Y(n_1453) );
INVx1_ASAP7_75t_L g1248 ( .A(n_185), .Y(n_1248) );
INVx1_ASAP7_75t_L g1621 ( .A(n_186), .Y(n_1621) );
INVx1_ASAP7_75t_L g419 ( .A(n_187), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g1299 ( .A1(n_188), .A2(n_335), .B1(n_1300), .B2(n_1301), .Y(n_1299) );
INVx1_ASAP7_75t_L g1419 ( .A(n_190), .Y(n_1419) );
OAI221xp5_ASAP7_75t_SL g1441 ( .A1(n_190), .A2(n_197), .B1(n_671), .B2(n_1442), .C(n_1443), .Y(n_1441) );
INVx1_ASAP7_75t_L g1970 ( .A(n_191), .Y(n_1970) );
OAI211xp5_ASAP7_75t_L g1981 ( .A1(n_191), .A2(n_1508), .B(n_1609), .C(n_1982), .Y(n_1981) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_192), .A2(n_219), .B1(n_1384), .B2(n_1387), .C(n_1388), .Y(n_1383) );
INVx1_ASAP7_75t_L g915 ( .A(n_193), .Y(n_915) );
INVx1_ASAP7_75t_L g1915 ( .A(n_194), .Y(n_1915) );
INVx1_ASAP7_75t_L g1367 ( .A(n_195), .Y(n_1367) );
INVx1_ASAP7_75t_L g1035 ( .A(n_196), .Y(n_1035) );
INVx1_ASAP7_75t_L g1420 ( .A(n_197), .Y(n_1420) );
INVx2_ASAP7_75t_L g1673 ( .A(n_198), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_198), .B(n_321), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_198), .B(n_1679), .Y(n_1681) );
AOI21xp5_ASAP7_75t_L g1379 ( .A1(n_199), .A2(n_424), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1407 ( .A(n_199), .Y(n_1407) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_200), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_200), .A2(n_336), .B1(n_879), .B2(n_880), .Y(n_878) );
INVx1_ASAP7_75t_L g1469 ( .A(n_201), .Y(n_1469) );
OAI211xp5_ASAP7_75t_L g1316 ( .A1(n_202), .A2(n_477), .B(n_1317), .C(n_1334), .Y(n_1316) );
INVx1_ASAP7_75t_L g599 ( .A(n_203), .Y(n_599) );
INVx1_ASAP7_75t_L g634 ( .A(n_205), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g1080 ( .A1(n_206), .A2(n_1065), .B(n_1081), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1112 ( .A1(n_206), .A2(n_305), .B1(n_1113), .B2(n_1114), .C(n_1115), .Y(n_1112) );
INVx1_ASAP7_75t_L g1888 ( .A(n_207), .Y(n_1888) );
INVx1_ASAP7_75t_L g994 ( .A(n_208), .Y(n_994) );
INVx1_ASAP7_75t_L g441 ( .A(n_209), .Y(n_441) );
INVx1_ASAP7_75t_L g1945 ( .A(n_210), .Y(n_1945) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_212), .Y(n_1030) );
INVx1_ASAP7_75t_L g1038 ( .A(n_213), .Y(n_1038) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_214), .Y(n_682) );
INVx1_ASAP7_75t_L g1364 ( .A(n_215), .Y(n_1364) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_216), .A2(n_639), .B(n_642), .C(n_657), .Y(n_638) );
INVx1_ASAP7_75t_L g1356 ( .A(n_217), .Y(n_1356) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_218), .A2(n_341), .B1(n_625), .B2(n_779), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_218), .A2(n_244), .B1(n_448), .B2(n_872), .C(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1408 ( .A(n_219), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_220), .A2(n_371), .B1(n_764), .B2(n_765), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_221), .A2(n_266), .B1(n_653), .B2(n_1088), .Y(n_1474) );
INVx2_ASAP7_75t_L g399 ( .A(n_222), .Y(n_399) );
INVx1_ASAP7_75t_L g429 ( .A(n_222), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_222), .B(n_397), .Y(n_458) );
INVxp67_ASAP7_75t_L g809 ( .A(n_223), .Y(n_809) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_224), .Y(n_1147) );
XOR2xp5_ASAP7_75t_L g1009 ( .A(n_225), .B(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1179 ( .A(n_226), .Y(n_1179) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_227), .A2(n_322), .B1(n_666), .B2(n_670), .C(n_675), .Y(n_665) );
INVx1_ASAP7_75t_L g706 ( .A(n_227), .Y(n_706) );
INVx1_ASAP7_75t_L g604 ( .A(n_228), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_228), .A2(n_343), .B1(n_630), .B2(n_632), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_229), .A2(n_331), .B1(n_600), .B2(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1071 ( .A(n_229), .Y(n_1071) );
INVx1_ASAP7_75t_L g1004 ( .A(n_230), .Y(n_1004) );
INVx1_ASAP7_75t_L g1540 ( .A(n_231), .Y(n_1540) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_232), .A2(n_351), .B1(n_653), .B2(n_654), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_232), .A2(n_276), .B1(n_424), .B2(n_727), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_233), .A2(n_290), .B1(n_727), .B2(n_808), .Y(n_1389) );
INVx1_ASAP7_75t_L g833 ( .A(n_234), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_234), .A2(n_371), .B1(n_874), .B2(n_876), .Y(n_875) );
BUFx3_ASAP7_75t_L g391 ( .A(n_235), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_236), .B(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1137 ( .A(n_237), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1708 ( .A1(n_238), .A2(n_246), .B1(n_1677), .B2(n_1680), .Y(n_1708) );
INVx1_ASAP7_75t_L g1082 ( .A(n_239), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_240), .A2(n_315), .B1(n_1250), .B2(n_1251), .C(n_1252), .Y(n_1249) );
OAI211xp5_ASAP7_75t_L g1257 ( .A1(n_240), .A2(n_1119), .B(n_1258), .C(n_1261), .Y(n_1257) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_241), .A2(n_699), .B(n_857), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_242), .Y(n_1235) );
OAI221xp5_ASAP7_75t_SL g1631 ( .A1(n_243), .A2(n_348), .B1(n_844), .B2(n_1632), .C(n_1634), .Y(n_1631) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_244), .A2(n_352), .B1(n_684), .B2(n_1097), .Y(n_1096) );
OAI21xp5_ASAP7_75t_L g920 ( .A1(n_245), .A2(n_921), .B(n_922), .Y(n_920) );
XOR2xp5_ASAP7_75t_L g635 ( .A(n_246), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_248), .A2(n_298), .B1(n_652), .B2(n_654), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g1505 ( .A1(n_249), .A2(n_1506), .B(n_1508), .C(n_1510), .Y(n_1505) );
INVx1_ASAP7_75t_L g1569 ( .A(n_249), .Y(n_1569) );
INVx1_ASAP7_75t_L g1914 ( .A(n_250), .Y(n_1914) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_251), .Y(n_697) );
INVx1_ASAP7_75t_L g460 ( .A(n_252), .Y(n_460) );
INVx1_ASAP7_75t_L g1918 ( .A(n_254), .Y(n_1918) );
INVx1_ASAP7_75t_L g1519 ( .A(n_255), .Y(n_1519) );
OAI211xp5_ASAP7_75t_SL g1560 ( .A1(n_255), .A2(n_1561), .B(n_1562), .C(n_1565), .Y(n_1560) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_256), .Y(n_1193) );
INVx1_ASAP7_75t_L g1335 ( .A(n_257), .Y(n_1335) );
INVx1_ASAP7_75t_L g853 ( .A(n_258), .Y(n_853) );
INVx1_ASAP7_75t_L g1373 ( .A(n_259), .Y(n_1373) );
OAI211xp5_ASAP7_75t_L g578 ( .A1(n_262), .A2(n_388), .B(n_412), .C(n_579), .Y(n_578) );
INVxp33_ASAP7_75t_SL g611 ( .A(n_262), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g1026 ( .A1(n_263), .A2(n_286), .B1(n_404), .B2(n_584), .C(n_712), .Y(n_1026) );
INVx1_ASAP7_75t_L g1278 ( .A(n_264), .Y(n_1278) );
INVx1_ASAP7_75t_L g485 ( .A(n_267), .Y(n_485) );
BUFx3_ASAP7_75t_L g498 ( .A(n_267), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g1784 ( .A(n_268), .Y(n_1784) );
AOI22xp5_ASAP7_75t_L g1684 ( .A1(n_269), .A2(n_291), .B1(n_1677), .B2(n_1680), .Y(n_1684) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_270), .Y(n_562) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_271), .A2(n_639), .B(n_846), .C(n_852), .Y(n_845) );
INVx1_ASAP7_75t_L g867 ( .A(n_271), .Y(n_867) );
INVx1_ASAP7_75t_L g1612 ( .A(n_273), .Y(n_1612) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_277), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g1391 ( .A(n_278), .Y(n_1391) );
OAI322xp33_ASAP7_75t_SL g1602 ( .A1(n_279), .A2(n_1551), .A3(n_1603), .B1(n_1607), .B2(n_1611), .C1(n_1618), .C2(n_1619), .Y(n_1602) );
OAI22xp33_ASAP7_75t_SL g1639 ( .A1(n_279), .A2(n_283), .B1(n_639), .B2(n_1640), .Y(n_1639) );
INVxp67_ASAP7_75t_SL g1074 ( .A(n_280), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_281), .Y(n_960) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_282), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_284), .Y(n_1244) );
INVx1_ASAP7_75t_L g1615 ( .A(n_285), .Y(n_1615) );
OA222x2_ASAP7_75t_L g1064 ( .A1(n_286), .A2(n_303), .B1(n_356), .B2(n_1065), .C1(n_1067), .C2(n_1068), .Y(n_1064) );
INVx1_ASAP7_75t_L g1954 ( .A(n_288), .Y(n_1954) );
INVx1_ASAP7_75t_L g932 ( .A(n_289), .Y(n_932) );
AOI32xp33_ASAP7_75t_L g1398 ( .A1(n_290), .A2(n_758), .A3(n_1399), .B1(n_1401), .B2(n_1999), .Y(n_1398) );
OAI21xp5_ASAP7_75t_L g1485 ( .A1(n_292), .A2(n_699), .B(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1138 ( .A(n_293), .Y(n_1138) );
XOR2x2_ASAP7_75t_L g826 ( .A(n_294), .B(n_827), .Y(n_826) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_295), .Y(n_679) );
OAI22xp5_ASAP7_75t_SL g1593 ( .A1(n_296), .A2(n_1594), .B1(n_1595), .B2(n_1641), .Y(n_1593) );
INVx1_ASAP7_75t_L g1641 ( .A(n_296), .Y(n_1641) );
AOI22xp5_ASAP7_75t_L g1643 ( .A1(n_296), .A2(n_1594), .B1(n_1595), .B2(n_1641), .Y(n_1643) );
AOI22xp5_ASAP7_75t_L g1694 ( .A1(n_299), .A2(n_362), .B1(n_1677), .B2(n_1680), .Y(n_1694) );
AO22x1_ASAP7_75t_L g1669 ( .A1(n_300), .A2(n_309), .B1(n_1670), .B2(n_1674), .Y(n_1669) );
INVx1_ASAP7_75t_L g394 ( .A(n_301), .Y(n_394) );
INVx1_ASAP7_75t_L g411 ( .A(n_301), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g847 ( .A1(n_302), .A2(n_336), .B1(n_758), .B2(n_848), .C(n_850), .Y(n_847) );
INVx1_ASAP7_75t_L g1025 ( .A(n_303), .Y(n_1025) );
INVx1_ASAP7_75t_L g1093 ( .A(n_304), .Y(n_1093) );
INVxp67_ASAP7_75t_SL g1120 ( .A(n_305), .Y(n_1120) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_306), .Y(n_1189) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_308), .Y(n_609) );
INVx1_ASAP7_75t_L g1542 ( .A(n_310), .Y(n_1542) );
INVxp67_ASAP7_75t_SL g1150 ( .A(n_311), .Y(n_1150) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_312), .A2(n_447), .B(n_448), .Y(n_446) );
INVxp67_ASAP7_75t_L g511 ( .A(n_312), .Y(n_511) );
INVx1_ASAP7_75t_L g1951 ( .A(n_313), .Y(n_1951) );
INVx1_ASAP7_75t_L g1543 ( .A(n_314), .Y(n_1543) );
INVx1_ASAP7_75t_L g1226 ( .A(n_316), .Y(n_1226) );
INVx1_ASAP7_75t_L g1536 ( .A(n_317), .Y(n_1536) );
INVxp33_ASAP7_75t_L g799 ( .A(n_318), .Y(n_799) );
INVx1_ASAP7_75t_L g812 ( .A(n_319), .Y(n_812) );
INVx1_ASAP7_75t_L g1423 ( .A(n_320), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_321), .B(n_1673), .Y(n_1672) );
INVx1_ASAP7_75t_L g1679 ( .A(n_321), .Y(n_1679) );
INVx1_ASAP7_75t_L g709 ( .A(n_322), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_323), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g1271 ( .A(n_324), .B(n_1272), .Y(n_1271) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_325), .A2(n_374), .B1(n_1499), .B2(n_1502), .Y(n_1498) );
OAI22xp33_ASAP7_75t_L g1581 ( .A1(n_325), .A2(n_374), .B1(n_1582), .B2(n_1584), .Y(n_1581) );
INVx1_ASAP7_75t_L g1330 ( .A(n_328), .Y(n_1330) );
AOI221xp5_ASAP7_75t_L g1343 ( .A1(n_328), .A2(n_375), .B1(n_807), .B2(n_1344), .C(n_1345), .Y(n_1343) );
INVx1_ASAP7_75t_L g1949 ( .A(n_329), .Y(n_1949) );
XOR2x2_ASAP7_75t_L g382 ( .A(n_330), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g1070 ( .A(n_331), .Y(n_1070) );
INVx1_ASAP7_75t_L g997 ( .A(n_332), .Y(n_997) );
INVx1_ASAP7_75t_L g897 ( .A(n_333), .Y(n_897) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_334), .Y(n_1395) );
INVx1_ASAP7_75t_L g1481 ( .A(n_337), .Y(n_1481) );
INVxp67_ASAP7_75t_SL g1637 ( .A(n_338), .Y(n_1637) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_341), .A2(n_351), .B1(n_727), .B2(n_940), .Y(n_1110) );
INVx1_ASAP7_75t_L g774 ( .A(n_342), .Y(n_774) );
INVx1_ASAP7_75t_L g595 ( .A(n_343), .Y(n_595) );
OAI211xp5_ASAP7_75t_L g1884 ( .A1(n_344), .A2(n_1885), .B(n_1886), .C(n_1887), .Y(n_1884) );
INVx1_ASAP7_75t_L g1902 ( .A(n_344), .Y(n_1902) );
INVx1_ASAP7_75t_L g1515 ( .A(n_345), .Y(n_1515) );
INVx1_ASAP7_75t_L g435 ( .A(n_346), .Y(n_435) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_347), .Y(n_488) );
INVxp67_ASAP7_75t_SL g1597 ( .A(n_348), .Y(n_1597) );
INVx1_ASAP7_75t_L g580 ( .A(n_349), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g1240 ( .A(n_350), .Y(n_1240) );
AOI21xp33_ASAP7_75t_L g1165 ( .A1(n_353), .A2(n_758), .B(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1610 ( .A(n_355), .Y(n_1610) );
INVx1_ASAP7_75t_L g1018 ( .A(n_356), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1186 ( .A(n_357), .Y(n_1186) );
INVx2_ASAP7_75t_L g473 ( .A(n_361), .Y(n_473) );
INVx1_ASAP7_75t_L g482 ( .A(n_361), .Y(n_482) );
INVx1_ASAP7_75t_L g551 ( .A(n_361), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g1446 ( .A1(n_363), .A2(n_364), .B1(n_687), .B2(n_758), .C(n_1158), .Y(n_1446) );
INVx1_ASAP7_75t_L g1153 ( .A(n_365), .Y(n_1153) );
INVx1_ASAP7_75t_L g1229 ( .A(n_366), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_367), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_368), .Y(n_754) );
OAI21xp33_ASAP7_75t_SL g571 ( .A1(n_369), .A2(n_477), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g576 ( .A(n_369), .Y(n_576) );
INVx1_ASAP7_75t_L g1955 ( .A(n_370), .Y(n_1955) );
INVx1_ASAP7_75t_L g1606 ( .A(n_372), .Y(n_1606) );
INVx1_ASAP7_75t_L g1538 ( .A(n_373), .Y(n_1538) );
INVx1_ASAP7_75t_L g1321 ( .A(n_375), .Y(n_1321) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_1648), .B(n_1661), .Y(n_376) );
XNOR2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_884), .Y(n_377) );
XNOR2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_748), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
XNOR2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_635), .Y(n_380) );
XNOR2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_569), .Y(n_381) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_491), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_453), .B(n_470), .C(n_474), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_400), .C(n_417), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g547 ( .A1(n_386), .A2(n_462), .B1(n_548), .B2(n_554), .C1(n_560), .C2(n_562), .Y(n_547) );
INVx2_ASAP7_75t_L g1117 ( .A(n_387), .Y(n_1117) );
AOI211xp5_ASAP7_75t_SL g1126 ( .A1(n_387), .A2(n_1127), .B(n_1128), .C(n_1129), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_387), .A2(n_1014), .B1(n_1208), .B2(n_1214), .C(n_1215), .Y(n_1213) );
AOI221xp5_ASAP7_75t_L g1247 ( .A1(n_387), .A2(n_1014), .B1(n_1248), .B2(n_1249), .C(n_1254), .Y(n_1247) );
AOI211xp5_ASAP7_75t_SL g1339 ( .A1(n_387), .A2(n_1335), .B(n_1340), .C(n_1341), .Y(n_1339) );
AOI211xp5_ASAP7_75t_SL g1366 ( .A1(n_387), .A2(n_1367), .B(n_1368), .C(n_1369), .Y(n_1366) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x6_ASAP7_75t_L g701 ( .A(n_388), .B(n_702), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_389), .B(n_395), .Y(n_388) );
INVx8_ASAP7_75t_L g425 ( .A(n_389), .Y(n_425) );
BUFx3_ASAP7_75t_L g451 ( .A(n_389), .Y(n_451) );
AND2x2_ASAP7_75t_L g465 ( .A(n_389), .B(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g720 ( .A(n_389), .Y(n_720) );
HB1xp67_ASAP7_75t_L g1458 ( .A(n_389), .Y(n_1458) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
AND2x4_ASAP7_75t_L g433 ( .A(n_390), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_391), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_391), .B(n_411), .Y(n_440) );
AND2x4_ASAP7_75t_L g469 ( .A(n_391), .B(n_410), .Y(n_469) );
OR2x2_ASAP7_75t_L g594 ( .A(n_391), .B(n_393), .Y(n_594) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
AND2x6_ASAP7_75t_L g402 ( .A(n_395), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g407 ( .A(n_395), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
AND2x4_ASAP7_75t_L g708 ( .A(n_395), .B(n_550), .Y(n_708) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_396), .B(n_429), .Y(n_428) );
NAND3x1_ASAP7_75t_L g734 ( .A(n_396), .B(n_429), .C(n_735), .Y(n_734) );
OR2x4_ASAP7_75t_L g1501 ( .A(n_396), .B(n_594), .Y(n_1501) );
INVx1_ASAP7_75t_L g1504 ( .A(n_396), .Y(n_1504) );
AND2x4_ASAP7_75t_L g1509 ( .A(n_396), .B(n_469), .Y(n_1509) );
OR2x6_ASAP7_75t_L g1525 ( .A(n_396), .B(n_811), .Y(n_1525) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g449 ( .A(n_397), .B(n_399), .Y(n_449) );
BUFx3_ASAP7_75t_L g589 ( .A(n_397), .Y(n_589) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g588 ( .A(n_399), .B(n_589), .Y(n_588) );
AND3x4_ASAP7_75t_L g715 ( .A(n_399), .B(n_472), .C(n_589), .Y(n_715) );
HB1xp67_ASAP7_75t_L g1494 ( .A(n_399), .Y(n_1494) );
INVx4_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_402), .A2(n_407), .B1(n_580), .B2(n_581), .Y(n_579) );
AND2x2_ASAP7_75t_L g707 ( .A(n_403), .B(n_708), .Y(n_707) );
NAND2x1_ASAP7_75t_L g825 ( .A(n_403), .B(n_708), .Y(n_825) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_403), .B(n_708), .Y(n_1468) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_405), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g452 ( .A(n_405), .B(n_409), .Y(n_452) );
BUFx2_ASAP7_75t_L g1514 ( .A(n_405), .Y(n_1514) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_407), .Y(n_1103) );
INVx1_ASAP7_75t_L g712 ( .A(n_408), .Y(n_712) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_411), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_412), .Y(n_1104) );
OR2x6_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g1143 ( .A(n_413), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1239 ( .A1(n_413), .A2(n_427), .B1(n_802), .B2(n_1240), .C(n_1241), .Y(n_1239) );
INVx1_ASAP7_75t_L g1387 ( .A(n_413), .Y(n_1387) );
INVx1_ASAP7_75t_L g1507 ( .A(n_413), .Y(n_1507) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_414), .Y(n_422) );
BUFx3_ASAP7_75t_L g990 ( .A(n_414), .Y(n_990) );
BUFx2_ASAP7_75t_L g1518 ( .A(n_415), .Y(n_1518) );
INVx1_ASAP7_75t_L g1027 ( .A(n_416), .Y(n_1027) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_430), .B(n_442), .Y(n_417) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_423), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_419), .A2(n_443), .B1(n_519), .B2(n_520), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_420), .A2(n_427), .B1(n_599), .B2(n_600), .C(n_601), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g1045 ( .A1(n_420), .A2(n_588), .B1(n_1046), .B2(n_1047), .C(n_1049), .Y(n_1045) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g1036 ( .A(n_421), .Y(n_1036) );
INVx2_ASAP7_75t_L g1135 ( .A(n_421), .Y(n_1135) );
INVx2_ASAP7_75t_L g1347 ( .A(n_421), .Y(n_1347) );
INVx1_ASAP7_75t_L g1928 ( .A(n_421), .Y(n_1928) );
INVx4_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_422), .Y(n_584) );
OR2x2_ASAP7_75t_L g700 ( .A(n_422), .B(n_695), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g1234 ( .A1(n_422), .A2(n_588), .B1(n_1235), .B2(n_1236), .C(n_1237), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1378 ( .A(n_422), .Y(n_1378) );
A2O1A1Ixp33_ASAP7_75t_L g988 ( .A1(n_424), .A2(n_708), .B(n_960), .C(n_989), .Y(n_988) );
INVx8_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g859 ( .A(n_425), .Y(n_859) );
INVx3_ASAP7_75t_L g879 ( .A(n_425), .Y(n_879) );
INVx2_ASAP7_75t_L g1289 ( .A(n_425), .Y(n_1289) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_427), .A2(n_1035), .B1(n_1036), .B2(n_1037), .C(n_1038), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_427), .B(n_1145), .Y(n_1144) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_427), .A2(n_600), .B1(n_990), .B2(n_1186), .C(n_1198), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g1345 ( .A1(n_427), .A2(n_800), .B1(n_1346), .B2(n_1347), .C(n_1348), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_427), .B(n_1389), .Y(n_1388) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_428), .B(n_496), .Y(n_1008) );
OR2x6_ASAP7_75t_L g1465 ( .A(n_428), .B(n_496), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_435), .B1(n_436), .B2(n_441), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g1350 ( .A1(n_431), .A2(n_588), .B1(n_1331), .B2(n_1347), .C(n_1351), .Y(n_1350) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g586 ( .A(n_432), .Y(n_586) );
INVx3_ASAP7_75t_L g730 ( .A(n_432), .Y(n_730) );
AND2x4_ASAP7_75t_L g743 ( .A(n_432), .B(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_432), .Y(n_876) );
BUFx8_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_433), .Y(n_447) );
INVx2_ASAP7_75t_L g459 ( .A(n_433), .Y(n_459) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_433), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_435), .A2(n_511), .B1(n_512), .B2(n_515), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_436), .A2(n_586), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g694 ( .A(n_438), .B(n_695), .Y(n_694) );
BUFx3_ASAP7_75t_L g795 ( .A(n_438), .Y(n_795) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_439), .Y(n_597) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g811 ( .A(n_440), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_441), .A2(n_506), .B1(n_523), .B2(n_525), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_446), .C(n_450), .Y(n_442) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g804 ( .A(n_445), .Y(n_804) );
INVx2_ASAP7_75t_L g1251 ( .A(n_445), .Y(n_1251) );
INVx5_ASAP7_75t_L g873 ( .A(n_447), .Y(n_873) );
INVx2_ASAP7_75t_SL g1023 ( .A(n_447), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_447), .Y(n_1032) );
INVx3_ASAP7_75t_L g1243 ( .A(n_447), .Y(n_1243) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g797 ( .A(n_449), .B(n_530), .Y(n_797) );
INVx1_ASAP7_75t_L g1219 ( .A(n_451), .Y(n_1219) );
AND2x4_ASAP7_75t_L g461 ( .A(n_452), .B(n_457), .Y(n_461) );
BUFx12f_ASAP7_75t_L g727 ( .A(n_452), .Y(n_727) );
INVx5_ASAP7_75t_L g732 ( .A(n_452), .Y(n_732) );
BUFx3_ASAP7_75t_L g874 ( .A(n_452), .Y(n_874) );
BUFx3_ASAP7_75t_L g1017 ( .A(n_452), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1344 ( .A(n_452), .Y(n_1344) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_460), .B1(n_461), .B2(n_462), .C(n_463), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
OR2x6_ASAP7_75t_SL g455 ( .A(n_456), .B(n_459), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_457), .Y(n_1015) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g466 ( .A(n_458), .Y(n_466) );
OR2x2_ASAP7_75t_L g695 ( .A(n_458), .B(n_530), .Y(n_695) );
BUFx2_ASAP7_75t_L g725 ( .A(n_459), .Y(n_725) );
INVx1_ASAP7_75t_L g793 ( .A(n_459), .Y(n_793) );
INVx3_ASAP7_75t_L g925 ( .A(n_459), .Y(n_925) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_459), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_460), .B(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g574 ( .A(n_461), .Y(n_574) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_465), .A2(n_468), .B1(n_576), .B2(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g468 ( .A(n_466), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g722 ( .A(n_469), .Y(n_722) );
BUFx2_ASAP7_75t_L g814 ( .A(n_469), .Y(n_814) );
BUFx2_ASAP7_75t_L g880 ( .A(n_469), .Y(n_880) );
INVx2_ASAP7_75t_L g1020 ( .A(n_469), .Y(n_1020) );
BUFx3_ASAP7_75t_L g1108 ( .A(n_469), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1463 ( .A(n_469), .Y(n_1463) );
BUFx2_ASAP7_75t_L g1617 ( .A(n_469), .Y(n_1617) );
INVx1_ASAP7_75t_L g788 ( .A(n_470), .Y(n_788) );
INVx1_ASAP7_75t_L g1484 ( .A(n_470), .Y(n_1484) );
BUFx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g690 ( .A(n_471), .Y(n_690) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_471), .Y(n_1255) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI31xp33_ASAP7_75t_SL g572 ( .A1(n_472), .A2(n_573), .A3(n_578), .B(n_582), .Y(n_572) );
INVx2_ASAP7_75t_SL g855 ( .A(n_472), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g1098 ( .A1(n_472), .A2(n_1099), .B1(n_1118), .B2(n_1120), .Y(n_1098) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g496 ( .A(n_473), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_473), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_478), .A2(n_564), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_478), .B(n_1078), .Y(n_1077) );
AOI211xp5_ASAP7_75t_L g1149 ( .A1(n_478), .A2(n_1150), .B(n_1151), .C(n_1155), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_478), .B(n_1211), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_478), .B(n_1253), .Y(n_1256) );
AO211x2_ASAP7_75t_L g1363 ( .A1(n_478), .A2(n_1364), .B(n_1365), .C(n_1392), .Y(n_1363) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
AND2x4_ASAP7_75t_L g564 ( .A(n_479), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g541 ( .A(n_480), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g613 ( .A(n_480), .B(n_542), .Y(n_613) );
INVxp67_ASAP7_75t_L g702 ( .A(n_480), .Y(n_702) );
INVx1_ASAP7_75t_L g1589 ( .A(n_480), .Y(n_1589) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g530 ( .A(n_481), .Y(n_530) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_483), .Y(n_660) );
INVx1_ASAP7_75t_L g770 ( .A(n_483), .Y(n_770) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_484), .B(n_551), .Y(n_556) );
AND2x2_ASAP7_75t_L g565 ( .A(n_484), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g640 ( .A(n_484), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g664 ( .A(n_484), .B(n_566), .Y(n_664) );
AND2x4_ASAP7_75t_SL g669 ( .A(n_484), .B(n_618), .Y(n_669) );
BUFx2_ASAP7_75t_L g962 ( .A(n_484), .Y(n_962) );
HB1xp67_ASAP7_75t_L g1577 ( .A(n_485), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_486), .B(n_537), .Y(n_553) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_486), .Y(n_621) );
INVx3_ASAP7_75t_L g631 ( .A(n_486), .Y(n_631) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
OR2x2_ASAP7_75t_L g514 ( .A(n_487), .B(n_490), .Y(n_514) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g504 ( .A(n_488), .B(n_490), .Y(n_504) );
INVx2_ASAP7_75t_L g509 ( .A(n_488), .Y(n_509) );
NAND2x1_ASAP7_75t_L g517 ( .A(n_488), .B(n_490), .Y(n_517) );
INVx1_ASAP7_75t_L g544 ( .A(n_488), .Y(n_544) );
AND2x2_ASAP7_75t_L g567 ( .A(n_488), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g619 ( .A(n_488), .B(n_490), .Y(n_619) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_490), .B(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g540 ( .A(n_490), .Y(n_540) );
AND2x2_ASAP7_75t_L g559 ( .A(n_490), .B(n_509), .Y(n_559) );
INVx2_ASAP7_75t_L g568 ( .A(n_490), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_547), .C(n_563), .Y(n_491) );
NOR2xp33_ASAP7_75t_SL g492 ( .A(n_493), .B(n_531), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_499), .A3(n_510), .B1(n_518), .B2(n_522), .B3(n_526), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g1183 ( .A1(n_494), .A2(n_1184), .A3(n_1188), .B1(n_1194), .B2(n_1199), .B3(n_1204), .Y(n_1183) );
OAI22xp5_ASAP7_75t_SL g1262 ( .A1(n_494), .A2(n_1263), .B1(n_1266), .B2(n_1267), .Y(n_1262) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx4_ASAP7_75t_L g623 ( .A(n_495), .Y(n_623) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_495), .Y(n_1053) );
AOI31xp33_ASAP7_75t_L g1085 ( .A1(n_495), .A2(n_607), .A3(n_1086), .B(n_1087), .Y(n_1085) );
INVx2_ASAP7_75t_L g1166 ( .A(n_495), .Y(n_1166) );
INVx2_ASAP7_75t_L g1529 ( .A(n_495), .Y(n_1529) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g919 ( .A(n_496), .Y(n_919) );
AND2x4_ASAP7_75t_L g528 ( .A(n_498), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g689 ( .A(n_498), .Y(n_689) );
BUFx2_ASAP7_75t_L g1568 ( .A(n_498), .Y(n_1568) );
AND2x4_ASAP7_75t_L g1572 ( .A(n_498), .B(n_543), .Y(n_1572) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_505), .B2(n_506), .Y(n_499) );
INVx2_ASAP7_75t_L g1328 ( .A(n_501), .Y(n_1328) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g524 ( .A(n_502), .Y(n_524) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_502), .Y(n_1056) );
BUFx3_ASAP7_75t_L g1171 ( .A(n_502), .Y(n_1171) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx4f_ASAP7_75t_L g678 ( .A(n_503), .Y(n_678) );
INVx2_ASAP7_75t_L g1162 ( .A(n_503), .Y(n_1162) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx8_ASAP7_75t_L g681 ( .A(n_507), .Y(n_681) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_507), .B(n_1568), .Y(n_1580) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_512), .A2(n_1033), .B1(n_1046), .B2(n_1060), .C(n_1062), .Y(n_1059) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g519 ( .A(n_514), .Y(n_519) );
INVx2_ASAP7_75t_L g835 ( .A(n_514), .Y(n_835) );
BUFx3_ASAP7_75t_L g901 ( .A(n_514), .Y(n_901) );
BUFx2_ASAP7_75t_L g958 ( .A(n_514), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_515), .A2(n_1030), .B1(n_1040), .B2(n_1056), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_515), .A2(n_1195), .B1(n_1197), .B2(n_1198), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1561 ( .A(n_515), .Y(n_1561) );
BUFx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g561 ( .A(n_516), .B(n_556), .Y(n_561) );
INVx2_ASAP7_75t_SL g832 ( .A(n_516), .Y(n_832) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_516), .B(n_556), .Y(n_1068) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_517), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_520), .A2(n_834), .B1(n_1235), .B2(n_1240), .C(n_1268), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_520), .A2(n_1538), .B1(n_1539), .B2(n_1540), .Y(n_1537) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x6_ASAP7_75t_L g545 ( .A(n_521), .B(n_546), .Y(n_545) );
BUFx4f_ASAP7_75t_L g896 ( .A(n_521), .Y(n_896) );
INVx4_ASAP7_75t_L g1191 ( .A(n_521), .Y(n_1191) );
BUFx4f_ASAP7_75t_L g1264 ( .A(n_521), .Y(n_1264) );
BUFx4f_ASAP7_75t_L g1896 ( .A(n_521), .Y(n_1896) );
BUFx4f_ASAP7_75t_L g1964 ( .A(n_521), .Y(n_1964) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_523), .A2(n_839), .B1(n_840), .B2(n_843), .Y(n_838) );
OAI221xp5_ASAP7_75t_L g1625 ( .A1(n_523), .A2(n_1606), .B1(n_1615), .B2(n_1626), .C(n_1628), .Y(n_1625) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g1204 ( .A(n_527), .Y(n_1204) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_528), .B(n_530), .Y(n_527) );
AND2x4_ASAP7_75t_L g626 ( .A(n_528), .B(n_627), .Y(n_626) );
INVx4_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
INVx4_ASAP7_75t_L g850 ( .A(n_528), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_528), .B(n_627), .Y(n_1266) );
AND2x4_ASAP7_75t_L g688 ( .A(n_529), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g1588 ( .A(n_529), .Y(n_1588) );
INVx1_ASAP7_75t_L g628 ( .A(n_530), .Y(n_628) );
HB1xp67_ASAP7_75t_L g1496 ( .A(n_530), .Y(n_1496) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g1090 ( .A(n_534), .Y(n_1090) );
NAND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_537), .B(n_543), .Y(n_542) );
AND2x6_ASAP7_75t_L g656 ( .A(n_537), .B(n_618), .Y(n_656) );
INVx1_ASAP7_75t_L g674 ( .A(n_537), .Y(n_674) );
AND2x2_ASAP7_75t_L g766 ( .A(n_537), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g673 ( .A(n_540), .Y(n_673) );
BUFx2_ASAP7_75t_L g767 ( .A(n_540), .Y(n_767) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_540), .B(n_1568), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1899 ( .A(n_540), .B(n_1568), .Y(n_1899) );
INVx1_ASAP7_75t_L g971 ( .A(n_542), .Y(n_971) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_545), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g1057 ( .A1(n_545), .A2(n_1058), .B(n_1059), .Y(n_1057) );
AOI332xp33_ASAP7_75t_L g614 ( .A1(n_548), .A2(n_615), .A3(n_620), .B1(n_622), .B2(n_624), .B3(n_626), .C1(n_629), .C2(n_633), .Y(n_614) );
AOI322xp5_ASAP7_75t_L g1156 ( .A1(n_548), .A2(n_626), .A3(n_1157), .B1(n_1159), .B2(n_1165), .C1(n_1167), .C2(n_1168), .Y(n_1156) );
AOI222xp33_ASAP7_75t_L g1206 ( .A1(n_548), .A2(n_554), .B1(n_560), .B2(n_1207), .C1(n_1208), .C2(n_1209), .Y(n_1206) );
AOI222xp33_ASAP7_75t_L g1334 ( .A1(n_548), .A2(n_554), .B1(n_560), .B2(n_1335), .C1(n_1336), .C2(n_1337), .Y(n_1334) );
AOI21xp33_ASAP7_75t_L g1411 ( .A1(n_548), .A2(n_607), .B(n_1412), .Y(n_1411) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
AOI332xp33_ASAP7_75t_L g1258 ( .A1(n_549), .A2(n_552), .A3(n_555), .B1(n_557), .B2(n_560), .B3(n_1248), .C1(n_1259), .C2(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g696 ( .A(n_550), .B(n_553), .Y(n_696) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g735 ( .A(n_551), .Y(n_735) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_554), .A2(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g1067 ( .A(n_554), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_554), .A2(n_560), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g632 ( .A(n_559), .Y(n_632) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_559), .Y(n_641) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_559), .Y(n_1088) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_560), .A2(n_581), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_564), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g1119 ( .A(n_564), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_564), .B(n_1147), .Y(n_1146) );
NAND2xp33_ASAP7_75t_SL g1225 ( .A(n_564), .B(n_1226), .Y(n_1225) );
HB1xp67_ASAP7_75t_L g1355 ( .A(n_564), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_564), .B(n_1391), .Y(n_1390) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
INVx2_ASAP7_75t_L g761 ( .A(n_566), .Y(n_761) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx3_ASAP7_75t_L g645 ( .A(n_567), .Y(n_645) );
INVx2_ASAP7_75t_L g780 ( .A(n_567), .Y(n_780) );
AND2x4_ASAP7_75t_L g1585 ( .A(n_567), .B(n_1577), .Y(n_1585) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_634), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_605), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_590), .B1(n_598), .B2(n_602), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_586), .B2(n_587), .C(n_588), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_584), .A2(n_802), .B1(n_994), .B2(n_995), .Y(n_993) );
HB1xp67_ASAP7_75t_L g1553 ( .A(n_584), .Y(n_1553) );
OAI22xp33_ASAP7_75t_L g1943 ( .A1(n_584), .A2(n_800), .B1(n_1944), .B2(n_1945), .Y(n_1943) );
INVx1_ASAP7_75t_L g940 ( .A(n_586), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_588), .A2(n_719), .B1(n_732), .B2(n_1137), .C(n_1138), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g1220 ( .A1(n_588), .A2(n_990), .B1(n_1002), .B2(n_1193), .C(n_1197), .Y(n_1220) );
INVx1_ASAP7_75t_L g1380 ( .A(n_588), .Y(n_1380) );
INVx3_ASAP7_75t_L g1513 ( .A(n_589), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_595), .B2(n_596), .Y(n_590) );
BUFx4f_ASAP7_75t_SL g1041 ( .A(n_592), .Y(n_1041) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g739 ( .A(n_593), .Y(n_739) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx3_ASAP7_75t_L g600 ( .A(n_594), .Y(n_600) );
BUFx4f_ASAP7_75t_L g802 ( .A(n_594), .Y(n_802) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_594), .Y(n_1037) );
OR2x4_ASAP7_75t_L g1522 ( .A(n_594), .B(n_1504), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_596), .A2(n_730), .B1(n_1189), .B2(n_1203), .Y(n_1223) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
CKINVDCx8_ASAP7_75t_R g1114 ( .A(n_597), .Y(n_1114) );
INVx3_ASAP7_75t_L g1245 ( .A(n_597), .Y(n_1245) );
INVx3_ASAP7_75t_L g1555 ( .A(n_597), .Y(n_1555) );
INVx1_ASAP7_75t_L g1386 ( .A(n_600), .Y(n_1386) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_606), .B(n_608), .C(n_610), .D(n_614), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g1261 ( .A(n_607), .B(n_1262), .C(n_1269), .Y(n_1261) );
NOR3xp33_ASAP7_75t_L g1317 ( .A(n_607), .B(n_1318), .C(n_1319), .Y(n_1317) );
AND2x4_ASAP7_75t_L g699 ( .A(n_613), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g921 ( .A(n_613), .B(n_700), .Y(n_921) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_613), .Y(n_1092) );
BUFx3_ASAP7_75t_L g1158 ( .A(n_616), .Y(n_1158) );
BUFx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx3_ASAP7_75t_L g625 ( .A(n_618), .Y(n_625) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_618), .Y(n_648) );
BUFx3_ASAP7_75t_L g758 ( .A(n_618), .Y(n_758) );
BUFx3_ASAP7_75t_L g776 ( .A(n_618), .Y(n_776) );
INVx1_ASAP7_75t_L g912 ( .A(n_618), .Y(n_912) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_618), .B(n_1564), .Y(n_1563) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g686 ( .A(n_619), .Y(n_686) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_621), .Y(n_653) );
INVx3_ASAP7_75t_L g966 ( .A(n_621), .Y(n_966) );
INVx1_ASAP7_75t_L g1912 ( .A(n_622), .Y(n_1912) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g1402 ( .A(n_623), .Y(n_1402) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_626), .Y(n_1058) );
NAND3xp33_ASAP7_75t_L g1094 ( .A(n_626), .B(n_1095), .C(n_1096), .Y(n_1094) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g764 ( .A(n_631), .Y(n_764) );
INVx2_ASAP7_75t_L g1300 ( .A(n_631), .Y(n_1300) );
INVx1_ASAP7_75t_L g1304 ( .A(n_631), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_632), .Y(n_765) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_632), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_632), .A2(n_758), .B1(n_960), .B2(n_961), .Y(n_959) );
BUFx3_ASAP7_75t_L g1301 ( .A(n_632), .Y(n_1301) );
NAND3xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_691), .C(n_703), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_665), .B(n_690), .Y(n_637) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_640), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g1297 ( .A1(n_640), .A2(n_656), .B1(n_1274), .B2(n_1298), .C(n_1299), .Y(n_1297) );
AOI221xp5_ASAP7_75t_L g1475 ( .A1(n_640), .A2(n_656), .B1(n_1453), .B2(n_1476), .C(n_1478), .Y(n_1475) );
INVx1_ASAP7_75t_L g655 ( .A(n_641), .Y(n_655) );
BUFx2_ASAP7_75t_L g979 ( .A(n_641), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_651), .B(n_656), .Y(n_642) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_648), .Y(n_1169) );
HB1xp67_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_656), .A2(n_773), .B1(n_774), .B2(n_775), .C(n_781), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_656), .A2(n_847), .B(n_851), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_656), .A2(n_910), .B(n_913), .Y(n_909) );
AOI21xp5_ASAP7_75t_SL g1434 ( .A1(n_656), .A2(n_1435), .B(n_1439), .Y(n_1434) );
INVx1_ASAP7_75t_L g1630 ( .A(n_656), .Y(n_1630) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_661), .B2(n_662), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g1294 ( .A1(n_659), .A2(n_784), .B1(n_1295), .B2(n_1296), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_660), .A2(n_784), .B1(n_853), .B2(n_854), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_660), .A2(n_664), .B1(n_915), .B2(n_916), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1480 ( .A1(n_660), .A2(n_664), .B1(n_1481), .B2(n_1482), .Y(n_1480) );
INVx1_ASAP7_75t_L g1640 ( .A(n_660), .Y(n_1640) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_662), .A2(n_769), .B1(n_1422), .B2(n_1423), .Y(n_1440) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_664), .Y(n_784) );
HB1xp67_ASAP7_75t_L g1633 ( .A(n_664), .Y(n_1633) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g894 ( .A(n_667), .Y(n_894) );
INVx1_ASAP7_75t_L g1442 ( .A(n_667), .Y(n_1442) );
INVx4_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g773 ( .A(n_669), .Y(n_773) );
BUFx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g844 ( .A(n_672), .Y(n_844) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g968 ( .A(n_674), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B1(n_680), .B2(n_682), .C(n_683), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g1443 ( .A1(n_676), .A2(n_1060), .B1(n_1444), .B2(n_1445), .C(n_1446), .Y(n_1443) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g904 ( .A(n_677), .Y(n_904) );
INVx2_ASAP7_75t_SL g1547 ( .A(n_677), .Y(n_1547) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g955 ( .A(n_678), .Y(n_955) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g842 ( .A(n_681), .Y(n_842) );
INVx1_ASAP7_75t_L g907 ( .A(n_681), .Y(n_907) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_681), .Y(n_1061) );
INVx2_ASAP7_75t_L g1173 ( .A(n_681), .Y(n_1173) );
INVx2_ASAP7_75t_SL g1187 ( .A(n_681), .Y(n_1187) );
INVx4_ASAP7_75t_L g1323 ( .A(n_681), .Y(n_1323) );
INVx2_ASAP7_75t_L g1916 ( .A(n_681), .Y(n_1916) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g1438 ( .A(n_685), .Y(n_1438) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g762 ( .A(n_688), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g895 ( .A1(n_688), .A2(n_896), .B1(n_897), .B2(n_898), .C(n_899), .Y(n_895) );
INVx3_ASAP7_75t_L g975 ( .A(n_688), .Y(n_975) );
INVx1_ASAP7_75t_L g1309 ( .A(n_688), .Y(n_1309) );
INVx1_ASAP7_75t_L g1564 ( .A(n_689), .Y(n_1564) );
INVxp67_ASAP7_75t_L g1583 ( .A(n_689), .Y(n_1583) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_697), .B(n_698), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_692), .A2(n_786), .B1(n_820), .B2(n_821), .C(n_822), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_692), .B(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_692), .B(n_928), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_692), .A2(n_820), .B1(n_1274), .B2(n_1275), .C(n_1276), .Y(n_1273) );
AOI221xp5_ASAP7_75t_L g1452 ( .A1(n_692), .A2(n_820), .B1(n_1453), .B2(n_1454), .C(n_1455), .Y(n_1452) );
AOI21xp5_ASAP7_75t_L g1620 ( .A1(n_692), .A2(n_1621), .B(n_1622), .Y(n_1620) );
INVx8_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g741 ( .A(n_695), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_695), .Y(n_744) );
INVx1_ASAP7_75t_L g1066 ( .A(n_696), .Y(n_1066) );
INVx2_ASAP7_75t_L g753 ( .A(n_699), .Y(n_753) );
INVx2_ASAP7_75t_L g985 ( .A(n_700), .Y(n_985) );
INVx3_ASAP7_75t_L g820 ( .A(n_701), .Y(n_820) );
INVx5_ASAP7_75t_L g868 ( .A(n_701), .Y(n_868) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_737), .C(n_745), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_713), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_709), .B2(n_710), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_707), .A2(n_710), .B1(n_864), .B2(n_865), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_707), .A2(n_710), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_707), .A2(n_710), .B1(n_1419), .B2(n_1420), .Y(n_1418) );
AND2x4_ASAP7_75t_L g710 ( .A(n_708), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g747 ( .A(n_708), .B(n_722), .Y(n_747) );
AND2x4_ASAP7_75t_SL g933 ( .A(n_708), .B(n_711), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_710), .A2(n_768), .B1(n_774), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_710), .A2(n_1467), .B1(n_1468), .B2(n_1469), .Y(n_1466) );
INVx1_ASAP7_75t_L g1601 ( .A(n_710), .Y(n_1601) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI33xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .A3(n_723), .B1(n_728), .B2(n_733), .B3(n_736), .Y(n_713) );
AOI33xp33_ASAP7_75t_L g869 ( .A1(n_714), .A2(n_870), .A3(n_871), .B1(n_875), .B2(n_877), .B3(n_878), .Y(n_869) );
INVx1_ASAP7_75t_L g1290 ( .A(n_714), .Y(n_1290) );
AOI33xp33_ASAP7_75t_L g1424 ( .A1(n_714), .A2(n_733), .A3(n_1425), .B1(n_1427), .B2(n_1428), .B3(n_1430), .Y(n_1424) );
BUFx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI33xp33_ASAP7_75t_L g936 ( .A1(n_715), .A2(n_937), .A3(n_938), .B1(n_939), .B2(n_941), .B3(n_942), .Y(n_936) );
AOI33xp33_ASAP7_75t_L g1456 ( .A1(n_715), .A2(n_1457), .A3(n_1459), .B1(n_1461), .B2(n_1462), .B3(n_1464), .Y(n_1456) );
BUFx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_720), .B(n_1253), .Y(n_1252) );
BUFx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_722), .A2(n_879), .B1(n_1078), .B2(n_1093), .Y(n_1115) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g1429 ( .A(n_732), .Y(n_1429) );
INVx2_ASAP7_75t_R g1460 ( .A(n_732), .Y(n_1460) );
INVx2_ASAP7_75t_L g1557 ( .A(n_733), .Y(n_1557) );
INVx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_L g817 ( .A(n_734), .Y(n_817) );
OR2x6_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g1558 ( .A1(n_739), .A2(n_804), .B1(n_1536), .B2(n_1543), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1619 ( .A(n_739), .B(n_740), .Y(n_1619) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g924 ( .A(n_741), .B(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g818 ( .A(n_743), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_743), .A2(n_853), .B1(n_854), .B2(n_858), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_743), .A2(n_858), .B1(n_1295), .B2(n_1296), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_743), .A2(n_858), .B1(n_1422), .B2(n_1423), .Y(n_1421) );
AND2x4_ASAP7_75t_L g858 ( .A(n_744), .B(n_859), .Y(n_858) );
AND2x4_ASAP7_75t_L g923 ( .A(n_744), .B(n_859), .Y(n_923) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
NAND3xp33_ASAP7_75t_SL g1276 ( .A(n_746), .B(n_1277), .C(n_1280), .Y(n_1276) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g881 ( .A(n_747), .Y(n_881) );
NOR3xp33_ASAP7_75t_L g1416 ( .A(n_747), .B(n_1417), .C(n_1431), .Y(n_1416) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_826), .B1(n_882), .B2(n_883), .Y(n_748) );
INVx1_ASAP7_75t_L g882 ( .A(n_749), .Y(n_882) );
XNOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_819), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_787), .C(n_789), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_772), .C(n_783), .Y(n_755) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_763), .B1(n_766), .B2(n_768), .C1(n_769), .C2(n_771), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g964 ( .A1(n_758), .A2(n_965), .B(n_967), .C(n_968), .Y(n_964) );
BUFx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g1308 ( .A(n_761), .Y(n_1308) );
INVx1_ASAP7_75t_L g837 ( .A(n_762), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g969 ( .A1(n_766), .A2(n_970), .B1(n_971), .B2(n_972), .Y(n_969) );
INVx1_ASAP7_75t_L g1311 ( .A(n_766), .Y(n_1311) );
AOI222xp33_ASAP7_75t_L g1472 ( .A1(n_766), .A2(n_773), .B1(n_1467), .B2(n_1469), .C1(n_1473), .C2(n_1474), .Y(n_1472) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI222xp33_ASAP7_75t_L g1302 ( .A1(n_773), .A2(n_1278), .B1(n_1279), .B2(n_1303), .C1(n_1305), .C2(n_1310), .Y(n_1302) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g849 ( .A(n_779), .Y(n_849) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g1477 ( .A(n_780), .Y(n_1477) );
A2O1A1Ixp33_ASAP7_75t_SL g1338 ( .A1(n_787), .A2(n_1339), .B(n_1342), .C(n_1353), .Y(n_1338) );
OAI21xp5_ASAP7_75t_L g1432 ( .A1(n_787), .A2(n_1433), .B(n_1441), .Y(n_1432) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B1(n_794), .B2(n_795), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g1605 ( .A(n_793), .Y(n_1605) );
OAI22xp5_ASAP7_75t_L g1950 ( .A1(n_795), .A2(n_1283), .B1(n_1951), .B2(n_1952), .Y(n_1950) );
OAI33xp33_ASAP7_75t_L g1926 ( .A1(n_796), .A2(n_1618), .A3(n_1927), .B1(n_1929), .B2(n_1930), .B3(n_1931), .Y(n_1926) );
BUFx8_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx4f_ASAP7_75t_L g992 ( .A(n_797), .Y(n_992) );
BUFx2_ASAP7_75t_L g1942 ( .A(n_797), .Y(n_1942) );
OAI22xp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_803), .B2(n_804), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g1953 ( .A1(n_800), .A2(n_1609), .B1(n_1954), .B2(n_1955), .Y(n_1953) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_802), .A2(n_990), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_809), .B1(n_810), .B2(n_812), .C(n_813), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g1374 ( .A(n_807), .Y(n_1374) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx6f_ASAP7_75t_L g1048 ( .A(n_808), .Y(n_1048) );
INVx2_ASAP7_75t_L g1113 ( .A(n_808), .Y(n_1113) );
INVx1_ASAP7_75t_L g1133 ( .A(n_808), .Y(n_1133) );
INVx2_ASAP7_75t_L g1237 ( .A(n_808), .Y(n_1237) );
AND2x4_ASAP7_75t_L g1503 ( .A(n_808), .B(n_1504), .Y(n_1503) );
INVx2_ASAP7_75t_L g1948 ( .A(n_808), .Y(n_1948) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_810), .A2(n_1030), .B1(n_1031), .B2(n_1033), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_810), .A2(n_1002), .B1(n_1540), .B2(n_1549), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g1603 ( .A1(n_810), .A2(n_1604), .B1(n_1605), .B2(n_1606), .Y(n_1603) );
OAI221xp5_ASAP7_75t_L g1611 ( .A1(n_810), .A2(n_1612), .B1(n_1613), .B2(n_1615), .C(n_1616), .Y(n_1611) );
BUFx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g999 ( .A(n_811), .Y(n_999) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
BUFx2_ASAP7_75t_L g877 ( .A(n_817), .Y(n_877) );
BUFx2_ASAP7_75t_L g942 ( .A(n_817), .Y(n_942) );
BUFx2_ASAP7_75t_L g1286 ( .A(n_817), .Y(n_1286) );
INVxp67_ASAP7_75t_L g1598 ( .A(n_818), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_820), .B(n_935), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_824), .A2(n_931), .B1(n_932), .B2(n_933), .Y(n_930) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g883 ( .A(n_826), .Y(n_883) );
NAND3x1_ASAP7_75t_L g827 ( .A(n_828), .B(n_860), .C(n_862), .Y(n_827) );
O2A1O1Ixp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_845), .B(n_855), .C(n_856), .Y(n_828) );
OAI221xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_833), .B1(n_834), .B2(n_836), .C(n_837), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g1541 ( .A1(n_831), .A2(n_1539), .B1(n_1542), .B2(n_1543), .Y(n_1541) );
INVx5_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_835), .Y(n_1196) );
INVx2_ASAP7_75t_L g1961 ( .A(n_835), .Y(n_1961) );
BUFx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVxp33_ASAP7_75t_L g1333 ( .A(n_842), .Y(n_1333) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g1097 ( .A(n_849), .Y(n_1097) );
A2O1A1Ixp33_ASAP7_75t_L g1125 ( .A1(n_855), .A2(n_1126), .B(n_1130), .C(n_1146), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_858), .B(n_982), .Y(n_981) );
AND4x1_ASAP7_75t_SL g862 ( .A(n_863), .B(n_866), .C(n_869), .D(n_881), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx8_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_873), .A2(n_997), .B1(n_998), .B2(n_1000), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1930 ( .A1(n_873), .A2(n_1043), .B1(n_1919), .B2(n_1925), .Y(n_1930) );
INVx1_ASAP7_75t_L g1618 ( .A(n_877), .Y(n_1618) );
A2O1A1Ixp33_ASAP7_75t_L g1024 ( .A1(n_879), .A2(n_1025), .B(n_1026), .C(n_1027), .Y(n_1024) );
AND4x1_ASAP7_75t_L g929 ( .A(n_881), .B(n_930), .C(n_934), .D(n_936), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g1455 ( .A(n_881), .B(n_1456), .C(n_1466), .Y(n_1455) );
AOI22x1_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_1359), .B1(n_1646), .B2(n_1647), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AO22x2_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_943), .B2(n_944), .Y(n_886) );
AO22x1_ASAP7_75t_L g1647 ( .A1(n_887), .A2(n_888), .B1(n_943), .B2(n_944), .Y(n_1647) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NOR2x1p5_ASAP7_75t_L g890 ( .A(n_891), .B(n_926), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
O2A1O1Ixp33_ASAP7_75t_SL g892 ( .A1(n_893), .A2(n_908), .B(n_917), .C(n_920), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g1920 ( .A1(n_896), .A2(n_1192), .B1(n_1921), .B2(n_1922), .Y(n_1920) );
OAI221xp5_ASAP7_75t_L g1329 ( .A1(n_899), .A2(n_1264), .B1(n_1330), .B2(n_1331), .C(n_1332), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g1917 ( .A1(n_899), .A2(n_1896), .B1(n_1918), .B2(n_1919), .Y(n_1917) );
OAI22xp5_ASAP7_75t_L g1963 ( .A1(n_899), .A2(n_1945), .B1(n_1955), .B2(n_1964), .Y(n_1963) );
INVx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_901), .A2(n_1236), .B1(n_1244), .B2(n_1264), .C(n_1265), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1546 ( .A1(n_906), .A2(n_1547), .B1(n_1548), .B2(n_1549), .Y(n_1546) );
BUFx3_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g1629 ( .A(n_912), .Y(n_1629) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_915), .A2(n_916), .B1(n_923), .B2(n_924), .Y(n_922) );
OAI31xp33_ASAP7_75t_L g1623 ( .A1(n_917), .A2(n_1624), .A3(n_1631), .B(n_1639), .Y(n_1623) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g1224 ( .A(n_918), .Y(n_1224) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
AOI21xp5_ASAP7_75t_SL g952 ( .A1(n_919), .A2(n_953), .B(n_973), .Y(n_952) );
INVx1_ASAP7_75t_L g1051 ( .A(n_919), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1486 ( .A1(n_923), .A2(n_924), .B1(n_1481), .B2(n_1482), .Y(n_1486) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_924), .A2(n_972), .B1(n_984), .B2(n_985), .Y(n_983) );
INVx2_ASAP7_75t_L g1002 ( .A(n_925), .Y(n_1002) );
INVx2_ASAP7_75t_L g1250 ( .A(n_925), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
XOR2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_1175), .Y(n_944) );
XNOR2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_1072), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
XNOR2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_1009), .Y(n_947) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OR2x2_ASAP7_75t_L g951 ( .A(n_952), .B(n_980), .Y(n_951) );
AOI21xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_962), .B(n_963), .Y(n_953) );
INVx2_ASAP7_75t_SL g1636 ( .A(n_955), .Y(n_1636) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx4_ASAP7_75t_L g1192 ( .A(n_957), .Y(n_1192) );
INVx2_ASAP7_75t_L g1539 ( .A(n_957), .Y(n_1539) );
INVx4_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_969), .Y(n_963) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g1479 ( .A(n_966), .Y(n_1479) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_974), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_973) );
NAND3xp33_ASAP7_75t_SL g980 ( .A(n_981), .B(n_983), .C(n_986), .Y(n_980) );
NOR2xp33_ASAP7_75t_SL g986 ( .A(n_987), .B(n_991), .Y(n_986) );
BUFx6f_ASAP7_75t_L g1609 ( .A(n_990), .Y(n_1609) );
OAI33xp33_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_993), .A3(n_996), .B1(n_1001), .B2(n_1005), .B3(n_1008), .Y(n_991) );
BUFx3_ASAP7_75t_L g1551 ( .A(n_992), .Y(n_1551) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_998), .A2(n_1002), .B1(n_1003), .B2(n_1004), .Y(n_1001) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
BUFx2_ASAP7_75t_L g1044 ( .A(n_999), .Y(n_1044) );
NAND4xp75_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1052), .C(n_1064), .D(n_1069), .Y(n_1010) );
OAI21x1_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1028), .B(n_1050), .Y(n_1011) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1016), .B(n_1024), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_1014), .A2(n_1082), .B1(n_1112), .B2(n_1116), .Y(n_1111) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
AOI221xp5_ASAP7_75t_SL g1016 ( .A1(n_1017), .A2(n_1018), .B1(n_1019), .B2(n_1021), .C(n_1022), .Y(n_1016) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1020), .Y(n_1284) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1020), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1554 ( .A1(n_1023), .A2(n_1538), .B1(n_1548), .B2(n_1555), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1034), .B1(n_1039), .B2(n_1045), .Y(n_1028) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1041), .B1(n_1042), .B2(n_1043), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1929 ( .A1(n_1043), .A2(n_1047), .B1(n_1918), .B2(n_1924), .Y(n_1929) );
INVx3_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
AOI211x1_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1054), .B(n_1057), .C(n_1063), .Y(n_1052) );
INVx1_ASAP7_75t_L g1959 ( .A(n_1056), .Y(n_1959) );
OAI33xp33_ASAP7_75t_L g1911 ( .A1(n_1058), .A2(n_1912), .A3(n_1913), .B1(n_1917), .B2(n_1920), .B3(n_1923), .Y(n_1911) );
INVx6_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx5_ASAP7_75t_L g1164 ( .A(n_1061), .Y(n_1164) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVxp67_ASAP7_75t_L g1394 ( .A(n_1067), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1122), .B1(n_1123), .B2(n_1174), .Y(n_1072) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1073), .Y(n_1174) );
OAI21x1_ASAP7_75t_SL g1073 ( .A1(n_1074), .A2(n_1075), .B(n_1121), .Y(n_1073) );
NAND4xp25_ASAP7_75t_L g1121 ( .A(n_1074), .B(n_1077), .C(n_1079), .D(n_1098), .Y(n_1121) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
NAND3xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1079), .C(n_1098), .Y(n_1076) );
NOR2xp33_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1084), .Y(n_1079) );
NAND3xp33_ASAP7_75t_SL g1084 ( .A(n_1085), .B(n_1089), .C(n_1094), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g1089 ( .A1(n_1090), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g1152 ( .A1(n_1090), .A2(n_1092), .B1(n_1153), .B2(n_1154), .Y(n_1152) );
AOI222xp33_ASAP7_75t_L g1393 ( .A1(n_1090), .A2(n_1092), .B1(n_1367), .B2(n_1394), .C1(n_1395), .C2(n_1396), .Y(n_1393) );
NAND3xp33_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1105), .C(n_1111), .Y(n_1099) );
NOR2xp33_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1104), .Y(n_1100) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
NOR3xp33_ASAP7_75t_L g1216 ( .A(n_1104), .B(n_1217), .C(n_1221), .Y(n_1216) );
NOR3xp33_ASAP7_75t_L g1232 ( .A(n_1104), .B(n_1233), .C(n_1238), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .B1(n_1109), .B2(n_1110), .Y(n_1105) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
NOR2x1_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1148), .Y(n_1124) );
NOR3xp33_ASAP7_75t_SL g1130 ( .A(n_1131), .B(n_1139), .C(n_1140), .Y(n_1130) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g1931 ( .A1(n_1135), .A2(n_1385), .B1(n_1915), .B2(n_1922), .Y(n_1931) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_1137), .A2(n_1171), .B1(n_1172), .B2(n_1173), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_1138), .A2(n_1161), .B1(n_1163), .B2(n_1164), .Y(n_1160) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1156), .Y(n_1148) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_1161), .A2(n_1185), .B1(n_1186), .B2(n_1187), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_1161), .A2(n_1164), .B1(n_1407), .B2(n_1408), .Y(n_1406) );
OAI22xp5_ASAP7_75t_L g1923 ( .A1(n_1161), .A2(n_1164), .B1(n_1924), .B2(n_1925), .Y(n_1923) );
BUFx4f_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVxp67_ASAP7_75t_L g1201 ( .A(n_1162), .Y(n_1201) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1162), .Y(n_1535) );
OR2x6_ASAP7_75t_L g1576 ( .A(n_1162), .B(n_1577), .Y(n_1576) );
OR2x6_ASAP7_75t_L g1582 ( .A(n_1162), .B(n_1583), .Y(n_1582) );
OAI22xp33_ASAP7_75t_L g1530 ( .A1(n_1164), .A2(n_1531), .B1(n_1532), .B2(n_1536), .Y(n_1530) );
OAI33xp33_ASAP7_75t_L g1956 ( .A1(n_1166), .A2(n_1544), .A3(n_1957), .B1(n_1960), .B2(n_1963), .B3(n_1965), .Y(n_1956) );
OAI22xp33_ASAP7_75t_L g1913 ( .A1(n_1171), .A2(n_1914), .B1(n_1915), .B2(n_1916), .Y(n_1913) );
XNOR2xp5_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1270), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
XNOR2x1_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1227), .Y(n_1177) );
XNOR2x1_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
NOR2x1_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1212), .Y(n_1180) );
NAND3xp33_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1206), .C(n_1210), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1205), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_1187), .A2(n_1200), .B1(n_1202), .B2(n_1203), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1190), .B1(n_1192), .B2(n_1193), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1962 ( .A(n_1190), .Y(n_1962) );
INVx2_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1191), .Y(n_1327) );
INVx4_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
A2O1A1Ixp33_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1216), .B(n_1224), .C(n_1225), .Y(n_1212) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
AOI21xp5_ASAP7_75t_L g1292 ( .A1(n_1224), .A2(n_1293), .B(n_1312), .Y(n_1292) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
XNOR2x1_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1230), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1257), .Y(n_1230) );
A2O1A1Ixp33_ASAP7_75t_L g1231 ( .A1(n_1232), .A2(n_1247), .B(n_1255), .C(n_1256), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_1243), .A2(n_1244), .B1(n_1245), .B2(n_1246), .Y(n_1242) );
INVx2_ASAP7_75t_L g1614 ( .A(n_1243), .Y(n_1614) );
OAI22xp5_ASAP7_75t_L g1946 ( .A1(n_1245), .A2(n_1947), .B1(n_1948), .B2(n_1949), .Y(n_1946) );
HB1xp67_ASAP7_75t_L g1885 ( .A(n_1251), .Y(n_1885) );
A2O1A1Ixp33_ASAP7_75t_SL g1365 ( .A1(n_1255), .A2(n_1366), .B(n_1370), .C(n_1390), .Y(n_1365) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1266), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_1271), .A2(n_1314), .B1(n_1357), .B2(n_1358), .Y(n_1270) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1271), .Y(n_1358) );
NAND2xp67_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1292), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1285), .B1(n_1288), .B2(n_1291), .Y(n_1280) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
NAND3xp33_ASAP7_75t_SL g1293 ( .A(n_1294), .B(n_1297), .C(n_1302), .Y(n_1293) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
HB1xp67_ASAP7_75t_L g1405 ( .A(n_1308), .Y(n_1405) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1314), .Y(n_1357) );
XOR2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1356), .Y(n_1314) );
NOR2x1_ASAP7_75t_SL g1315 ( .A(n_1316), .B(n_1338), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1329), .Y(n_1319) );
OAI211xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1322), .B(n_1324), .C(n_1325), .Y(n_1320) );
OAI22xp5_ASAP7_75t_SL g1957 ( .A1(n_1322), .A2(n_1944), .B1(n_1954), .B2(n_1958), .Y(n_1957) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx2_ASAP7_75t_L g1627 ( .A(n_1323), .Y(n_1627) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
NOR3xp33_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1349), .C(n_1352), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1355), .Y(n_1353) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1359), .Y(n_1646) );
AOI22xp5_ASAP7_75t_SL g1359 ( .A1(n_1360), .A2(n_1447), .B1(n_1644), .B2(n_1645), .Y(n_1359) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1360), .Y(n_1644) );
OA22x2_ASAP7_75t_L g1360 ( .A1(n_1361), .A2(n_1362), .B1(n_1413), .B2(n_1414), .Y(n_1360) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
NOR3xp33_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1382), .C(n_1383), .Y(n_1370) );
NOR3xp33_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1375), .C(n_1381), .Y(n_1371) );
NOR2xp33_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1374), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1404 ( .A(n_1373), .B(n_1400), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1379), .Y(n_1375) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
OAI22xp33_ASAP7_75t_L g1552 ( .A1(n_1385), .A2(n_1531), .B1(n_1542), .B2(n_1553), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g1607 ( .A1(n_1385), .A2(n_1608), .B1(n_1609), .B2(n_1610), .Y(n_1607) );
OAI22xp33_ASAP7_75t_L g1927 ( .A1(n_1385), .A2(n_1914), .B1(n_1921), .B2(n_1928), .Y(n_1927) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
NAND3xp33_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1397), .C(n_1411), .Y(n_1392) );
AOI22xp5_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1403), .B1(n_1409), .B2(n_1410), .Y(n_1397) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_1399), .A2(n_1404), .B1(n_1405), .B2(n_1406), .Y(n_1403) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1432), .Y(n_1415) );
NAND3xp33_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1421), .C(n_1424), .Y(n_1417) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1447), .Y(n_1645) );
XOR2xp5_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1487), .Y(n_1447) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
HB1xp67_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1470), .Y(n_1451) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1468), .Y(n_1600) );
AOI21xp5_ASAP7_75t_L g1470 ( .A1(n_1471), .A2(n_1483), .B(n_1485), .Y(n_1470) );
NAND3xp33_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1475), .C(n_1480), .Y(n_1471) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
AOI22x1_ASAP7_75t_L g1487 ( .A1(n_1488), .A2(n_1489), .B1(n_1592), .B2(n_1642), .Y(n_1487) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1490), .Y(n_1590) );
OAI211xp5_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1497), .B(n_1526), .C(n_1559), .Y(n_1490) );
CKINVDCx14_ASAP7_75t_R g1491 ( .A(n_1492), .Y(n_1491) );
OAI31xp33_ASAP7_75t_L g1879 ( .A1(n_1492), .A2(n_1880), .A3(n_1884), .B(n_1890), .Y(n_1879) );
AND2x4_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1495), .Y(n_1492) );
AND2x2_ASAP7_75t_SL g1990 ( .A(n_1493), .B(n_1495), .Y(n_1990) );
INVx1_ASAP7_75t_SL g1493 ( .A(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
NOR3xp33_ASAP7_75t_SL g1497 ( .A(n_1498), .B(n_1505), .C(n_1520), .Y(n_1497) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx2_ASAP7_75t_SL g1500 ( .A(n_1501), .Y(n_1500) );
INVx2_ASAP7_75t_SL g1882 ( .A(n_1501), .Y(n_1882) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx2_ASAP7_75t_L g1883 ( .A(n_1503), .Y(n_1883) );
INVx2_ASAP7_75t_L g1980 ( .A(n_1503), .Y(n_1980) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
CKINVDCx8_ASAP7_75t_R g1508 ( .A(n_1509), .Y(n_1508) );
CKINVDCx8_ASAP7_75t_R g1886 ( .A(n_1509), .Y(n_1886) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_1511), .A2(n_1515), .B1(n_1516), .B2(n_1519), .Y(n_1510) );
AOI22xp33_ASAP7_75t_SL g1887 ( .A1(n_1511), .A2(n_1517), .B1(n_1888), .B2(n_1889), .Y(n_1887) );
BUFx3_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
BUFx3_ASAP7_75t_L g1983 ( .A(n_1512), .Y(n_1983) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1514), .Y(n_1512) );
AND2x4_ASAP7_75t_L g1517 ( .A(n_1513), .B(n_1518), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_1515), .A2(n_1566), .B1(n_1569), .B2(n_1570), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1982 ( .A1(n_1516), .A2(n_1969), .B1(n_1983), .B2(n_1984), .Y(n_1982) );
BUFx6f_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
BUFx2_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
BUFx3_ASAP7_75t_L g1891 ( .A(n_1522), .Y(n_1891) );
INVx2_ASAP7_75t_SL g1987 ( .A(n_1522), .Y(n_1987) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVx2_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1525), .Y(n_1893) );
BUFx3_ASAP7_75t_L g1988 ( .A(n_1525), .Y(n_1988) );
NOR2xp33_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1550), .Y(n_1526) );
OAI33xp33_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1530), .A3(n_1537), .B1(n_1541), .B2(n_1544), .B3(n_1546), .Y(n_1527) );
BUFx6f_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx2_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
OAI33xp33_ASAP7_75t_L g1550 ( .A1(n_1551), .A2(n_1552), .A3(n_1554), .B1(n_1556), .B2(n_1557), .B3(n_1558), .Y(n_1550) );
OAI31xp33_ASAP7_75t_L g1559 ( .A1(n_1560), .A2(n_1573), .A3(n_1581), .B(n_1586), .Y(n_1559) );
INVx3_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1897 ( .A(n_1563), .Y(n_1897) );
BUFx3_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
AOI22xp33_ASAP7_75t_L g1968 ( .A1(n_1567), .A2(n_1969), .B1(n_1970), .B2(n_1971), .Y(n_1968) );
INVx2_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx2_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx2_ASAP7_75t_L g1901 ( .A(n_1572), .Y(n_1901) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
BUFx2_ASAP7_75t_L g1904 ( .A(n_1576), .Y(n_1904) );
HB1xp67_ASAP7_75t_L g1973 ( .A(n_1576), .Y(n_1973) );
HB1xp67_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
BUFx2_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx2_ASAP7_75t_L g1906 ( .A(n_1580), .Y(n_1906) );
INVx3_ASAP7_75t_L g1660 ( .A(n_1582), .Y(n_1660) );
CKINVDCx16_ASAP7_75t_R g1584 ( .A(n_1585), .Y(n_1584) );
INVx4_ASAP7_75t_L g1908 ( .A(n_1585), .Y(n_1908) );
INVx3_ASAP7_75t_SL g1977 ( .A(n_1585), .Y(n_1977) );
OAI31xp33_ASAP7_75t_L g1966 ( .A1(n_1586), .A2(n_1967), .A3(n_1972), .B(n_1975), .Y(n_1966) );
BUFx3_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
BUFx2_ASAP7_75t_SL g1909 ( .A(n_1587), .Y(n_1909) );
AND2x4_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1589), .Y(n_1587) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1588), .Y(n_1659) );
NOR2xp33_ASAP7_75t_L g1934 ( .A(n_1588), .B(n_1651), .Y(n_1934) );
INVxp67_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AND3x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1620), .C(n_1623), .Y(n_1595) );
AOI211xp5_ASAP7_75t_SL g1596 ( .A1(n_1597), .A2(n_1598), .B(n_1599), .C(n_1602), .Y(n_1596) );
OAI221xp5_ASAP7_75t_L g1634 ( .A1(n_1608), .A2(n_1626), .B1(n_1635), .B2(n_1637), .C(n_1638), .Y(n_1634) );
INVx2_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
OAI33xp33_ASAP7_75t_L g1941 ( .A1(n_1618), .A2(n_1942), .A3(n_1943), .B1(n_1946), .B2(n_1950), .B3(n_1953), .Y(n_1941) );
OAI22xp5_ASAP7_75t_L g1965 ( .A1(n_1626), .A2(n_1949), .B1(n_1952), .B2(n_1958), .Y(n_1965) );
INVx2_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
INVxp67_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
INVx2_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
BUFx3_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
INVx3_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1657), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
NOR2xp33_ASAP7_75t_L g1652 ( .A(n_1653), .B(n_1655), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1993 ( .A(n_1653), .B(n_1656), .Y(n_1993) );
INVx1_ASAP7_75t_L g1995 ( .A(n_1653), .Y(n_1995) );
HB1xp67_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
NOR2xp33_ASAP7_75t_L g1997 ( .A(n_1656), .B(n_1995), .Y(n_1997) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1660), .Y(n_1658) );
AND2x4_ASAP7_75t_SL g1933 ( .A(n_1660), .B(n_1934), .Y(n_1933) );
INVx1_ASAP7_75t_L g1976 ( .A(n_1660), .Y(n_1976) );
OAI221xp5_ASAP7_75t_L g1661 ( .A1(n_1662), .A2(n_1875), .B1(n_1877), .B2(n_1932), .C(n_1935), .Y(n_1661) );
AOI21xp5_ASAP7_75t_L g1662 ( .A1(n_1663), .A2(n_1786), .B(n_1845), .Y(n_1662) );
NAND5xp2_ASAP7_75t_L g1663 ( .A(n_1664), .B(n_1729), .C(n_1749), .D(n_1762), .E(n_1772), .Y(n_1663) );
O2A1O1Ixp33_ASAP7_75t_L g1664 ( .A1(n_1665), .A2(n_1696), .B(n_1703), .C(n_1714), .Y(n_1664) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1665), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1666), .B(n_1686), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1666), .B(n_1693), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1666), .B(n_1688), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1666), .B(n_1687), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1798 ( .A(n_1666), .B(n_1799), .Y(n_1798) );
NAND2xp5_ASAP7_75t_L g1834 ( .A(n_1666), .B(n_1700), .Y(n_1834) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1666), .Y(n_1857) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1667), .B(n_1682), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1667), .B(n_1728), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1667), .B(n_1687), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1667), .B(n_1683), .Y(n_1748) );
AND3x1_ASAP7_75t_L g1822 ( .A(n_1667), .B(n_1683), .C(n_1687), .Y(n_1822) );
OR2x2_ASAP7_75t_L g1863 ( .A(n_1667), .B(n_1728), .Y(n_1863) );
INVx2_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1668), .B(n_1682), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1753 ( .A(n_1668), .B(n_1683), .Y(n_1753) );
OR2x2_ASAP7_75t_L g1668 ( .A(n_1669), .B(n_1676), .Y(n_1668) );
INVx2_ASAP7_75t_L g1783 ( .A(n_1670), .Y(n_1783) );
AND2x6_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1672), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1671), .B(n_1675), .Y(n_1674) );
AND2x4_ASAP7_75t_L g1677 ( .A(n_1671), .B(n_1678), .Y(n_1677) );
AND2x6_ASAP7_75t_L g1680 ( .A(n_1671), .B(n_1681), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1671), .B(n_1675), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1671), .B(n_1675), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1673), .B(n_1679), .Y(n_1678) );
INVxp67_ASAP7_75t_L g1785 ( .A(n_1674), .Y(n_1785) );
HB1xp67_ASAP7_75t_L g1876 ( .A(n_1674), .Y(n_1876) );
OAI21xp5_ASAP7_75t_L g1994 ( .A1(n_1675), .A2(n_1995), .B(n_1996), .Y(n_1994) );
AND2x2_ASAP7_75t_L g1825 ( .A(n_1682), .B(n_1728), .Y(n_1825) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
OR2x2_ASAP7_75t_L g1758 ( .A(n_1683), .B(n_1728), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1819 ( .A(n_1683), .B(n_1728), .Y(n_1819) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1685), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1686), .B(n_1748), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1833 ( .A(n_1686), .B(n_1753), .Y(n_1833) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1686), .Y(n_1860) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1692), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1768 ( .A(n_1687), .B(n_1702), .Y(n_1768) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1687), .B(n_1771), .Y(n_1770) );
INVx2_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1688), .B(n_1702), .Y(n_1701) );
OAI322xp33_ASAP7_75t_L g1714 ( .A1(n_1688), .A2(n_1710), .A3(n_1715), .B1(n_1721), .B2(n_1723), .C1(n_1725), .C2(n_1726), .Y(n_1714) );
BUFx2_ASAP7_75t_L g1728 ( .A(n_1688), .Y(n_1728) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1688), .B(n_1752), .Y(n_1751) );
AOI321xp33_ASAP7_75t_L g1772 ( .A1(n_1688), .A2(n_1773), .A3(n_1774), .B1(n_1775), .B2(n_1777), .C(n_1779), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1810 ( .A(n_1688), .B(n_1753), .Y(n_1810) );
OR2x2_ASAP7_75t_L g1871 ( .A(n_1688), .B(n_1805), .Y(n_1871) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1692), .B(n_1704), .Y(n_1767) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_1692), .B(n_1753), .Y(n_1771) );
NOR2xp33_ASAP7_75t_L g1777 ( .A(n_1692), .B(n_1778), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1820 ( .A(n_1692), .B(n_1744), .Y(n_1820) );
NAND2xp5_ASAP7_75t_L g1844 ( .A(n_1692), .B(n_1702), .Y(n_1844) );
OAI21xp33_ASAP7_75t_L g1865 ( .A1(n_1692), .A2(n_1844), .B(n_1866), .Y(n_1865) );
INVx2_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1693), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1693), .B(n_1706), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1693), .B(n_1710), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1797 ( .A(n_1693), .B(n_1728), .Y(n_1797) );
NAND2xp5_ASAP7_75t_L g1805 ( .A(n_1693), .B(n_1753), .Y(n_1805) );
NAND2xp5_ASAP7_75t_L g1853 ( .A(n_1693), .B(n_1718), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1695), .Y(n_1693) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1701), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1827 ( .A(n_1698), .B(n_1763), .Y(n_1827) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1699), .B(n_1716), .Y(n_1715) );
NOR2xp33_ASAP7_75t_L g1757 ( .A(n_1699), .B(n_1758), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1699), .B(n_1790), .Y(n_1789) );
AND2x2_ASAP7_75t_L g1821 ( .A(n_1699), .B(n_1822), .Y(n_1821) );
AND2x2_ASAP7_75t_L g1829 ( .A(n_1699), .B(n_1768), .Y(n_1829) );
INVx2_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1799 ( .A(n_1700), .B(n_1716), .Y(n_1799) );
O2A1O1Ixp33_ASAP7_75t_L g1873 ( .A1(n_1700), .A2(n_1842), .B(n_1843), .C(n_1874), .Y(n_1873) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1701), .Y(n_1874) );
OR2x2_ASAP7_75t_L g1773 ( .A(n_1702), .B(n_1748), .Y(n_1773) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1702), .Y(n_1843) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1709), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1776 ( .A(n_1704), .B(n_1710), .Y(n_1776) );
INVx2_ASAP7_75t_L g1794 ( .A(n_1704), .Y(n_1794) );
A2O1A1O1Ixp25_ASAP7_75t_L g1839 ( .A1(n_1704), .A2(n_1718), .B(n_1796), .C(n_1840), .D(n_1841), .Y(n_1839) );
OR2x2_ASAP7_75t_L g1854 ( .A(n_1704), .B(n_1855), .Y(n_1854) );
INVx2_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1705), .B(n_1709), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1705), .B(n_1718), .Y(n_1732) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1706), .B(n_1718), .Y(n_1717) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1706), .B(n_1745), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1832 ( .A(n_1706), .B(n_1718), .Y(n_1832) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1708), .Y(n_1706) );
NAND2xp5_ASAP7_75t_L g1725 ( .A(n_1709), .B(n_1716), .Y(n_1725) );
NOR2xp33_ASAP7_75t_L g1756 ( .A(n_1709), .B(n_1717), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_1709), .B(n_1744), .Y(n_1791) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1709), .B(n_1718), .Y(n_1801) );
OR2x2_ASAP7_75t_L g1812 ( .A(n_1709), .B(n_1718), .Y(n_1812) );
CKINVDCx6p67_ASAP7_75t_R g1709 ( .A(n_1710), .Y(n_1709) );
OR2x2_ASAP7_75t_L g1755 ( .A(n_1710), .B(n_1718), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1710), .B(n_1718), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1836 ( .A(n_1710), .B(n_1837), .Y(n_1836) );
CKINVDCx5p33_ASAP7_75t_R g1858 ( .A(n_1710), .Y(n_1858) );
OR2x2_ASAP7_75t_L g1861 ( .A(n_1710), .B(n_1731), .Y(n_1861) );
OR2x6_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1713), .Y(n_1710) );
OR2x2_ASAP7_75t_L g1814 ( .A(n_1711), .B(n_1713), .Y(n_1814) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1715), .Y(n_1847) );
NAND2xp5_ASAP7_75t_L g1741 ( .A(n_1716), .B(n_1722), .Y(n_1741) );
INVx2_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
INVx3_ASAP7_75t_L g1736 ( .A(n_1718), .Y(n_1736) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1718), .Y(n_1745) );
AOI22xp5_ASAP7_75t_L g1762 ( .A1(n_1718), .A2(n_1763), .B1(n_1764), .B2(n_1769), .Y(n_1762) );
AND2x4_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1720), .Y(n_1718) );
INVxp67_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1724), .B(n_1761), .Y(n_1760) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1725), .Y(n_1872) );
CKINVDCx14_ASAP7_75t_R g1726 ( .A(n_1727), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1802 ( .A(n_1728), .B(n_1748), .Y(n_1802) );
NOR2xp33_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1742), .Y(n_1729) );
OAI211xp5_ASAP7_75t_L g1730 ( .A1(n_1731), .A2(n_1733), .B(n_1734), .C(n_1741), .Y(n_1730) );
AOI21xp33_ASAP7_75t_L g1803 ( .A1(n_1731), .A2(n_1804), .B(n_1805), .Y(n_1803) );
CKINVDCx6p67_ASAP7_75t_R g1731 ( .A(n_1732), .Y(n_1731) );
AOI21xp33_ASAP7_75t_L g1867 ( .A1(n_1733), .A2(n_1808), .B(n_1868), .Y(n_1867) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1735), .B(n_1737), .Y(n_1734) );
CKINVDCx14_ASAP7_75t_R g1735 ( .A(n_1736), .Y(n_1735) );
AOI221xp5_ASAP7_75t_L g1869 ( .A1(n_1737), .A2(n_1763), .B1(n_1870), .B2(n_1872), .C(n_1873), .Y(n_1869) );
NOR2xp33_ASAP7_75t_L g1737 ( .A(n_1738), .B(n_1740), .Y(n_1737) );
CKINVDCx14_ASAP7_75t_R g1738 ( .A(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1740), .Y(n_1837) );
NOR2xp33_ASAP7_75t_L g1742 ( .A(n_1743), .B(n_1746), .Y(n_1742) );
AOI21xp5_ASAP7_75t_L g1848 ( .A1(n_1743), .A2(n_1849), .B(n_1850), .Y(n_1848) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1748), .Y(n_1778) );
AOI221xp5_ASAP7_75t_L g1749 ( .A1(n_1750), .A2(n_1754), .B1(n_1756), .B2(n_1757), .C(n_1759), .Y(n_1749) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_1751), .B(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1753), .B(n_1797), .Y(n_1796) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1755), .B(n_1761), .Y(n_1804) );
OAI221xp5_ASAP7_75t_L g1841 ( .A1(n_1755), .A2(n_1779), .B1(n_1842), .B2(n_1843), .C(n_1844), .Y(n_1841) );
AOI221xp5_ASAP7_75t_L g1851 ( .A1(n_1756), .A2(n_1790), .B1(n_1852), .B2(n_1858), .C(n_1859), .Y(n_1851) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
AOI222xp33_ASAP7_75t_L g1815 ( .A1(n_1763), .A2(n_1816), .B1(n_1820), .B2(n_1821), .C1(n_1823), .C2(n_1826), .Y(n_1815) );
NAND2xp5_ASAP7_75t_L g1842 ( .A(n_1763), .B(n_1794), .Y(n_1842) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
NOR2xp33_ASAP7_75t_L g1813 ( .A(n_1765), .B(n_1814), .Y(n_1813) );
NAND2xp5_ASAP7_75t_L g1765 ( .A(n_1766), .B(n_1768), .Y(n_1765) );
OAI21xp33_ASAP7_75t_L g1800 ( .A1(n_1766), .A2(n_1801), .B(n_1802), .Y(n_1800) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1768), .Y(n_1817) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
AOI211xp5_ASAP7_75t_SL g1859 ( .A1(n_1771), .A2(n_1860), .B(n_1861), .C(n_1862), .Y(n_1859) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
OAI22xp5_ASAP7_75t_L g1830 ( .A1(n_1776), .A2(n_1831), .B1(n_1833), .B2(n_1834), .Y(n_1830) );
INVx2_ASAP7_75t_SL g1779 ( .A(n_1780), .Y(n_1779) );
OAI22xp5_ASAP7_75t_SL g1781 ( .A1(n_1782), .A2(n_1783), .B1(n_1784), .B2(n_1785), .Y(n_1781) );
NAND5xp2_ASAP7_75t_L g1786 ( .A(n_1787), .B(n_1806), .C(n_1815), .D(n_1828), .E(n_1839), .Y(n_1786) );
AOI211xp5_ASAP7_75t_L g1787 ( .A1(n_1788), .A2(n_1791), .B(n_1792), .C(n_1803), .Y(n_1787) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
AOI221xp5_ASAP7_75t_L g1864 ( .A1(n_1791), .A2(n_1821), .B1(n_1832), .B2(n_1865), .C(n_1867), .Y(n_1864) );
OAI211xp5_ASAP7_75t_L g1792 ( .A1(n_1793), .A2(n_1795), .B(n_1798), .C(n_1800), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1793), .B(n_1809), .Y(n_1808) );
INVx2_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1797), .Y(n_1856) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1799), .Y(n_1838) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1801), .Y(n_1868) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1802), .Y(n_1866) );
INVxp67_ASAP7_75t_SL g1840 ( .A(n_1804), .Y(n_1840) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1805), .Y(n_1809) );
O2A1O1Ixp33_ASAP7_75t_SL g1806 ( .A1(n_1807), .A2(n_1810), .B(n_1811), .C(n_1813), .Y(n_1806) );
INVxp67_ASAP7_75t_SL g1807 ( .A(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1810), .Y(n_1850) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
AOI211xp5_ASAP7_75t_L g1828 ( .A1(n_1814), .A2(n_1829), .B(n_1830), .C(n_1835), .Y(n_1828) );
A2O1A1Ixp33_ASAP7_75t_L g1846 ( .A1(n_1814), .A2(n_1819), .B(n_1847), .C(n_1848), .Y(n_1846) );
NAND2xp5_ASAP7_75t_SL g1816 ( .A(n_1817), .B(n_1818), .Y(n_1816) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
AOI21xp33_ASAP7_75t_L g1835 ( .A1(n_1824), .A2(n_1836), .B(n_1838), .Y(n_1835) );
OAI21xp33_ASAP7_75t_L g1852 ( .A1(n_1824), .A2(n_1853), .B(n_1854), .Y(n_1852) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVxp67_ASAP7_75t_SL g1826 ( .A(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1849 ( .A(n_1829), .Y(n_1849) );
INVx2_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
NAND4xp25_ASAP7_75t_L g1845 ( .A(n_1846), .B(n_1851), .C(n_1864), .D(n_1869), .Y(n_1845) );
OR2x2_ASAP7_75t_L g1855 ( .A(n_1856), .B(n_1857), .Y(n_1855) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1863), .Y(n_1862) );
INVx1_ASAP7_75t_L g1870 ( .A(n_1871), .Y(n_1870) );
INVx4_ASAP7_75t_L g1875 ( .A(n_1876), .Y(n_1875) );
NAND3xp33_ASAP7_75t_L g1878 ( .A(n_1879), .B(n_1894), .C(n_1910), .Y(n_1878) );
INVx2_ASAP7_75t_SL g1881 ( .A(n_1882), .Y(n_1881) );
AOI22xp33_ASAP7_75t_L g1898 ( .A1(n_1888), .A2(n_1899), .B1(n_1900), .B2(n_1902), .Y(n_1898) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1893), .Y(n_1892) );
OAI31xp33_ASAP7_75t_L g1894 ( .A1(n_1895), .A2(n_1903), .A3(n_1907), .B(n_1909), .Y(n_1894) );
INVx2_ASAP7_75t_L g1900 ( .A(n_1901), .Y(n_1900) );
INVx2_ASAP7_75t_L g1971 ( .A(n_1901), .Y(n_1971) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1906), .Y(n_1905) );
INVx2_ASAP7_75t_L g1974 ( .A(n_1906), .Y(n_1974) );
NOR2xp33_ASAP7_75t_L g1910 ( .A(n_1911), .B(n_1926), .Y(n_1910) );
INVx3_ASAP7_75t_L g1932 ( .A(n_1933), .Y(n_1932) );
INVxp33_ASAP7_75t_L g1936 ( .A(n_1937), .Y(n_1936) );
HB1xp67_ASAP7_75t_L g1938 ( .A(n_1939), .Y(n_1938) );
NAND3xp33_ASAP7_75t_L g1939 ( .A(n_1940), .B(n_1966), .C(n_1978), .Y(n_1939) );
NOR2xp33_ASAP7_75t_L g1940 ( .A(n_1941), .B(n_1956), .Y(n_1940) );
OAI22xp5_ASAP7_75t_L g1960 ( .A1(n_1947), .A2(n_1951), .B1(n_1961), .B2(n_1962), .Y(n_1960) );
INVx2_ASAP7_75t_L g1958 ( .A(n_1959), .Y(n_1958) );
OAI31xp33_ASAP7_75t_L g1978 ( .A1(n_1979), .A2(n_1981), .A3(n_1985), .B(n_1989), .Y(n_1978) );
INVx1_ASAP7_75t_L g1986 ( .A(n_1987), .Y(n_1986) );
BUFx2_ASAP7_75t_L g1989 ( .A(n_1990), .Y(n_1989) );
HB1xp67_ASAP7_75t_L g1991 ( .A(n_1992), .Y(n_1991) );
BUFx3_ASAP7_75t_L g1992 ( .A(n_1993), .Y(n_1992) );
INVx1_ASAP7_75t_L g1996 ( .A(n_1997), .Y(n_1996) );
endmodule