module real_jpeg_14193_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_0),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_0),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_10),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_12),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_2),
.B(n_12),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_8),
.B(n_13),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

NOR5xp2_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_16),
.C(n_28),
.D(n_38),
.E(n_41),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_17),
.B1(n_24),
.B2(n_26),
.Y(n_16)
);

OR2x2_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_11),
.B(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_15),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_25),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_23),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_30),
.B(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);


endmodule