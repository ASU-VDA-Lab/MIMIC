module fake_jpeg_29778_n_219 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_53),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_20),
.B1(n_18),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_77),
.B1(n_20),
.B2(n_17),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_38),
.B(n_27),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_46),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_31),
.B1(n_24),
.B2(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_56),
.B1(n_43),
.B2(n_22),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_94),
.B1(n_98),
.B2(n_55),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_52),
.B1(n_54),
.B2(n_50),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_88),
.B1(n_100),
.B2(n_67),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_91),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_75),
.B1(n_68),
.B2(n_69),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_42),
.B1(n_28),
.B2(n_25),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_102),
.B1(n_101),
.B2(n_97),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_78),
.B1(n_71),
.B2(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_25),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_101),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_28),
.B1(n_22),
.B2(n_34),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_99),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_55),
.B1(n_38),
.B2(n_29),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_21),
.B1(n_23),
.B2(n_31),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_74),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_110),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_66),
.C(n_72),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_114),
.C(n_100),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_92),
.B(n_87),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_92),
.B(n_85),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_21),
.C(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_78),
.B1(n_67),
.B2(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_86),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_125),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_100),
.B(n_88),
.C(n_86),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_127),
.B(n_115),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_128),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_88),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_82),
.C(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_133),
.B1(n_113),
.B2(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_107),
.A3(n_113),
.B1(n_115),
.B2(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_150),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_117),
.C(n_62),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_121),
.B1(n_136),
.B2(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_110),
.B1(n_95),
.B2(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_109),
.B1(n_118),
.B2(n_106),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_126),
.C(n_128),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_160),
.C(n_164),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_130),
.B(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_165),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_136),
.C(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_166),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_135),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_151),
.B1(n_145),
.B2(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_155),
.B1(n_106),
.B2(n_103),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_139),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_146),
.C(n_138),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_165),
.C(n_161),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_147),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_155),
.B1(n_158),
.B2(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_24),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_81),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.C(n_173),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_74),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_170),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_186),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_176),
.B1(n_174),
.B2(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_193),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_62),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_199),
.Y(n_202)
);

NAND4xp25_ASAP7_75t_SL g200 ( 
.A(n_188),
.B(n_16),
.C(n_15),
.D(n_14),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_180),
.B(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_179),
.B1(n_192),
.B2(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_204),
.B(n_205),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_190),
.B1(n_62),
.B2(n_16),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_14),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_10),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_11),
.B(n_1),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_209),
.B(n_2),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_2),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_204),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_212),
.A2(n_213),
.B(n_5),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_5),
.B(n_7),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_214),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_9),
.B(n_10),
.Y(n_219)
);


endmodule