module fake_jpeg_20502_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_0),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_6),
.A2(n_5),
.B1(n_0),
.B2(n_1),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_19),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_8),
.B1(n_16),
.B2(n_19),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_10),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_12),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_15),
.C(n_11),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_11),
.B1(n_8),
.B2(n_13),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_32),
.B1(n_34),
.B2(n_28),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_33),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_25),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_30),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_44),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.C(n_40),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_47),
.C(n_43),
.Y(n_49)
);


endmodule