module fake_jpeg_20004_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_62),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_33),
.B(n_28),
.C(n_35),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_59),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_28),
.B1(n_33),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_68),
.B1(n_77),
.B2(n_31),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_21),
.B1(n_34),
.B2(n_19),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_21),
.B1(n_34),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_29),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_17),
.B1(n_36),
.B2(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_26),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_0),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_35),
.B1(n_29),
.B2(n_30),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_65),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_40),
.B1(n_20),
.B2(n_36),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_94),
.B1(n_99),
.B2(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_20),
.B1(n_32),
.B2(n_17),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_105),
.B1(n_106),
.B2(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_120),
.B1(n_76),
.B2(n_60),
.Y(n_138)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_37),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_109),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_37),
.B1(n_26),
.B2(n_9),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_61),
.A2(n_37),
.B1(n_26),
.B2(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_0),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_112),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_1),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_81),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_2),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_2),
.Y(n_125)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_53),
.B1(n_75),
.B2(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_121),
.B(n_123),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_124),
.B(n_128),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g169 ( 
.A1(n_125),
.A2(n_138),
.B(n_151),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_80),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_72),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_136),
.C(n_140),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_146),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_58),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_13),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_79),
.B1(n_53),
.B2(n_76),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_151),
.B1(n_98),
.B2(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_153),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_109),
.B(n_11),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_10),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_108),
.B(n_95),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_103),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_71),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_94),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_92),
.A2(n_65),
.B1(n_64),
.B2(n_58),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_90),
.A2(n_64),
.B1(n_10),
.B2(n_5),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_112),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_169),
.B(n_134),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_172),
.B1(n_177),
.B2(n_178),
.Y(n_214)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_146),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_126),
.A2(n_138),
.B1(n_129),
.B2(n_131),
.Y(n_172)
);

NAND2x1p5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_129),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_215)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_126),
.A2(n_102),
.B1(n_108),
.B2(n_101),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_87),
.B1(n_117),
.B2(n_110),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_115),
.B1(n_111),
.B2(n_87),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_132),
.B1(n_135),
.B2(n_139),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_111),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_188),
.Y(n_199)
);

INVx2_ASAP7_75t_R g185 ( 
.A(n_125),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_8),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_152),
.Y(n_186)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_201),
.B1(n_168),
.B2(n_172),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_210),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_160),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_134),
.B(n_140),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_198),
.B(n_200),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_134),
.B(n_135),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_137),
.B1(n_152),
.B2(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_122),
.B(n_153),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_97),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_215),
.Y(n_221)
);

XOR2x2_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_180),
.Y(n_220)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_97),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_176),
.B(n_7),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_212),
.B(n_15),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_3),
.B(n_4),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_217),
.B1(n_191),
.B2(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_234),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_177),
.B1(n_164),
.B2(n_163),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_190),
.B1(n_214),
.B2(n_201),
.Y(n_250)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_167),
.A3(n_156),
.B1(n_162),
.B2(n_182),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_226),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_165),
.C(n_156),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_240),
.C(n_227),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_199),
.B(n_187),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_238),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_178),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_205),
.B(n_216),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_165),
.C(n_179),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_196),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_229),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_252),
.B(n_254),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_259),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_239),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_221),
.B1(n_231),
.B2(n_230),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_197),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_197),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_192),
.C(n_195),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_257),
.C(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_193),
.C(n_203),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_222),
.B1(n_232),
.B2(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_203),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_223),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_208),
.C(n_166),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_219),
.B1(n_230),
.B2(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_270),
.Y(n_282)
);

HB1xp67_ASAP7_75t_SL g267 ( 
.A(n_244),
.Y(n_267)
);

AOI31xp33_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_269),
.A3(n_262),
.B(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_277),
.B1(n_278),
.B2(n_249),
.Y(n_279)
);

AND2x4_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_243),
.B(n_228),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_259),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_250),
.A2(n_236),
.B1(n_220),
.B2(n_237),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_280),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_287),
.C(n_264),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_246),
.B1(n_237),
.B2(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_257),
.C(n_255),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_260),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_273),
.CI(n_274),
.CON(n_296),
.SN(n_296)
);

OAI322xp33_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_283),
.A3(n_284),
.B1(n_207),
.B2(n_286),
.C1(n_215),
.C2(n_282),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_291),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_277),
.B1(n_269),
.B2(n_276),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_297),
.B1(n_291),
.B2(n_288),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_281),
.C(n_280),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_202),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_274),
.B1(n_268),
.B2(n_208),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_207),
.C(n_287),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_210),
.B(n_215),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_158),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_305),
.B1(n_296),
.B2(n_293),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_303),
.A3(n_308),
.B1(n_300),
.B2(n_292),
.C1(n_294),
.C2(n_296),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_306),
.B(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_158),
.C(n_202),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_202),
.B(n_11),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_310),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_293),
.B(n_294),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_313),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_186),
.B(n_7),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_12),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

OAI311xp33_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_186),
.A3(n_12),
.B1(n_13),
.C1(n_4),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_315),
.C(n_318),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_3),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_4),
.Y(n_322)
);


endmodule