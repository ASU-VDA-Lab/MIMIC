module fake_jpeg_9435_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

HAxp5_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_22),
.CON(n_24),
.SN(n_24)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_20),
.A2(n_17),
.B1(n_13),
.B2(n_12),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_23),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_1),
.B(n_3),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_13),
.B1(n_16),
.B2(n_14),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_29),
.B1(n_13),
.B2(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_21),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_14),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_11),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_33),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_38),
.C(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_31),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_28),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_27),
.B1(n_34),
.B2(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_39),
.B1(n_30),
.B2(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_47),
.C(n_45),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_48),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_63),
.C(n_64),
.Y(n_66)
);

AOI321xp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_53),
.A3(n_9),
.B1(n_17),
.B2(n_29),
.C(n_12),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_60),
.B1(n_61),
.B2(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_6),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_71),
.B1(n_6),
.B2(n_8),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_1),
.B(n_3),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_74),
.B(n_3),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);


endmodule