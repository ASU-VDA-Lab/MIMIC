module fake_jpeg_5523_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_4),
.B(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_51)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_31),
.B1(n_29),
.B2(n_23),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_57),
.B1(n_58),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_49),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_16),
.C(n_20),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_55),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_53),
.B(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_23),
.B1(n_25),
.B2(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_28),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_71),
.Y(n_92)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_63),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_38),
.Y(n_78)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_87),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_69),
.B1(n_19),
.B2(n_73),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_50),
.B1(n_56),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_105),
.B1(n_79),
.B2(n_97),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_36),
.B1(n_42),
.B2(n_52),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_103),
.Y(n_128)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_36),
.B1(n_42),
.B2(n_32),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_63),
.B1(n_42),
.B2(n_36),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_15),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_15),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_39),
.B1(n_61),
.B2(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_70),
.C(n_69),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_125),
.C(n_126),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_84),
.B1(n_39),
.B2(n_60),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_129),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_81),
.C(n_75),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_76),
.C(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_15),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_84),
.B1(n_68),
.B2(n_64),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_92),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_89),
.B1(n_102),
.B2(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_2),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_144),
.B(n_150),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_99),
.C(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_125),
.C(n_111),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_88),
.B(n_87),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_140),
.B(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_148),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_86),
.B(n_107),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_84),
.B1(n_93),
.B2(n_95),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_110),
.B1(n_112),
.B2(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_149),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_104),
.B(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_159),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_110),
.B1(n_124),
.B2(n_130),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_169),
.B1(n_143),
.B2(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_114),
.C(n_115),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_112),
.B(n_129),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_146),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_132),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_160),
.C(n_150),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_175),
.Y(n_187)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_181),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_143),
.B1(n_135),
.B2(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_136),
.B1(n_142),
.B2(n_164),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_189),
.B(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_155),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_192),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_158),
.B(n_138),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_168),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_183),
.B(n_170),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_202),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_187),
.B(n_149),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_181),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_14),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_205),
.B(n_14),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_170),
.C(n_179),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_194),
.A3(n_157),
.B1(n_201),
.B2(n_189),
.C1(n_205),
.C2(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_3),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_172),
.C(n_190),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_208),
.B(n_210),
.C(n_3),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_11),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_199),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_3),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_6),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_214),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_224),
.B(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_7),
.C(n_9),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_222),
.B1(n_7),
.B2(n_11),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);


endmodule