module fake_jpeg_14665_n_217 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_24),
.B1(n_27),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_59),
.B1(n_63),
.B2(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_27),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_38),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_18),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_23),
.B1(n_0),
.B2(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_63),
.B1(n_26),
.B2(n_29),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_22),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_26),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_38),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_88),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_103),
.B1(n_71),
.B2(n_84),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_43),
.B1(n_56),
.B2(n_35),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_41),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_64),
.C(n_70),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_41),
.B1(n_53),
.B2(n_51),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_53),
.B1(n_62),
.B2(n_47),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_47),
.B1(n_44),
.B2(n_61),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_66),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_88),
.B1(n_104),
.B2(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_15),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_105),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_47),
.B1(n_101),
.B2(n_57),
.Y(n_137)
);

OAI221xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_125),
.B1(n_106),
.B2(n_118),
.C(n_84),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_117),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_81),
.B(n_80),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_111),
.B1(n_115),
.B2(n_50),
.C(n_25),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_78),
.B1(n_76),
.B2(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_85),
.B1(n_99),
.B2(n_91),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_74),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_126),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_85),
.C(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_67),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_94),
.B(n_92),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_141),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_113),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_140),
.C(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

OA21x2_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_108),
.B(n_110),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_42),
.C(n_34),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_57),
.B(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_25),
.B1(n_19),
.B2(n_17),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_25),
.B1(n_28),
.B2(n_19),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_19),
.B(n_17),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_116),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_148),
.C(n_151),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_158),
.B(n_160),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_115),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_114),
.C(n_124),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_114),
.C(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_119),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_132),
.B1(n_128),
.B2(n_144),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_1),
.B(n_3),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_42),
.C(n_34),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_1),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_17),
.C(n_28),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_133),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_171),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_164),
.B(n_173),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

AO221x1_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_132),
.B1(n_128),
.B2(n_141),
.C(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_175),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_153),
.B(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_181),
.B1(n_28),
.B2(n_5),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_147),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_187),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_166),
.B(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_3),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_7),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_172),
.B1(n_168),
.B2(n_165),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_191),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_172),
.C(n_165),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_195),
.C(n_9),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_7),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_186),
.A3(n_181),
.B1(n_180),
.B2(n_11),
.C1(n_12),
.C2(n_8),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_10),
.C(n_11),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_10),
.C(n_11),
.Y(n_203)
);

AOI31xp67_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_10),
.A3(n_13),
.B(n_14),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_194),
.B(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_13),
.B(n_14),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_13),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_213),
.B(n_28),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_207),
.B(n_28),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_215),
.Y(n_217)
);


endmodule