module fake_jpeg_19013_n_155 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_71),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_63),
.B1(n_70),
.B2(n_69),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_66),
.B1(n_65),
.B2(n_64),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_61),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_48),
.B1(n_73),
.B2(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_89),
.B1(n_82),
.B2(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_101),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_50),
.C(n_52),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_59),
.C(n_55),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_73),
.B1(n_54),
.B2(n_57),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_89),
.B1(n_66),
.B2(n_65),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_60),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_0),
.CI(n_1),
.CON(n_103),
.SN(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_1),
.Y(n_105)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_119),
.B(n_116),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_109),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_64),
.B1(n_68),
.B2(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_113),
.B1(n_106),
.B2(n_118),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_130),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_51),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_126),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_3),
.B(n_4),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_24),
.B(n_27),
.Y(n_139)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_23),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_134),
.B(n_136),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_7),
.B1(n_11),
.B2(n_14),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_138),
.B(n_139),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_120),
.B(n_128),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_132),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_123),
.B(n_136),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_121),
.B(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_28),
.B(n_30),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_31),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_38),
.B(n_39),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_41),
.B(n_43),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_44),
.Y(n_155)
);


endmodule