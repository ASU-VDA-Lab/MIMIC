module fake_jpeg_350_n_433 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_433);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_5),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_56),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_26),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_5),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_59),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_64),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_69),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_83),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_79),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_82),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_1),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_91),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

BUFx12f_ASAP7_75t_SL g93 ( 
.A(n_34),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_15),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_95),
.Y(n_138)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_36),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_115),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_15),
.B1(n_39),
.B2(n_32),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_134),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_70),
.B(n_83),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_40),
.B1(n_20),
.B2(n_19),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_121),
.B1(n_140),
.B2(n_61),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_20),
.B1(n_40),
.B2(n_42),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_42),
.B1(n_36),
.B2(n_14),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_86),
.B1(n_78),
.B2(n_73),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_53),
.A2(n_34),
.B1(n_36),
.B2(n_14),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_11),
.B(n_12),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_46),
.B(n_58),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_52),
.B(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_136),
.B(n_4),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_14),
.B1(n_36),
.B2(n_34),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_49),
.B(n_14),
.C(n_36),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_65),
.C(n_51),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_28),
.B(n_21),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_47),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_76),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_44),
.A2(n_14),
.B1(n_36),
.B2(n_41),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_47),
.B1(n_68),
.B2(n_74),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_8),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_4),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_163),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_170),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_91),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_158),
.C(n_162),
.Y(n_225)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_177),
.B1(n_191),
.B2(n_99),
.Y(n_211)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_50),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_164),
.Y(n_198)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_172),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_1),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_179),
.Y(n_214)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_99),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_2),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_185),
.Y(n_220)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_2),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_187),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_98),
.B(n_80),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_189),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_101),
.B(n_62),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_141),
.B(n_60),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_2),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_150),
.C(n_131),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_151),
.A2(n_46),
.B1(n_28),
.B2(n_21),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_194),
.B1(n_99),
.B2(n_126),
.Y(n_202)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_163),
.CI(n_171),
.CON(n_197),
.SN(n_197)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_197),
.B(n_103),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_132),
.B1(n_111),
.B2(n_146),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_213),
.B1(n_217),
.B2(n_119),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_202),
.A2(n_126),
.B1(n_167),
.B2(n_119),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_205),
.B(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_153),
.A2(n_146),
.B1(n_125),
.B2(n_127),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_139),
.C(n_124),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_130),
.C(n_103),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_158),
.A2(n_145),
.B1(n_127),
.B2(n_147),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_112),
.B(n_131),
.C(n_71),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_149),
.B(n_130),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_139),
.B1(n_133),
.B2(n_104),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_179),
.B1(n_187),
.B2(n_160),
.Y(n_227)
);

NOR2x1_ASAP7_75t_R g226 ( 
.A(n_174),
.B(n_112),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_231),
.B1(n_235),
.B2(n_237),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_174),
.C(n_156),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_233),
.C(n_245),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_238),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_162),
.B(n_154),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_214),
.B(n_201),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_156),
.B1(n_157),
.B2(n_172),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_161),
.C(n_168),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_167),
.B(n_176),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_202),
.B(n_221),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_192),
.B1(n_145),
.B2(n_194),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_182),
.B1(n_169),
.B2(n_155),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_243),
.B1(n_198),
.B2(n_209),
.Y(n_269)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_178),
.B1(n_165),
.B2(n_164),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_246),
.B1(n_211),
.B2(n_223),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_169),
.B1(n_155),
.B2(n_100),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_196),
.C(n_216),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_128),
.B1(n_100),
.B2(n_191),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_219),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_205),
.Y(n_278)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_261),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_258),
.C(n_270),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_221),
.B(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_200),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_200),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_236),
.B1(n_235),
.B2(n_232),
.Y(n_281)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_197),
.Y(n_275)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_238),
.B(n_224),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_277),
.B(n_215),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_205),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_287),
.B1(n_289),
.B2(n_296),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_245),
.C(n_228),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_301),
.C(n_259),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_250),
.B1(n_230),
.B2(n_236),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_293),
.B1(n_258),
.B2(n_254),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_253),
.B1(n_242),
.B2(n_227),
.Y(n_287)
);

XOR2x2_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_231),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_278),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_253),
.B1(n_251),
.B2(n_246),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_263),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_257),
.A2(n_239),
.B1(n_237),
.B2(n_247),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_256),
.B1(n_276),
.B2(n_274),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_251),
.B1(n_241),
.B2(n_226),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_273),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_271),
.B1(n_255),
.B2(n_264),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_215),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_252),
.C(n_244),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_291),
.B1(n_289),
.B2(n_279),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_317),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_309),
.C(n_313),
.Y(n_335)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_284),
.C(n_266),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_259),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_315),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_280),
.C(n_282),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_280),
.A2(n_270),
.B(n_259),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_261),
.C(n_270),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_264),
.C(n_255),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_265),
.C(n_268),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_321),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_265),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_272),
.B1(n_262),
.B2(n_269),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_322),
.A2(n_291),
.B1(n_293),
.B2(n_286),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_272),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_326),
.Y(n_340)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_268),
.B(n_218),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_325),
.A2(n_292),
.B(n_282),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_218),
.C(n_204),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_310),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_337),
.A2(n_347),
.B1(n_311),
.B2(n_315),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_338),
.B(n_343),
.Y(n_357)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_324),
.Y(n_341)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_307),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_348),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_303),
.A2(n_287),
.B1(n_292),
.B2(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_365),
.Y(n_369)
);

BUFx12f_ASAP7_75t_SL g351 ( 
.A(n_328),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_351),
.A2(n_355),
.B(n_361),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_306),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_354),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_319),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_339),
.A2(n_313),
.B(n_320),
.Y(n_355)
);

BUFx12_ASAP7_75t_L g360 ( 
.A(n_346),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_360),
.B(n_367),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_309),
.B(n_300),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_198),
.Y(n_362)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_362),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_363),
.A2(n_329),
.B1(n_331),
.B2(n_344),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_333),
.A2(n_332),
.B(n_341),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_204),
.Y(n_366)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_366),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_209),
.C(n_203),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_347),
.B1(n_337),
.B2(n_332),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_372),
.A2(n_97),
.B1(n_184),
.B2(n_186),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_335),
.C(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_373),
.B(n_375),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_327),
.C(n_345),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_342),
.C(n_336),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_379),
.C(n_381),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_380),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_329),
.C(n_331),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_213),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_203),
.C(n_128),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_356),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_8),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_365),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_396),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_394),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_371),
.A2(n_363),
.B(n_356),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_388),
.A2(n_390),
.B(n_368),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_377),
.A2(n_351),
.B(n_360),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_373),
.B(n_358),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_391),
.B(n_397),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_369),
.A2(n_364),
.B1(n_358),
.B2(n_360),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_392),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_369),
.A2(n_181),
.B1(n_108),
.B2(n_149),
.Y(n_394)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_97),
.C(n_159),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_370),
.C(n_381),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_402),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_370),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_384),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_397),
.C(n_384),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_374),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_380),
.C(n_71),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_405),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_387),
.A2(n_388),
.B(n_389),
.Y(n_405)
);

AOI31xp67_ASAP7_75t_L g409 ( 
.A1(n_386),
.A2(n_9),
.A3(n_11),
.B(n_14),
.Y(n_409)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_409),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_400),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_392),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_414),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_415),
.B1(n_418),
.B2(n_403),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_395),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_394),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_403),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_421),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_416),
.B(n_399),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_423),
.B(n_2),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_9),
.Y(n_423)
);

A2O1A1O1Ixp25_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_84),
.B(n_67),
.C(n_25),
.D(n_24),
.Y(n_424)
);

AOI321xp33_ASAP7_75t_L g427 ( 
.A1(n_424),
.A2(n_28),
.A3(n_25),
.B1(n_41),
.B2(n_23),
.C(n_9),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_412),
.C(n_25),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_426),
.B(n_427),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_420),
.Y(n_430)
);

XOR2x2_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_425),
.Y(n_431)
);

AOI221xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_429),
.B1(n_41),
.B2(n_23),
.C(n_3),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_23),
.C(n_180),
.Y(n_433)
);


endmodule