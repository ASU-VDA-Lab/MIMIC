module fake_netlist_5_2273_n_1566 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1566);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1566;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_1529;
wire n_526;
wire n_677;
wire n_372;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_783;
wire n_555;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_980;
wire n_698;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_1540;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_74),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_82),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_201),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_15),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_270),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_88),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_196),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_312),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_264),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_162),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_30),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_65),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_165),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_255),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_25),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_121),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_324),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_126),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_87),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_274),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_218),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_319),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_328),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_315),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_307),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_71),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_299),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_57),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_89),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_235),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_183),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_203),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_217),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_21),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_273),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_128),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_35),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_254),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_120),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_2),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_338),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_11),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_105),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_137),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_46),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_9),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_5),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_146),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_138),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_241),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_226),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_310),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_181),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_243),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_11),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_48),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_283),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_34),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_213),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_22),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_303),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_109),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_191),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_330),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_271),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_2),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_327),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_282),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_197),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_304),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_169),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_289),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_253),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_230),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_143),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_34),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_15),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_267),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_26),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_228),
.B(n_200),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_309),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_1),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_62),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_131),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_248),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_110),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_12),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_257),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_305),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_250),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_123),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_91),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_168),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_215),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_130),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_221),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_252),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_78),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_186),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_287),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_275),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_268),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_10),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_301),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_56),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_236),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_153),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_149),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_61),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_326),
.B(n_297),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_247),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_163),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_212),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_190),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_288),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_35),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_70),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_229),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_249),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_251),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_292),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_214),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_158),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_174),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_256),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_189),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_147),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_198),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_175),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_127),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_171),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_284),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_210),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_331),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_49),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_232),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_47),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_10),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_302),
.Y(n_487)
);

BUFx5_ASAP7_75t_L g488 ( 
.A(n_205),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_98),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_296),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_337),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_225),
.Y(n_492)
);

INVxp33_ASAP7_75t_R g493 ( 
.A(n_227),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_141),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_14),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_280),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_150),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_58),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_151),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_92),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_68),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_95),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_140),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_103),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_233),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_111),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_244),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_199),
.Y(n_508)
);

CKINVDCx14_ASAP7_75t_R g509 ( 
.A(n_313),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_269),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_194),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_114),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_220),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_122),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_50),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_240),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_135),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_329),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_258),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_142),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_160),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_7),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_260),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_335),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_172),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_336),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_306),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_63),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_180),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_277),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_21),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_293),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_184),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_43),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_51),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_42),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_32),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_222),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_0),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_22),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_155),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_276),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_125),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_242),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_108),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_266),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_224),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_295),
.Y(n_548)
);

BUFx8_ASAP7_75t_SL g549 ( 
.A(n_341),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_36),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_52),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_170),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_115),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_219),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_178),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_148),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_112),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_285),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_102),
.Y(n_559)
);

BUFx5_ASAP7_75t_L g560 ( 
.A(n_24),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_298),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_81),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_202),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_239),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_300),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_290),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_157),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_234),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_18),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_90),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_24),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_107),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_272),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_132),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_144),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_80),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_207),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_145),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_344),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_560),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_560),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_344),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_349),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_413),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_349),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_391),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_349),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_560),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_R g589 ( 
.A1(n_345),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_589)
);

OAI22x1_ASAP7_75t_R g590 ( 
.A1(n_353),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_391),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_438),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_359),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_560),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_500),
.B(n_4),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_411),
.B(n_498),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_560),
.Y(n_597)
);

OA21x2_ASAP7_75t_L g598 ( 
.A1(n_348),
.A2(n_361),
.B(n_358),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_560),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_391),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_385),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_412),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_602)
);

BUFx12f_ASAP7_75t_L g603 ( 
.A(n_357),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_538),
.B(n_6),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_390),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_509),
.B(n_8),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_9),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_359),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_392),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_403),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_366),
.B(n_12),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_433),
.B(n_472),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_461),
.B(n_13),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_426),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_480),
.Y(n_615)
);

CKINVDCx6p67_ASAP7_75t_R g616 ( 
.A(n_387),
.Y(n_616)
);

BUFx8_ASAP7_75t_SL g617 ( 
.A(n_549),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_488),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_382),
.B(n_13),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_435),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_468),
.B(n_14),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

OA21x2_ASAP7_75t_L g624 ( 
.A1(n_368),
.A2(n_16),
.B(n_17),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_525),
.B(n_16),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_355),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_359),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_500),
.B(n_17),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_393),
.Y(n_629)
);

INVx6_ASAP7_75t_L g630 ( 
.A(n_393),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_393),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_488),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_373),
.B(n_18),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_451),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_381),
.B(n_515),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_542),
.B(n_19),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_379),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_545),
.B(n_557),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_488),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_441),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_441),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_485),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_351),
.B(n_19),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_441),
.Y(n_645)
);

BUFx8_ASAP7_75t_SL g646 ( 
.A(n_401),
.Y(n_646)
);

INVx6_ASAP7_75t_L g647 ( 
.A(n_491),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_424),
.B(n_20),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_405),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_407),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_423),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_350),
.B(n_20),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_491),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_495),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_429),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_534),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_464),
.B(n_23),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_491),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_377),
.B(n_23),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_486),
.Y(n_660)
);

AOI22x1_ASAP7_75t_SL g661 ( 
.A1(n_531),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_506),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_522),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_506),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_473),
.B(n_28),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_514),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_383),
.B(n_408),
.Y(n_668)
);

OAI22x1_ASAP7_75t_R g669 ( 
.A1(n_537),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_514),
.Y(n_670)
);

BUFx8_ASAP7_75t_L g671 ( 
.A(n_427),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_370),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_514),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_530),
.Y(n_674)
);

BUFx8_ASAP7_75t_SL g675 ( 
.A(n_374),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_536),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_342),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_539),
.B(n_31),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_540),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_378),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_384),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_550),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_343),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_346),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_440),
.B(n_32),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_569),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_530),
.Y(n_687)
);

OA21x2_ASAP7_75t_L g688 ( 
.A1(n_402),
.A2(n_33),
.B(n_36),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_530),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_571),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_469),
.B(n_37),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_548),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_347),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_496),
.B(n_511),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_548),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_513),
.B(n_38),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_409),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_548),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_SL g699 ( 
.A1(n_395),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_388),
.B(n_39),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_415),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_416),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_352),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_418),
.Y(n_704)
);

CKINVDCx11_ASAP7_75t_R g705 ( 
.A(n_399),
.Y(n_705)
);

NOR2x1_ASAP7_75t_L g706 ( 
.A(n_419),
.B(n_53),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_420),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_388),
.B(n_471),
.Y(n_708)
);

OAI22x1_ASAP7_75t_SL g709 ( 
.A1(n_404),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_354),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_471),
.B(n_43),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_578),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_425),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_434),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_356),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_439),
.Y(n_716)
);

BUFx8_ASAP7_75t_SL g717 ( 
.A(n_414),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_447),
.A2(n_44),
.B(n_45),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_448),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_452),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_460),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_360),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_466),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_467),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_470),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_477),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_508),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_512),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_520),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_521),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_527),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_532),
.Y(n_732)
);

BUFx12f_ASAP7_75t_L g733 ( 
.A(n_362),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_544),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_551),
.B(n_47),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_363),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_516),
.B(n_48),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_516),
.B(n_54),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_579),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_630),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_583),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_583),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_630),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_647),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_617),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_647),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_658),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_583),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_R g749 ( 
.A(n_684),
.B(n_431),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_R g750 ( 
.A(n_626),
.B(n_437),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_675),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_717),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_705),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_693),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_613),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_733),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_R g757 ( 
.A(n_649),
.B(n_364),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_646),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_677),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_683),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_585),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_585),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_703),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_722),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_612),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_603),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_585),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_658),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_582),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_600),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_650),
.Y(n_771)
);

BUFx10_ASAP7_75t_L g772 ( 
.A(n_622),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_710),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_655),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_715),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_587),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_715),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_660),
.B(n_443),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_715),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_736),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_676),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_587),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_736),
.Y(n_783)
);

CKINVDCx8_ASAP7_75t_R g784 ( 
.A(n_607),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_637),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_593),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_682),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_596),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_638),
.B(n_553),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_736),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_593),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_616),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_592),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_615),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_R g795 ( 
.A(n_660),
.B(n_446),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_593),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_584),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_608),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_686),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_608),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_708),
.B(n_578),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_679),
.Y(n_802)
);

CKINVDCx16_ASAP7_75t_R g803 ( 
.A(n_606),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_651),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_635),
.B(n_558),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_679),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_671),
.Y(n_807)
);

XNOR2x2_ASAP7_75t_SL g808 ( 
.A(n_619),
.B(n_493),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_608),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_694),
.B(n_365),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_629),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_629),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_671),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_629),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_727),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_728),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_631),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_729),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_631),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_731),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_604),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_R g822 ( 
.A(n_611),
.B(n_449),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_633),
.B(n_563),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_631),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_627),
.B(n_568),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_716),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_716),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_716),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_672),
.B(n_367),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_640),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_640),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_R g832 ( 
.A(n_737),
.B(n_457),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_640),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_720),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_738),
.B(n_570),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_641),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_720),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_641),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_720),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_641),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_788),
.B(n_602),
.C(n_652),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_749),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_835),
.B(n_627),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_769),
.B(n_657),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_762),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_801),
.B(n_700),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_801),
.B(n_598),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_823),
.B(n_598),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_803),
.B(n_648),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_785),
.B(n_666),
.C(n_625),
.Y(n_850)
);

BUFx6f_ASAP7_75t_SL g851 ( 
.A(n_755),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_767),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_759),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_810),
.B(n_711),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_810),
.B(n_627),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_802),
.B(n_678),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_815),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_776),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_832),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_805),
.B(n_628),
.C(n_595),
.Y(n_860)
);

AO221x1_ASAP7_75t_L g861 ( 
.A1(n_804),
.A2(n_712),
.B1(n_699),
.B2(n_576),
.C(n_577),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_809),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_778),
.B(n_795),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_826),
.B(n_645),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_833),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_806),
.B(n_636),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_757),
.A2(n_502),
.B1(n_533),
.B2(n_510),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_836),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_748),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_748),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_816),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_761),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_829),
.A2(n_668),
.B(n_594),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_761),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_796),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_789),
.B(n_581),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_827),
.B(n_828),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_773),
.B(n_607),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_796),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_800),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_829),
.B(n_597),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_L g882 ( 
.A(n_834),
.B(n_691),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_784),
.B(n_685),
.C(n_659),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_837),
.B(n_599),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_800),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_839),
.B(n_645),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_793),
.B(n_643),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_838),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_794),
.B(n_643),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_760),
.B(n_735),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_818),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_820),
.B(n_696),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_786),
.B(n_645),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_739),
.B(n_586),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_838),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_791),
.B(n_653),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_798),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_770),
.B(n_681),
.C(n_680),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_741),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_811),
.B(n_812),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_741),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_797),
.B(n_735),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_763),
.B(n_697),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_764),
.Y(n_904)
);

BUFx6f_ASAP7_75t_SL g905 ( 
.A(n_755),
.Y(n_905)
);

INVx3_ASAP7_75t_R g906 ( 
.A(n_787),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_799),
.B(n_690),
.C(n_664),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_814),
.B(n_653),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_772),
.B(n_696),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_817),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_819),
.B(n_702),
.C(n_701),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_824),
.B(n_653),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_772),
.B(n_665),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_775),
.B(n_369),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_777),
.B(n_665),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_779),
.B(n_714),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_742),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_742),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_830),
.B(n_580),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_822),
.B(n_561),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_831),
.B(n_580),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_742),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_821),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_740),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_743),
.B(n_591),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_840),
.B(n_662),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_782),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_782),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_780),
.B(n_719),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_782),
.B(n_588),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_744),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_746),
.Y(n_933)
);

NOR2x1p5_ASAP7_75t_L g934 ( 
.A(n_807),
.B(n_601),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_853),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_846),
.B(n_783),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_844),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_860),
.B(n_765),
.C(n_702),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_859),
.B(n_771),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_904),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_854),
.B(n_790),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_860),
.A2(n_575),
.B1(n_781),
.B2(n_774),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_842),
.B(n_745),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_859),
.B(n_750),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_894),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_857),
.B(n_747),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_931),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_933),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_918),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_926),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_856),
.B(n_792),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_931),
.Y(n_952)
);

OAI22xp33_ASAP7_75t_L g953 ( 
.A1(n_867),
.A2(n_881),
.B1(n_883),
.B2(n_884),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_903),
.B(n_813),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_881),
.B(n_572),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_847),
.A2(n_688),
.B1(n_718),
.B2(n_624),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_914),
.B(n_866),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_924),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_918),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_876),
.B(n_721),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_871),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_920),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_878),
.B(n_753),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_863),
.B(n_706),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_851),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_891),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_918),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_920),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_847),
.A2(n_848),
.B1(n_850),
.B2(n_876),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_848),
.A2(n_688),
.B(n_624),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_884),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_922),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_855),
.A2(n_662),
.B(n_588),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_933),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_SL g975 ( 
.A1(n_906),
.A2(n_758),
.B1(n_751),
.B2(n_752),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_909),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_922),
.Y(n_977)
);

NOR2xp67_ASAP7_75t_L g978 ( 
.A(n_883),
.B(n_754),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_902),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_845),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_890),
.B(n_756),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_843),
.B(n_723),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_902),
.B(n_882),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_852),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_900),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_862),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_841),
.A2(n_458),
.B1(n_372),
.B2(n_375),
.Y(n_987)
);

BUFx4f_ASAP7_75t_L g988 ( 
.A(n_933),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_868),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_925),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_873),
.B(n_730),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_861),
.A2(n_718),
.B1(n_726),
.B2(n_618),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_869),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_917),
.B(n_930),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_870),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_919),
.B(n_732),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_887),
.B(n_768),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_864),
.B(n_726),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_SL g999 ( 
.A(n_849),
.B(n_589),
.C(n_766),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_899),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_889),
.B(n_371),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_892),
.B(n_376),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_858),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_865),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_886),
.B(n_701),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_901),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_874),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_897),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_910),
.B(n_704),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_907),
.A2(n_623),
.B1(n_632),
.B2(n_620),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_913),
.B(n_704),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_923),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_928),
.B(n_707),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_929),
.Y(n_1014)
);

CKINVDCx8_ASAP7_75t_R g1015 ( 
.A(n_916),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_932),
.A2(n_808),
.B1(n_669),
.B2(n_590),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_879),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_885),
.Y(n_1018)
);

BUFx8_ASAP7_75t_L g1019 ( 
.A(n_851),
.Y(n_1019)
);

NOR2x1p5_ASAP7_75t_L g1020 ( 
.A(n_898),
.B(n_605),
.Y(n_1020)
);

INVx5_ASAP7_75t_L g1021 ( 
.A(n_888),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_872),
.B(n_614),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_875),
.B(n_707),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_880),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_934),
.B(n_656),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_895),
.B(n_713),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_877),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_921),
.A2(n_386),
.B1(n_389),
.B2(n_380),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_905),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_915),
.B(n_394),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_893),
.B(n_896),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_908),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_912),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_979),
.B(n_911),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_SL g1035 ( 
.A1(n_957),
.A2(n_927),
.B(n_734),
.C(n_713),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_953),
.A2(n_734),
.B(n_689),
.C(n_695),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_970),
.A2(n_991),
.B(n_983),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_947),
.A2(n_662),
.B(n_663),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_936),
.B(n_941),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_1027),
.B(n_396),
.Y(n_1040)
);

BUFx5_ASAP7_75t_L g1041 ( 
.A(n_952),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_962),
.B(n_397),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1031),
.A2(n_667),
.B(n_663),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_SL g1044 ( 
.A1(n_955),
.A2(n_911),
.B(n_898),
.C(n_644),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_937),
.B(n_994),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1011),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_975),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_980),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_968),
.A2(n_639),
.B(n_400),
.C(n_406),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_938),
.B(n_661),
.C(n_410),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_935),
.Y(n_1052)
);

OAI22x1_ASAP7_75t_L g1053 ( 
.A1(n_942),
.A2(n_661),
.B1(n_709),
.B2(n_905),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_961),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_972),
.B(n_398),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_971),
.B(n_417),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_956),
.A2(n_667),
.B(n_663),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_977),
.A2(n_969),
.B(n_960),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_966),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_940),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_SL g1061 ( 
.A(n_939),
.B(n_422),
.C(n_421),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1032),
.A2(n_673),
.B(n_667),
.Y(n_1062)
);

AO31x2_ASAP7_75t_L g1063 ( 
.A1(n_982),
.A2(n_698),
.A3(n_670),
.B(n_610),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_954),
.A2(n_654),
.B(n_610),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_985),
.A2(n_725),
.B1(n_724),
.B2(n_430),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_996),
.A2(n_674),
.B(n_673),
.Y(n_1066)
);

INVx8_ASAP7_75t_L g1067 ( 
.A(n_1025),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1010),
.B(n_428),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_944),
.B(n_621),
.C(n_609),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1027),
.B(n_988),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_998),
.A2(n_674),
.B(n_673),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_976),
.A2(n_609),
.B(n_621),
.C(n_634),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1027),
.A2(n_507),
.B1(n_436),
.B2(n_442),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_959),
.A2(n_687),
.B(n_674),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1009),
.A2(n_634),
.B(n_642),
.C(n_591),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_964),
.A2(n_505),
.B1(n_444),
.B2(n_445),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_981),
.B(n_432),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_986),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1015),
.B(n_450),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_SL g1080 ( 
.A(n_943),
.B(n_965),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1005),
.B(n_453),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_949),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1033),
.B(n_454),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_974),
.B(n_455),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_950),
.B(n_642),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_987),
.B(n_456),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_SL g1087 ( 
.A1(n_1001),
.A2(n_574),
.B(n_573),
.C(n_567),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_989),
.A2(n_825),
.B(n_55),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_1008),
.A2(n_517),
.B(n_462),
.C(n_566),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1022),
.B(n_59),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_L g1091 ( 
.A(n_1025),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_992),
.A2(n_725),
.B1(n_724),
.B2(n_519),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_959),
.A2(n_692),
.B(n_687),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1013),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_958),
.B(n_724),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_949),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1022),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_951),
.B(n_459),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_967),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_R g1100 ( 
.A(n_963),
.B(n_463),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1024),
.A2(n_523),
.B(n_475),
.C(n_476),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1003),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1033),
.B(n_474),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_959),
.A2(n_692),
.B(n_687),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1004),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_993),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1000),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1014),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1017),
.A2(n_524),
.B1(n_479),
.B2(n_565),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_967),
.Y(n_1110)
);

O2A1O1Ixp5_ASAP7_75t_SL g1111 ( 
.A1(n_1002),
.A2(n_725),
.B(n_526),
.C(n_564),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1033),
.B(n_478),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_1019),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_974),
.B(n_692),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_984),
.B(n_481),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_995),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1023),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_974),
.A2(n_483),
.B(n_482),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1054),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1059),
.Y(n_1120)
);

BUFx5_ASAP7_75t_L g1121 ( 
.A(n_1090),
.Y(n_1121)
);

NAND2x1p5_ASAP7_75t_L g1122 ( 
.A(n_1110),
.B(n_948),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_1048),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1047),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1037),
.A2(n_1018),
.B(n_1007),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1090),
.B(n_990),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1041),
.Y(n_1127)
);

OA21x2_ASAP7_75t_L g1128 ( 
.A1(n_1058),
.A2(n_1026),
.B(n_973),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1052),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1057),
.A2(n_1039),
.B(n_1050),
.Y(n_1130)
);

BUFx2_ASAP7_75t_SL g1131 ( 
.A(n_1060),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1102),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_1113),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1088),
.A2(n_997),
.B(n_1028),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1086),
.A2(n_1020),
.B1(n_1012),
.B2(n_978),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1110),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1045),
.B(n_1016),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1041),
.B(n_967),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1111),
.A2(n_1006),
.B(n_1021),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1083),
.A2(n_1012),
.B(n_946),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1110),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1105),
.Y(n_1142)
);

BUFx12f_ASAP7_75t_L g1143 ( 
.A(n_1096),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1096),
.Y(n_1144)
);

AOI22x1_ASAP7_75t_L g1145 ( 
.A1(n_1046),
.A2(n_1029),
.B1(n_541),
.B2(n_535),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1096),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1067),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1036),
.A2(n_1006),
.B(n_1021),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1041),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1095),
.B(n_946),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1085),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1043),
.A2(n_1006),
.B(n_1021),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1041),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1067),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1049),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1078),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1085),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1099),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1106),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1035),
.A2(n_1030),
.B(n_999),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1034),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1116),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1034),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1107),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1117),
.B(n_484),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1097),
.B(n_60),
.Y(n_1166)
);

AO21x2_ASAP7_75t_L g1167 ( 
.A1(n_1044),
.A2(n_1112),
.B(n_1103),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1056),
.B(n_487),
.Y(n_1168)
);

AO21x2_ASAP7_75t_L g1169 ( 
.A1(n_1042),
.A2(n_490),
.B(n_489),
.Y(n_1169)
);

AO21x2_ASAP7_75t_L g1170 ( 
.A1(n_1055),
.A2(n_494),
.B(n_492),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1092),
.A2(n_499),
.B(n_497),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1108),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1072),
.Y(n_1173)
);

BUFx8_ASAP7_75t_SL g1174 ( 
.A(n_1091),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1082),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1089),
.A2(n_64),
.B(n_66),
.Y(n_1176)
);

BUFx2_ASAP7_75t_R g1177 ( 
.A(n_1070),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1101),
.A2(n_1081),
.B(n_1068),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1063),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1062),
.A2(n_67),
.B(n_69),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1066),
.A2(n_503),
.B(n_501),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1094),
.B(n_1019),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1071),
.A2(n_72),
.B(n_73),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1040),
.B(n_75),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1063),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1061),
.B(n_76),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1084),
.B(n_1038),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1114),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1075),
.Y(n_1189)
);

BUFx10_ASAP7_75t_L g1190 ( 
.A(n_1079),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1115),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_SL g1192 ( 
.A(n_1143),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1137),
.B(n_1069),
.Y(n_1193)
);

BUFx10_ASAP7_75t_L g1194 ( 
.A(n_1186),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1127),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1132),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1161),
.A2(n_1077),
.B1(n_1051),
.B2(n_1098),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1136),
.B(n_1074),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1142),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1150),
.B(n_1064),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1136),
.B(n_1093),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1129),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1120),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1156),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1124),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1156),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1159),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1162),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1164),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1129),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1163),
.A2(n_1065),
.B1(n_1109),
.B2(n_1076),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1127),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1124),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1151),
.B(n_1053),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1172),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1155),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1174),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1155),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1163),
.A2(n_1135),
.B1(n_1126),
.B2(n_1166),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1161),
.A2(n_1100),
.B1(n_1073),
.B2(n_1080),
.Y(n_1220)
);

CKINVDCx14_ASAP7_75t_R g1221 ( 
.A(n_1133),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1121),
.A2(n_552),
.B1(n_518),
.B2(n_562),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1125),
.A2(n_1104),
.B(n_1118),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1163),
.A2(n_547),
.B1(n_528),
.B2(n_559),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1163),
.A2(n_1135),
.B1(n_1126),
.B2(n_1166),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1173),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1176),
.A2(n_1063),
.B(n_554),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1143),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1122),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1122),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1126),
.A2(n_556),
.B1(n_555),
.B2(n_546),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1119),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1123),
.A2(n_543),
.B1(n_529),
.B2(n_504),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1149),
.Y(n_1234)
);

INVx4_ASAP7_75t_SL g1235 ( 
.A(n_1166),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1168),
.B(n_77),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1147),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1146),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1147),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1133),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1153),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1153),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1152),
.A2(n_1087),
.B(n_83),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1141),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1136),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1121),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_SL g1247 ( 
.A(n_1154),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1174),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1136),
.Y(n_1249)
);

BUFx8_ASAP7_75t_L g1250 ( 
.A(n_1157),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1176),
.A2(n_86),
.B(n_93),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1144),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1138),
.B(n_94),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1190),
.B(n_96),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1144),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1157),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1123),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1121),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1152),
.A2(n_101),
.B(n_104),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1171),
.A2(n_1121),
.B1(n_1191),
.B2(n_1160),
.Y(n_1260)
);

OR2x6_ASAP7_75t_L g1261 ( 
.A(n_1131),
.B(n_106),
.Y(n_1261)
);

INVx4_ASAP7_75t_SL g1262 ( 
.A(n_1186),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1165),
.B(n_113),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1261),
.B(n_1154),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_R g1265 ( 
.A(n_1192),
.B(n_1190),
.Y(n_1265)
);

AOI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1197),
.A2(n_1178),
.B(n_1169),
.Y(n_1266)
);

CKINVDCx16_ASAP7_75t_R g1267 ( 
.A(n_1217),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1209),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1241),
.A2(n_1130),
.B(n_1138),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1257),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1223),
.A2(n_1134),
.B(n_1180),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1245),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1193),
.B(n_1200),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1199),
.Y(n_1274)
);

NAND2xp33_ASAP7_75t_R g1275 ( 
.A(n_1203),
.B(n_1186),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1209),
.B(n_1160),
.Y(n_1276)
);

INVxp33_ASAP7_75t_SL g1277 ( 
.A(n_1238),
.Y(n_1277)
);

OR2x6_ASAP7_75t_L g1278 ( 
.A(n_1261),
.B(n_1182),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1204),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1219),
.B(n_1140),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1232),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1213),
.B(n_1158),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_1248),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1213),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1219),
.A2(n_1121),
.B1(n_1182),
.B2(n_1189),
.Y(n_1285)
);

NOR2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1202),
.B(n_1188),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_R g1287 ( 
.A(n_1228),
.B(n_1121),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_SL g1288 ( 
.A(n_1220),
.B(n_1184),
.C(n_1187),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1210),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1214),
.B(n_1175),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1240),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1196),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1215),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1233),
.A2(n_1184),
.B1(n_1169),
.B2(n_1170),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1221),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1205),
.B(n_1170),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1206),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1236),
.B(n_1175),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1218),
.B(n_1177),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1233),
.A2(n_1145),
.B1(n_1178),
.B2(n_1130),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_R g1301 ( 
.A(n_1254),
.B(n_1181),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1207),
.B(n_1208),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1252),
.B(n_1188),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1235),
.B(n_1237),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1239),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_R g1306 ( 
.A(n_1261),
.B(n_1181),
.Y(n_1306)
);

AND3x1_ASAP7_75t_L g1307 ( 
.A(n_1260),
.B(n_1179),
.C(n_1185),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1226),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1234),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1225),
.A2(n_1187),
.B1(n_1185),
.B2(n_1179),
.Y(n_1310)
);

OR2x6_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_1183),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1211),
.A2(n_1134),
.B(n_1180),
.C(n_1183),
.Y(n_1312)
);

NOR3xp33_ASAP7_75t_SL g1313 ( 
.A(n_1231),
.B(n_1181),
.C(n_1167),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1216),
.B(n_1167),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1235),
.B(n_1148),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1242),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_L g1317 ( 
.A(n_1258),
.B(n_1128),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1252),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1255),
.B(n_1128),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1231),
.B(n_1139),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1244),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1211),
.A2(n_1148),
.B1(n_1139),
.B2(n_118),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1195),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1263),
.B(n_340),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1262),
.B(n_116),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1250),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1249),
.B(n_1229),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1266),
.A2(n_1243),
.B(n_1259),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1273),
.B(n_1262),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1286),
.B(n_1262),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1305),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1319),
.Y(n_1332)
);

NAND2xp33_ASAP7_75t_R g1333 ( 
.A(n_1287),
.B(n_1251),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1289),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1284),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1296),
.B(n_1212),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1308),
.B(n_1212),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1289),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1277),
.B(n_1194),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1268),
.B(n_1194),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1264),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1298),
.B(n_1230),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1292),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1303),
.B(n_1245),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1293),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1285),
.B(n_1222),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1302),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1299),
.B(n_1245),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1285),
.B(n_1222),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1318),
.B(n_1274),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1279),
.B(n_1246),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1297),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1309),
.B(n_1253),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1321),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1314),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1317),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1316),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1281),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1280),
.B(n_1253),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1282),
.B(n_1227),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1264),
.B(n_1323),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1327),
.B(n_1198),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1280),
.B(n_1227),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1280),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1304),
.B(n_1247),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1317),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1307),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1294),
.B(n_1224),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1307),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1320),
.B(n_1251),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1304),
.Y(n_1372)
);

OAI211xp5_ASAP7_75t_L g1373 ( 
.A1(n_1300),
.A2(n_1256),
.B(n_1247),
.C(n_1250),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1272),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1271),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1272),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1315),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1278),
.B(n_1201),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1288),
.B(n_117),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1265),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1311),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1310),
.Y(n_1382)
);

AND2x4_ASAP7_75t_SL g1383 ( 
.A(n_1315),
.B(n_1311),
.Y(n_1383)
);

NAND2x1_ASAP7_75t_L g1384 ( 
.A(n_1269),
.B(n_119),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1322),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1322),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1324),
.B(n_124),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1325),
.Y(n_1388)
);

NAND4xp25_ASAP7_75t_L g1389 ( 
.A(n_1275),
.B(n_129),
.C(n_133),
.D(n_134),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1270),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1312),
.B(n_136),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1267),
.Y(n_1392)
);

INVx5_ASAP7_75t_L g1393 ( 
.A(n_1306),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1344),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1346),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1355),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1356),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1359),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1334),
.B(n_1313),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1383),
.B(n_1326),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1345),
.B(n_1267),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1383),
.B(n_1301),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1332),
.B(n_1283),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1336),
.B(n_1283),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1381),
.B(n_1295),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1336),
.B(n_1291),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1332),
.B(n_139),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1337),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1357),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1365),
.B(n_152),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1348),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1388),
.B(n_1368),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1381),
.B(n_1370),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1361),
.B(n_154),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1359),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1393),
.B(n_156),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1377),
.B(n_1342),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1342),
.B(n_159),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1382),
.B(n_161),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1357),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1362),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1351),
.B(n_164),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1343),
.B(n_166),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1367),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1375),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1353),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1393),
.B(n_167),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1338),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1393),
.B(n_1367),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1358),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1338),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1393),
.B(n_173),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1364),
.B(n_176),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1331),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1363),
.B(n_177),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1341),
.B(n_179),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1385),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1371),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1371),
.B(n_182),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1342),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1396),
.Y(n_1442)
);

NAND2xp33_ASAP7_75t_R g1443 ( 
.A(n_1402),
.B(n_1330),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1413),
.B(n_1386),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1396),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1439),
.B(n_1360),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1394),
.Y(n_1447)
);

AOI211x1_ASAP7_75t_L g1448 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1373),
.C(n_1369),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1430),
.B(n_1378),
.Y(n_1449)
);

AND2x4_ASAP7_75t_SL g1450 ( 
.A(n_1402),
.B(n_1330),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1409),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1395),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1425),
.B(n_1392),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1430),
.B(n_1329),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1408),
.B(n_1347),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1420),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1421),
.B(n_1349),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1435),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1423),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1397),
.B(n_1350),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1402),
.B(n_1350),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1426),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1398),
.B(n_1331),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1412),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1425),
.B(n_1352),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1416),
.B(n_1342),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1403),
.B(n_1379),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1415),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1399),
.B(n_1369),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1412),
.B(n_1429),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1432),
.B(n_1341),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1438),
.B(n_1411),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1427),
.B(n_1431),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1459),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1465),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1460),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1470),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1442),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1445),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1447),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1473),
.B(n_1427),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1462),
.B(n_1431),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1452),
.Y(n_1485)
);

NOR2x1p5_ASAP7_75t_L g1486 ( 
.A(n_1471),
.B(n_1390),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1453),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1446),
.B(n_1426),
.Y(n_1488)
);

NOR2x1p5_ASAP7_75t_SL g1489 ( 
.A(n_1459),
.B(n_1461),
.Y(n_1489)
);

XNOR2xp5_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_1390),
.Y(n_1490)
);

XOR2x2_ASAP7_75t_L g1491 ( 
.A(n_1448),
.B(n_1401),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1461),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1462),
.B(n_1440),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1464),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1464),
.Y(n_1495)
);

OA222x2_ASAP7_75t_L g1496 ( 
.A1(n_1466),
.A2(n_1434),
.B1(n_1419),
.B2(n_1372),
.C1(n_1391),
.C2(n_1333),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1467),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1491),
.A2(n_1468),
.B1(n_1416),
.B2(n_1443),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1486),
.A2(n_1468),
.B1(n_1443),
.B2(n_1463),
.Y(n_1499)
);

AOI21xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1490),
.A2(n_1406),
.B(n_1469),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1483),
.A2(n_1391),
.B(n_1373),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1480),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1493),
.A2(n_1455),
.B(n_1472),
.Y(n_1503)
);

AOI31xp33_ASAP7_75t_L g1504 ( 
.A1(n_1478),
.A2(n_1400),
.A3(n_1405),
.B(n_1340),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1481),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1496),
.A2(n_1418),
.B(n_1400),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1479),
.A2(n_1418),
.B1(n_1405),
.B2(n_1450),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1482),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1485),
.Y(n_1509)
);

OAI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1484),
.A2(n_1437),
.B1(n_1340),
.B2(n_1422),
.C(n_1436),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_1418),
.B1(n_1449),
.B2(n_1454),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1503),
.B(n_1487),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1508),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1509),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1502),
.Y(n_1515)
);

BUFx2_ASAP7_75t_SL g1516 ( 
.A(n_1498),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_SL g1518 ( 
.A1(n_1500),
.A2(n_1335),
.B(n_1339),
.C(n_1492),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1505),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1501),
.A2(n_1433),
.B1(n_1428),
.B2(n_1424),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1506),
.A2(n_1441),
.B1(n_1474),
.B2(n_1444),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1510),
.B(n_1407),
.C(n_1414),
.D(n_1410),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1504),
.B(n_1380),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1511),
.Y(n_1524)
);

AOI221x1_ASAP7_75t_L g1525 ( 
.A1(n_1516),
.A2(n_1374),
.B1(n_1376),
.B2(n_1475),
.C(n_1407),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1524),
.B(n_1494),
.Y(n_1526)
);

AOI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1521),
.A2(n_1507),
.B(n_1387),
.C(n_1366),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1517),
.B(n_1476),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1518),
.A2(n_1366),
.B(n_1492),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1523),
.B(n_1488),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1515),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1520),
.A2(n_1384),
.B(n_1451),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1531),
.B(n_1530),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1532),
.B(n_1513),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1527),
.A2(n_1522),
.B(n_1519),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1525),
.B(n_1514),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1529),
.A2(n_1526),
.B(n_1533),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1528),
.B(n_1489),
.Y(n_1539)
);

AOI221x1_ASAP7_75t_L g1540 ( 
.A1(n_1538),
.A2(n_1458),
.B1(n_1456),
.B2(n_1417),
.C(n_1354),
.Y(n_1540)
);

AOI321xp33_ASAP7_75t_L g1541 ( 
.A1(n_1534),
.A2(n_1417),
.A3(n_185),
.B1(n_187),
.B2(n_188),
.C(n_192),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1536),
.A2(n_1328),
.B1(n_193),
.B2(n_195),
.Y(n_1542)
);

AOI222xp33_ASAP7_75t_L g1543 ( 
.A1(n_1535),
.A2(n_204),
.B1(n_206),
.B2(n_208),
.C1(n_209),
.C2(n_211),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1537),
.B(n_216),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1540),
.B(n_1539),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1544),
.B(n_1328),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1542),
.A2(n_231),
.B1(n_237),
.B2(n_238),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1541),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_SL g1549 ( 
.A(n_1548),
.B(n_1543),
.C(n_245),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1545),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1550),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1549),
.Y(n_1552)
);

AO22x2_ASAP7_75t_L g1553 ( 
.A1(n_1551),
.A2(n_1546),
.B1(n_1547),
.B2(n_261),
.Y(n_1553)
);

OA22x2_ASAP7_75t_L g1554 ( 
.A1(n_1552),
.A2(n_246),
.B1(n_259),
.B2(n_262),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1554),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1553),
.B(n_263),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1555),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1556),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1557),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1558),
.Y(n_1560)
);

AOI21xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1559),
.A2(n_291),
.B(n_294),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1560),
.B(n_308),
.C(n_311),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1561),
.A2(n_314),
.B1(n_316),
.B2(n_318),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1562),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1563),
.B(n_325),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1565),
.A2(n_1564),
.B1(n_332),
.B2(n_333),
.Y(n_1566)
);


endmodule