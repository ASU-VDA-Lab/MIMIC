module fake_netlist_5_664_n_1606 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1606);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1606;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_67),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_58),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_19),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_27),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_75),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_26),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_38),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_37),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_61),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_91),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_30),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_63),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_35),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_111),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_98),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_81),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_34),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_88),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_38),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_44),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_72),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_25),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_77),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_59),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_26),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_36),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_43),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_104),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_90),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_20),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_56),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_83),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_141),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_28),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_15),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_117),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_140),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_85),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_79),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_44),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_37),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_40),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_73),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_133),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_151),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_106),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_93),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_118),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_96),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_39),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_47),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_49),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_121),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_57),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_54),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_55),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_60),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_12),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_84),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_5),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_41),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_86),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_22),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_45),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_112),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_105),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_20),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_48),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_1),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_27),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_41),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_134),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_24),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_11),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_64),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_19),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_21),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_132),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_107),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_16),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_42),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_122),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_13),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_11),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_46),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_51),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_13),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_39),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_46),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_144),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_68),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_4),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_135),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_65),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_191),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_200),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_203),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_172),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_207),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_214),
.B(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_208),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_194),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_198),
.B(n_4),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_202),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_213),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_219),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_222),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_284),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_229),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_156),
.B(n_7),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

BUFx6f_ASAP7_75t_SL g335 ( 
.A(n_166),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_231),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_288),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_184),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_243),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_247),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_159),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_216),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_216),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_227),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_248),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_179),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_180),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_187),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_185),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_196),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_156),
.B(n_7),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_190),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_227),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_246),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_256),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_220),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_209),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_249),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_186),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_206),
.B(n_8),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_189),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_193),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_195),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_260),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_258),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_273),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_206),
.B(n_8),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_255),
.B(n_306),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_259),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_276),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_220),
.B(n_10),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_199),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_262),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_287),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_234),
.B(n_10),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_293),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_264),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_201),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_204),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_160),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_234),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_196),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_238),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_371),
.A2(n_294),
.B(n_285),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_311),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_152),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_320),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_338),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_384),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_350),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_152),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_360),
.B(n_210),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_363),
.B(n_211),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_307),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_364),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_255),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_365),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_332),
.B(n_306),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_285),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_322),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_313),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_387),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_316),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_382),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_383),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_307),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_317),
.B(n_153),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_329),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_308),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_308),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_310),
.B(n_294),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_352),
.B(n_361),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_309),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_356),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_309),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_312),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_337),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_312),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_319),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_319),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_323),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_323),
.Y(n_454)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_386),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_324),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_324),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_379),
.B(n_154),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_326),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_326),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_416),
.B(n_358),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_416),
.B(n_421),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_390),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_424),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_409),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_435),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_381),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_434),
.A2(n_321),
.B1(n_318),
.B2(n_370),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_390),
.B(n_331),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_394),
.B(n_318),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

NOR2x1p5_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_331),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_351),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_409),
.B(n_336),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_413),
.B(n_336),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_432),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_401),
.B(n_333),
.C(n_362),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_397),
.B(n_339),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_397),
.B(n_339),
.Y(n_484)
);

BUFx6f_ASAP7_75t_SL g485 ( 
.A(n_412),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_422),
.B(n_340),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_422),
.B(n_340),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_433),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_388),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_401),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_388),
.A2(n_374),
.B1(n_378),
.B2(n_296),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_430),
.B(n_265),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx4_ASAP7_75t_SL g499 ( 
.A(n_399),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_458),
.B(n_265),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_388),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_429),
.B(n_345),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_405),
.B(n_345),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_455),
.B(n_314),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_430),
.B(n_265),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_393),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_458),
.A2(n_299),
.B(n_298),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_403),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_443),
.B(n_359),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_458),
.A2(n_412),
.B1(n_441),
.B2(n_451),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_435),
.B(n_265),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_395),
.B(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_395),
.B(n_368),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_400),
.B(n_368),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_372),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_438),
.B(n_265),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_438),
.B(n_157),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_412),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_400),
.B(n_372),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_438),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_441),
.A2(n_303),
.B1(n_335),
.B2(n_304),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_455),
.B(n_224),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_406),
.B(n_376),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_406),
.B(n_376),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_441),
.B(n_242),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_439),
.B(n_380),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_441),
.A2(n_335),
.B1(n_192),
.B2(n_275),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_439),
.B(n_380),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_455),
.B(n_162),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_398),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_407),
.Y(n_544)
);

OAI21xp33_ASAP7_75t_SL g545 ( 
.A1(n_425),
.A2(n_427),
.B(n_426),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_437),
.B(n_375),
.Y(n_546)
);

AND3x2_ASAP7_75t_L g547 ( 
.A(n_442),
.B(n_188),
.C(n_167),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_442),
.A2(n_335),
.B1(n_181),
.B2(n_176),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_407),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_170),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_398),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_456),
.A2(n_181),
.B1(n_176),
.B2(n_174),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_456),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_402),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_389),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_455),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_439),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_455),
.A2(n_297),
.B1(n_301),
.B2(n_305),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_402),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_451),
.A2(n_197),
.B1(n_177),
.B2(n_205),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_448),
.B(n_212),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_407),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_415),
.B(n_217),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_448),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_451),
.B(n_160),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_431),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_448),
.B(n_215),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_402),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_417),
.B(n_218),
.Y(n_574)
);

NOR2x1p5_ASAP7_75t_L g575 ( 
.A(n_449),
.B(n_163),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_452),
.B(n_153),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_448),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_411),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_453),
.B(n_280),
.Y(n_579)
);

INVxp33_ASAP7_75t_L g580 ( 
.A(n_404),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_450),
.A2(n_232),
.B1(n_237),
.B2(n_263),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_425),
.B(n_166),
.Y(n_582)
);

OAI21xp33_ASAP7_75t_SL g583 ( 
.A1(n_426),
.A2(n_251),
.B(n_257),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_454),
.B(n_305),
.C(n_292),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_457),
.B(n_459),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_411),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_460),
.B(n_155),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_450),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_450),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_446),
.B(n_221),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_450),
.B(n_223),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_446),
.B(n_169),
.C(n_292),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_411),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_427),
.B(n_166),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_418),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_464),
.B(n_225),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_392),
.C(n_420),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_467),
.A2(n_494),
.B1(n_465),
.B2(n_492),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_469),
.B(n_396),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_482),
.B(n_226),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_471),
.B(n_155),
.Y(n_602)
);

AND2x6_ASAP7_75t_SL g603 ( 
.A(n_502),
.B(n_233),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_461),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_484),
.B(n_431),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_511),
.B(n_408),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_508),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_525),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_511),
.B(n_410),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_469),
.B(n_477),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_491),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_556),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_486),
.B(n_158),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_509),
.Y(n_614)
);

BUFx6f_ASAP7_75t_SL g615 ( 
.A(n_556),
.Y(n_615)
);

AO221x1_ASAP7_75t_L g616 ( 
.A1(n_561),
.A2(n_283),
.B1(n_250),
.B2(n_418),
.C(n_446),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_513),
.B(n_431),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_487),
.B(n_230),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_463),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_515),
.B(n_158),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_477),
.B(n_235),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_479),
.B(n_419),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_465),
.A2(n_494),
.B1(n_501),
.B2(n_490),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_537),
.B(n_236),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_480),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_537),
.B(n_239),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_479),
.B(n_240),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_473),
.B(n_163),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_491),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_517),
.B(n_161),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_519),
.B(n_161),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_470),
.B(n_164),
.C(n_168),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_539),
.B(n_233),
.Y(n_633)
);

INVxp33_ASAP7_75t_L g634 ( 
.A(n_473),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_489),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_558),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_538),
.A2(n_254),
.B1(n_241),
.B2(n_244),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_465),
.A2(n_494),
.B1(n_507),
.B2(n_550),
.Y(n_638)
);

INVx8_ASAP7_75t_L g639 ( 
.A(n_506),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_580),
.B(n_168),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_498),
.B(n_245),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_526),
.B(n_534),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_504),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_493),
.B(n_250),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_507),
.A2(n_550),
.B1(n_493),
.B2(n_500),
.Y(n_645)
);

BUFx8_ASAP7_75t_L g646 ( 
.A(n_585),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_550),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_535),
.B(n_174),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_576),
.B(n_269),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_590),
.B(n_252),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_570),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_582),
.B(n_269),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_590),
.B(n_253),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_566),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_559),
.B(n_278),
.Y(n_656)
);

AO221x1_ASAP7_75t_L g657 ( 
.A1(n_566),
.A2(n_283),
.B1(n_233),
.B2(n_277),
.C(n_175),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_587),
.B(n_278),
.Y(n_658)
);

INVx8_ASAP7_75t_L g659 ( 
.A(n_506),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_590),
.B(n_261),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_550),
.A2(n_282),
.B1(n_171),
.B2(n_175),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_582),
.B(n_266),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_570),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_538),
.B(n_169),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_594),
.B(n_300),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_530),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_595),
.B(n_594),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_550),
.B(n_302),
.Y(n_669)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_476),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_506),
.A2(n_281),
.B1(n_178),
.B2(n_182),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_595),
.B(n_283),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_541),
.B(n_171),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_182),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_567),
.B(n_183),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_545),
.B(n_282),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_550),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_574),
.B(n_183),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_476),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_591),
.B(n_268),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_510),
.A2(n_444),
.B(n_423),
.C(n_414),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_466),
.Y(n_682)
);

AND2x6_ASAP7_75t_SL g683 ( 
.A(n_512),
.B(n_277),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_518),
.B(n_281),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_485),
.A2(n_481),
.B1(n_506),
.B2(n_542),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_528),
.B(n_271),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_522),
.A2(n_551),
.B(n_568),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_466),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_472),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_543),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_527),
.B(n_286),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_554),
.B(n_274),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_472),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_536),
.B(n_274),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_536),
.B(n_279),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_503),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_542),
.B(n_80),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_500),
.A2(n_291),
.B1(n_290),
.B2(n_289),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_505),
.B(n_286),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_555),
.B(n_289),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_539),
.B(n_497),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_529),
.B(n_277),
.Y(n_702)
);

NOR2x1p5_ASAP7_75t_L g703 ( 
.A(n_546),
.B(n_592),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g704 ( 
.A(n_521),
.B(n_391),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_546),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_548),
.B(n_17),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_579),
.B(n_17),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_552),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_503),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_540),
.B(n_22),
.C(n_23),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_557),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_557),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_485),
.A2(n_69),
.B1(n_146),
.B2(n_139),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_475),
.B(n_25),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_542),
.B(n_62),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_583),
.B(n_28),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_563),
.A2(n_560),
.B(n_553),
.C(n_589),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_532),
.B(n_29),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_485),
.B(n_29),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_542),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_532),
.B(n_31),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_500),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_575),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_532),
.B(n_33),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_462),
.B(n_94),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_562),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_532),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_468),
.B(n_483),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_462),
.B(n_549),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_581),
.A2(n_92),
.B1(n_136),
.B2(n_129),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_562),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_547),
.B(n_102),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_614),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_614),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_617),
.A2(n_565),
.B(n_520),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_642),
.B(n_531),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_642),
.B(n_531),
.Y(n_737)
);

OAI21xp33_ASAP7_75t_L g738 ( 
.A1(n_602),
.A2(n_692),
.B(n_699),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_638),
.A2(n_588),
.B(n_577),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_623),
.A2(n_572),
.B1(n_564),
.B2(n_523),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_598),
.B(n_593),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_598),
.B(n_593),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_676),
.A2(n_572),
.B(n_564),
.C(n_524),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_623),
.B(n_586),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_629),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_722),
.A2(n_514),
.B1(n_523),
.B2(n_569),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_722),
.A2(n_514),
.B1(n_578),
.B2(n_573),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_644),
.A2(n_586),
.B1(n_578),
.B2(n_573),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_644),
.A2(n_474),
.B1(n_549),
.B2(n_533),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_613),
.A2(n_500),
.B1(n_524),
.B2(n_478),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_613),
.B(n_649),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_729),
.A2(n_468),
.B(n_488),
.Y(n_752)
);

OAI22x1_ASAP7_75t_L g753 ( 
.A1(n_706),
.A2(n_40),
.B1(n_42),
.B2(n_47),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_665),
.A2(n_478),
.B(n_549),
.C(n_533),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_612),
.B(n_500),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_687),
.A2(n_488),
.B(n_571),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_611),
.B(n_652),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_638),
.A2(n_478),
.B(n_531),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_639),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_649),
.B(n_533),
.Y(n_760)
);

AOI21x1_ASAP7_75t_L g761 ( 
.A1(n_711),
.A2(n_726),
.B(n_712),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_692),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.C(n_52),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_676),
.A2(n_500),
.B(n_52),
.C(n_53),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_636),
.Y(n_764)
);

OAI21xp33_ASAP7_75t_L g765 ( 
.A1(n_699),
.A2(n_50),
.B(n_53),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_701),
.B(n_499),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_664),
.B(n_499),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_706),
.A2(n_661),
.B1(n_665),
.B2(n_673),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_673),
.A2(n_571),
.B(n_544),
.C(n_496),
.Y(n_769)
);

AND2x6_ASAP7_75t_L g770 ( 
.A(n_697),
.B(n_108),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_647),
.A2(n_680),
.B(n_717),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_655),
.A2(n_571),
.B(n_544),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_658),
.B(n_620),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_618),
.B(n_496),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_SL g775 ( 
.A(n_606),
.B(n_495),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_645),
.A2(n_495),
.B(n_115),
.Y(n_776)
);

AOI21x1_ASAP7_75t_L g777 ( 
.A1(n_731),
.A2(n_495),
.B(n_119),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_674),
.A2(n_110),
.B(n_120),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_SL g779 ( 
.A(n_609),
.B(n_127),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_674),
.A2(n_149),
.B(n_648),
.C(n_630),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_604),
.B(n_619),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_599),
.B(n_631),
.Y(n_782)
);

INVx11_ASAP7_75t_L g783 ( 
.A(n_646),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_639),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_631),
.A2(n_648),
.B1(n_601),
.B2(n_607),
.Y(n_785)
);

BUFx8_ASAP7_75t_SL g786 ( 
.A(n_615),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_625),
.B(n_635),
.Y(n_787)
);

BUFx4f_ASAP7_75t_SL g788 ( 
.A(n_646),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_663),
.Y(n_789)
);

CKINVDCx10_ASAP7_75t_R g790 ( 
.A(n_615),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_633),
.B(n_679),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_663),
.B(n_643),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_622),
.B(n_670),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_632),
.B(n_596),
.C(n_705),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_650),
.B(n_608),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_675),
.B(n_678),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_671),
.B(n_656),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_667),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_651),
.A2(n_654),
.B(n_660),
.Y(n_799)
);

AO21x1_ASAP7_75t_L g800 ( 
.A1(n_624),
.A2(n_626),
.B(n_725),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_661),
.A2(n_698),
.B1(n_718),
.B2(n_697),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_720),
.Y(n_802)
);

OAI321xp33_ASAP7_75t_L g803 ( 
.A1(n_710),
.A2(n_698),
.A3(n_707),
.B1(n_716),
.B2(n_628),
.C(n_721),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_686),
.B(n_695),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_694),
.B(n_700),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_715),
.A2(n_685),
.B1(n_720),
.B2(n_721),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_690),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_634),
.B(n_640),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_639),
.B(n_659),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_721),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_641),
.A2(n_669),
.B(n_672),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_659),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_621),
.Y(n_813)
);

OAI321xp33_ASAP7_75t_L g814 ( 
.A1(n_600),
.A2(n_702),
.A3(n_714),
.B1(n_626),
.B2(n_624),
.C(n_621),
.Y(n_814)
);

AOI33xp33_ASAP7_75t_L g815 ( 
.A1(n_723),
.A2(n_681),
.A3(n_724),
.B1(n_732),
.B2(n_637),
.B3(n_715),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_682),
.A2(n_688),
.B(n_696),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_708),
.B(n_689),
.Y(n_817)
);

OAI21xp33_ASAP7_75t_L g818 ( 
.A1(n_653),
.A2(n_600),
.B(n_627),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_627),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_693),
.A2(n_709),
.B(n_708),
.Y(n_820)
);

AO21x1_ASAP7_75t_L g821 ( 
.A1(n_730),
.A2(n_684),
.B(n_691),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_727),
.B(n_703),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_662),
.A2(n_666),
.B(n_677),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_704),
.B(n_719),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_713),
.A2(n_732),
.B(n_616),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_L g827 ( 
.A1(n_597),
.A2(n_657),
.B(n_683),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_603),
.B(n_642),
.Y(n_828)
);

AO21x1_ASAP7_75t_L g829 ( 
.A1(n_602),
.A2(n_673),
.B(n_665),
.Y(n_829)
);

OAI21xp33_ASAP7_75t_L g830 ( 
.A1(n_602),
.A2(n_470),
.B(n_692),
.Y(n_830)
);

AOI221xp5_ASAP7_75t_SL g831 ( 
.A1(n_676),
.A2(n_434),
.B1(n_470),
.B2(n_467),
.C(n_510),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_642),
.B(n_464),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_642),
.B(n_464),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_642),
.B(n_416),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_629),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_676),
.A2(n_434),
.B(n_664),
.C(n_652),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_642),
.B(n_464),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_642),
.B(n_598),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_676),
.A2(n_434),
.B(n_664),
.C(n_652),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_642),
.B(n_598),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_617),
.A2(n_668),
.B(n_605),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_610),
.B(n_559),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_642),
.B(n_416),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_617),
.A2(n_668),
.B(n_605),
.Y(n_844)
);

AOI21x1_ASAP7_75t_L g845 ( 
.A1(n_728),
.A2(n_605),
.B(n_668),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_610),
.B(n_469),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_617),
.A2(n_668),
.B(n_605),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_642),
.B(n_464),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_642),
.B(n_464),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_642),
.B(n_464),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_642),
.B(n_464),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_602),
.B(n_416),
.C(n_387),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_602),
.A2(n_642),
.B(n_673),
.C(n_665),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_599),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_676),
.A2(n_434),
.B(n_664),
.C(n_652),
.Y(n_855)
);

NAND2x2_ASAP7_75t_L g856 ( 
.A(n_703),
.B(n_475),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_629),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_642),
.B(n_464),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_617),
.A2(n_668),
.B(n_605),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_602),
.B(n_416),
.C(n_387),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_642),
.B(n_416),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_623),
.A2(n_598),
.B1(n_722),
.B2(n_470),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_617),
.A2(n_668),
.B(n_605),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_617),
.A2(n_668),
.B(n_605),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_604),
.B(n_511),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_642),
.B(n_416),
.Y(n_866)
);

OAI21xp33_ASAP7_75t_L g867 ( 
.A1(n_602),
.A2(n_470),
.B(n_692),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_642),
.A2(n_602),
.B1(n_610),
.B2(n_464),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_642),
.B(n_598),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_663),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_602),
.A2(n_642),
.B(n_673),
.C(n_665),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_642),
.B(n_464),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_701),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_642),
.B(n_464),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_873),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_764),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_834),
.B(n_843),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_807),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_832),
.B(n_833),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_853),
.A2(n_871),
.B(n_751),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_861),
.B(n_866),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_768),
.A2(n_738),
.B1(n_830),
.B2(n_867),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_859),
.A2(n_864),
.B(n_863),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_789),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_770),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_741),
.A2(n_742),
.B(n_774),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_846),
.B(n_791),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_768),
.A2(n_773),
.B1(n_862),
.B2(n_782),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_837),
.B(n_850),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_733),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_838),
.A2(n_869),
.B(n_840),
.C(n_862),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_798),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_759),
.B(n_784),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_734),
.Y(n_896)
);

AOI21xp33_ASAP7_75t_L g897 ( 
.A1(n_829),
.A2(n_801),
.B(n_796),
.Y(n_897)
);

NOR2x1_ASAP7_75t_R g898 ( 
.A(n_825),
.B(n_854),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_819),
.A2(n_813),
.B1(n_818),
.B2(n_869),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_838),
.A2(n_840),
.B(n_736),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_793),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_851),
.B(n_858),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_857),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_872),
.A2(n_874),
.B(n_765),
.C(n_868),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_789),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_822),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_770),
.B(n_780),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_737),
.A2(n_742),
.B(n_741),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_744),
.A2(n_740),
.B(n_739),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_789),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_845),
.A2(n_771),
.B(n_816),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_744),
.A2(n_740),
.B(n_799),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_811),
.A2(n_760),
.B(n_805),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_848),
.B(n_849),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_786),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_759),
.B(n_784),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_852),
.B(n_860),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_822),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_804),
.B(n_831),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_820),
.A2(n_756),
.B(n_758),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_SL g921 ( 
.A(n_812),
.B(n_870),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_762),
.A2(n_803),
.B(n_855),
.C(n_839),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_776),
.A2(n_754),
.B(n_746),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_814),
.B(n_785),
.Y(n_924)
);

AND3x4_ASAP7_75t_L g925 ( 
.A(n_781),
.B(n_865),
.C(n_842),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_842),
.B(n_792),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_870),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_817),
.A2(n_777),
.B(n_772),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_745),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_802),
.Y(n_930)
);

AO31x2_ASAP7_75t_L g931 ( 
.A1(n_800),
.A2(n_821),
.A3(n_748),
.B(n_769),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_836),
.A2(n_815),
.B(n_743),
.C(n_824),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_792),
.B(n_787),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_795),
.B(n_766),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_808),
.A2(n_835),
.B(n_753),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_812),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_746),
.A2(n_747),
.B(n_749),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_870),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_806),
.A2(n_794),
.B1(n_797),
.B2(n_750),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_802),
.B(n_810),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_802),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_757),
.Y(n_942)
);

AOI21x1_ASAP7_75t_SL g943 ( 
.A1(n_755),
.A2(n_826),
.B(n_778),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_775),
.A2(n_806),
.B(n_779),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_767),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_770),
.B(n_823),
.Y(n_946)
);

INVx4_ASAP7_75t_SL g947 ( 
.A(n_770),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_770),
.B(n_828),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_763),
.A2(n_827),
.B(n_856),
.C(n_809),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_812),
.B(n_809),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_809),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_790),
.A2(n_783),
.B(n_788),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_853),
.A2(n_871),
.B(n_751),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_798),
.Y(n_954)
);

OAI222xp33_ASAP7_75t_L g955 ( 
.A1(n_768),
.A2(n_862),
.B1(n_751),
.B2(n_773),
.C1(n_801),
.C2(n_840),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_789),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_853),
.A2(n_871),
.B(n_751),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_853),
.B(n_871),
.Y(n_959)
);

OAI22x1_ASAP7_75t_L g960 ( 
.A1(n_834),
.A2(n_843),
.B1(n_866),
.B2(n_861),
.Y(n_960)
);

AOI21xp33_ASAP7_75t_L g961 ( 
.A1(n_738),
.A2(n_843),
.B(n_834),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_832),
.B(n_872),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_832),
.B(n_872),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_968)
);

AND3x2_ASAP7_75t_L g969 ( 
.A(n_762),
.B(n_719),
.C(n_834),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_832),
.B(n_872),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_972)
);

OAI21x1_ASAP7_75t_SL g973 ( 
.A1(n_824),
.A2(n_799),
.B(n_800),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_SL g974 ( 
.A1(n_862),
.A2(n_871),
.B(n_853),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_853),
.A2(n_871),
.B(n_751),
.Y(n_977)
);

AO31x2_ASAP7_75t_L g978 ( 
.A1(n_829),
.A2(n_768),
.A3(n_800),
.B(n_853),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_980)
);

OAI22xp33_ASAP7_75t_L g981 ( 
.A1(n_862),
.A2(n_768),
.B1(n_751),
.B2(n_773),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_807),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_759),
.B(n_784),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_807),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_751),
.B(n_773),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_738),
.A2(n_853),
.B(n_871),
.C(n_867),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_768),
.A2(n_862),
.B1(n_867),
.B2(n_830),
.Y(n_988)
);

BUFx4f_ASAP7_75t_SL g989 ( 
.A(n_812),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_853),
.A2(n_871),
.B(n_830),
.C(n_867),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_832),
.B(n_872),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_995)
);

AO21x1_ASAP7_75t_L g996 ( 
.A1(n_768),
.A2(n_751),
.B(n_773),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_798),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_768),
.A2(n_751),
.B(n_773),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_735),
.A2(n_761),
.B(n_752),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_834),
.Y(n_1000)
);

BUFx8_ASAP7_75t_L g1001 ( 
.A(n_810),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_841),
.A2(n_847),
.B(n_844),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_857),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_875),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_1000),
.B(n_877),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_887),
.B(n_921),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_878),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_882),
.B(n_902),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_889),
.B(n_901),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_902),
.B(n_986),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_961),
.B(n_884),
.C(n_988),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_986),
.B(n_880),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1000),
.B(n_960),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_917),
.B(n_891),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_981),
.A2(n_890),
.B1(n_925),
.B2(n_988),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_962),
.B(n_965),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_971),
.B(n_994),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_936),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_903),
.Y(n_1020)
);

AO21x1_ASAP7_75t_L g1021 ( 
.A1(n_981),
.A2(n_924),
.B(n_959),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_876),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_895),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_933),
.B(n_893),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_875),
.B(n_926),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_982),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_1004),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_906),
.B(n_929),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_1003),
.A2(n_879),
.B(n_995),
.Y(n_1029)
);

OA21x2_ASAP7_75t_L g1030 ( 
.A1(n_923),
.A2(n_937),
.B(n_912),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_936),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_984),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_895),
.B(n_916),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_987),
.A2(n_991),
.B1(n_881),
.B2(n_953),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_940),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_989),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_936),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_1002),
.A2(n_979),
.B(n_995),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_929),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_892),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_930),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_925),
.A2(n_907),
.B1(n_969),
.B2(n_948),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_996),
.B(n_998),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_991),
.B(n_900),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_896),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_887),
.B(n_916),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_899),
.B(n_914),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_894),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_954),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_983),
.B(n_918),
.Y(n_1050)
);

OA21x2_ASAP7_75t_L g1051 ( 
.A1(n_909),
.A2(n_967),
.B(n_966),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_941),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_997),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_969),
.A2(n_939),
.B1(n_935),
.B2(n_914),
.Y(n_1054)
);

BUFx12f_ASAP7_75t_L g1055 ( 
.A(n_1001),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_958),
.B(n_977),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_922),
.A2(n_955),
.B(n_924),
.C(n_959),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_904),
.B(n_934),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_1001),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_989),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_SL g1061 ( 
.A(n_887),
.B(n_946),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_887),
.B(n_955),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_904),
.B(n_919),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_942),
.A2(n_944),
.B1(n_922),
.B2(n_951),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_945),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_983),
.B(n_941),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_886),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_974),
.A2(n_908),
.B1(n_932),
.B2(n_913),
.Y(n_1068)
);

AO21x1_ASAP7_75t_L g1069 ( 
.A1(n_885),
.A2(n_979),
.B(n_972),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_949),
.B(n_967),
.C(n_972),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_910),
.B(n_938),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_910),
.B(n_938),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_SL g1073 ( 
.A(n_950),
.B(n_888),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_927),
.B(n_978),
.Y(n_1074)
);

BUFx2_ASAP7_75t_R g1075 ( 
.A(n_915),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_927),
.B(n_978),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_978),
.B(n_898),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_886),
.A2(n_905),
.B1(n_957),
.B2(n_968),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_949),
.A2(n_970),
.B(n_920),
.C(n_911),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_905),
.A2(n_957),
.B1(n_947),
.B2(n_973),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_978),
.B(n_947),
.Y(n_1081)
);

INVx5_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_931),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_931),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_931),
.B(n_928),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_931),
.A2(n_952),
.B(n_883),
.C(n_956),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_963),
.B(n_964),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_975),
.Y(n_1088)
);

AOI21xp33_ASAP7_75t_L g1089 ( 
.A1(n_976),
.A2(n_980),
.B(n_985),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_990),
.B(n_992),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_993),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_999),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_887),
.B(n_921),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_882),
.B(n_834),
.Y(n_1094)
);

O2A1O1Ixp5_ASAP7_75t_SL g1095 ( 
.A1(n_924),
.A2(n_959),
.B(n_768),
.C(n_897),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_902),
.B(n_986),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_878),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_871),
.B(n_853),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_895),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_875),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_961),
.B(n_867),
.C(n_830),
.Y(n_1101)
);

OAI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_877),
.A2(n_751),
.B1(n_773),
.B2(n_461),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_L g1103 ( 
.A(n_960),
.B(n_853),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_981),
.A2(n_768),
.B(n_960),
.Y(n_1104)
);

INVx8_ASAP7_75t_L g1105 ( 
.A(n_895),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1004),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_878),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_1001),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_923),
.A2(n_937),
.B(n_912),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_902),
.B(n_986),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_878),
.Y(n_1111)
);

NOR2x1_ASAP7_75t_SL g1112 ( 
.A(n_887),
.B(n_862),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_876),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_902),
.B(n_986),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_991),
.A2(n_871),
.B(n_853),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_989),
.B(n_389),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_991),
.A2(n_871),
.B(n_853),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_944),
.B(n_809),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_878),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_882),
.B(n_877),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_1001),
.Y(n_1121)
);

OR2x2_ASAP7_75t_SL g1122 ( 
.A(n_877),
.B(n_917),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_902),
.B(n_986),
.Y(n_1123)
);

AOI222xp33_ASAP7_75t_L g1124 ( 
.A1(n_1012),
.A2(n_1034),
.B1(n_1098),
.B2(n_1115),
.C1(n_1117),
.C2(n_1015),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_1020),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1016),
.B(n_1101),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1008),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1017),
.A2(n_1018),
.B1(n_1009),
.B2(n_1122),
.Y(n_1128)
);

OAI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1062),
.A2(n_1054),
.B1(n_1017),
.B2(n_1018),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1094),
.B(n_1010),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1105),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1019),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1042),
.A2(n_1102),
.B1(n_1006),
.B2(n_1047),
.Y(n_1133)
);

CKINVDCx8_ASAP7_75t_R g1134 ( 
.A(n_1113),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1120),
.A2(n_1064),
.B1(n_1096),
.B2(n_1123),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1011),
.B(n_1096),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1055),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1104),
.A2(n_1034),
.B1(n_1117),
.B2(n_1115),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1032),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1011),
.A2(n_1123),
.B1(n_1114),
.B2(n_1110),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1039),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1062),
.A2(n_1056),
.B1(n_1098),
.B2(n_1110),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1019),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1097),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_1108),
.Y(n_1145)
);

OAI22xp33_ASAP7_75t_R g1146 ( 
.A1(n_1028),
.A2(n_1005),
.B1(n_1100),
.B2(n_1106),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1107),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1114),
.A2(n_1077),
.B1(n_1056),
.B2(n_1013),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1111),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_1118),
.B(n_1086),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1119),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1040),
.Y(n_1152)
);

AO21x2_ASAP7_75t_L g1153 ( 
.A1(n_1089),
.A2(n_1038),
.B(n_1029),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1045),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1065),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1035),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1025),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1118),
.B(n_1033),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1103),
.A2(n_1109),
.B1(n_1030),
.B2(n_1116),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1013),
.A2(n_1024),
.B1(n_1058),
.B2(n_1118),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1024),
.B(n_1057),
.Y(n_1161)
);

BUFx8_ASAP7_75t_L g1162 ( 
.A(n_1121),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1030),
.A2(n_1109),
.B1(n_1014),
.B2(n_1112),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1104),
.A2(n_1021),
.B1(n_1068),
.B2(n_1063),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1049),
.Y(n_1165)
);

INVx6_ASAP7_75t_L g1166 ( 
.A(n_1105),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1105),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1053),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1051),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1051),
.Y(n_1170)
);

CKINVDCx11_ASAP7_75t_R g1171 ( 
.A(n_1060),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1027),
.B(n_1044),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_SL g1173 ( 
.A1(n_1068),
.A2(n_1070),
.B1(n_1022),
.B2(n_1082),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1081),
.B(n_1074),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1043),
.A2(n_1048),
.B1(n_1082),
.B2(n_1083),
.Y(n_1175)
);

INVx6_ASAP7_75t_L g1176 ( 
.A(n_1033),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1076),
.B(n_1043),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1071),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1072),
.Y(n_1179)
);

CKINVDCx11_ASAP7_75t_R g1180 ( 
.A(n_1059),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1082),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1041),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1052),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1073),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1041),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1007),
.A2(n_1093),
.B1(n_1080),
.B2(n_1099),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1036),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1095),
.B(n_1084),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1023),
.A2(n_1099),
.B1(n_1082),
.B2(n_1050),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1061),
.A2(n_1083),
.B1(n_1050),
.B2(n_1078),
.Y(n_1190)
);

BUFx8_ASAP7_75t_SL g1191 ( 
.A(n_1031),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1083),
.A2(n_1078),
.B1(n_1046),
.B2(n_1066),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1067),
.A2(n_1037),
.B1(n_1090),
.B2(n_1087),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1067),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1085),
.A2(n_1092),
.B1(n_1091),
.B2(n_1088),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1079),
.B(n_1069),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1197)
);

INVx6_ASAP7_75t_L g1198 ( 
.A(n_1019),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1116),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_1104),
.A2(n_768),
.B(n_981),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1118),
.B(n_974),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_1113),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1015),
.A2(n_830),
.B1(n_867),
.B2(n_738),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1020),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1101),
.A2(n_768),
.B1(n_867),
.B2(n_830),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1094),
.B(n_1010),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1016),
.B(n_1101),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1105),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1105),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1020),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1007),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1026),
.Y(n_1212)
);

INVx8_ASAP7_75t_L g1213 ( 
.A(n_1105),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1015),
.B(n_882),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1020),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1026),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1025),
.B(n_1120),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1039),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1015),
.B(n_882),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1015),
.A2(n_834),
.B1(n_861),
.B2(n_843),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1026),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1113),
.Y(n_1223)
);

OAI22x1_ASAP7_75t_L g1224 ( 
.A1(n_1054),
.A2(n_1016),
.B1(n_884),
.B2(n_890),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1157),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1219),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1215),
.B(n_1220),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1169),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1200),
.A2(n_1196),
.A3(n_1224),
.B(n_1170),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1174),
.B(n_1136),
.Y(n_1230)
);

OAI21xp33_ASAP7_75t_L g1231 ( 
.A1(n_1221),
.A2(n_1203),
.B(n_1205),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1201),
.B(n_1158),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1185),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1177),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1174),
.B(n_1136),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1201),
.B(n_1150),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1148),
.B(n_1140),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1188),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1205),
.A2(n_1124),
.B(n_1173),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1183),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1126),
.B(n_1207),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1141),
.Y(n_1242)
);

AO21x1_ASAP7_75t_SL g1243 ( 
.A1(n_1175),
.A2(n_1164),
.B(n_1138),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1126),
.B(n_1207),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1201),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1163),
.B(n_1138),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1172),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1159),
.B(n_1224),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1153),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1160),
.B(n_1128),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1182),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1184),
.A2(n_1181),
.B(n_1164),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1171),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1130),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1153),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1189),
.A2(n_1175),
.B(n_1186),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1150),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1155),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1127),
.Y(n_1259)
);

NOR3xp33_ASAP7_75t_L g1260 ( 
.A(n_1129),
.B(n_1135),
.C(n_1133),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1166),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1139),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1194),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1144),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_1161),
.B2(n_1142),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1147),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1149),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1195),
.A2(n_1142),
.B(n_1151),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1166),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1152),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1154),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1178),
.A2(n_1179),
.B(n_1206),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1218),
.B(n_1222),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1195),
.A2(n_1165),
.B(n_1168),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1204),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1212),
.B(n_1217),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1125),
.B(n_1216),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1190),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1197),
.B(n_1192),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1210),
.B(n_1214),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1193),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1211),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1171),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1228),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1275),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1238),
.B(n_1156),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1260),
.A2(n_1132),
.B(n_1143),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1247),
.B(n_1132),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1234),
.B(n_1229),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1274),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1234),
.B(n_1229),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1229),
.B(n_1167),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1229),
.B(n_1167),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1274),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1229),
.B(n_1249),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1245),
.B(n_1236),
.Y(n_1296)
);

OR2x6_ASAP7_75t_L g1297 ( 
.A(n_1236),
.B(n_1213),
.Y(n_1297)
);

AND2x4_ASAP7_75t_SL g1298 ( 
.A(n_1236),
.B(n_1223),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1229),
.B(n_1176),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1249),
.B(n_1187),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1230),
.B(n_1176),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1249),
.B(n_1223),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1255),
.B(n_1223),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1237),
.B(n_1198),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1255),
.B(n_1202),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1239),
.A2(n_1199),
.B1(n_1134),
.B2(n_1198),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1255),
.B(n_1202),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1236),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1235),
.B(n_1131),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1235),
.B(n_1245),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1236),
.B(n_1268),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1274),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1268),
.B(n_1202),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1237),
.B(n_1199),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1285),
.B(n_1225),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1314),
.B(n_1227),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1306),
.A2(n_1231),
.B1(n_1265),
.B2(n_1248),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1285),
.B(n_1233),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1310),
.B(n_1248),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1288),
.B(n_1241),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1310),
.B(n_1257),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1306),
.A2(n_1231),
.B1(n_1278),
.B2(n_1244),
.Y(n_1322)
);

NAND4xp25_ASAP7_75t_L g1323 ( 
.A(n_1314),
.B(n_1272),
.C(n_1244),
.D(n_1277),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1302),
.B(n_1257),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1302),
.B(n_1240),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1297),
.A2(n_1250),
.B(n_1268),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1313),
.A2(n_1250),
.B(n_1246),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1287),
.B(n_1232),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1313),
.A2(n_1232),
.B1(n_1246),
.B2(n_1278),
.Y(n_1329)
);

AND2x2_ASAP7_75t_SL g1330 ( 
.A(n_1308),
.B(n_1232),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1301),
.B(n_1254),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1284),
.Y(n_1332)
);

AOI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1313),
.A2(n_1281),
.B(n_1279),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1302),
.B(n_1226),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1301),
.B(n_1283),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1303),
.B(n_1251),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1303),
.B(n_1257),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1313),
.B(n_1281),
.C(n_1242),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1287),
.B(n_1263),
.C(n_1273),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1303),
.B(n_1273),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1303),
.B(n_1267),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1290),
.B(n_1282),
.C(n_1279),
.Y(n_1342)
);

OA211x2_ASAP7_75t_L g1343 ( 
.A1(n_1304),
.A2(n_1243),
.B(n_1283),
.C(n_1162),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1305),
.B(n_1267),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1305),
.B(n_1232),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1305),
.B(n_1267),
.Y(n_1346)
);

OAI21xp33_ASAP7_75t_L g1347 ( 
.A1(n_1311),
.A2(n_1276),
.B(n_1256),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1305),
.B(n_1275),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_L g1349 ( 
.A(n_1290),
.B(n_1280),
.C(n_1266),
.Y(n_1349)
);

OAI21xp33_ASAP7_75t_L g1350 ( 
.A1(n_1311),
.A2(n_1276),
.B(n_1256),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_L g1351 ( 
.A1(n_1294),
.A2(n_1270),
.B1(n_1271),
.B2(n_1266),
.C(n_1264),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1294),
.B(n_1280),
.C(n_1262),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1307),
.B(n_1258),
.Y(n_1353)
);

OAI221xp5_ASAP7_75t_L g1354 ( 
.A1(n_1304),
.A2(n_1253),
.B1(n_1134),
.B2(n_1261),
.C(n_1187),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1307),
.B(n_1252),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1299),
.B(n_1252),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1299),
.B(n_1259),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1286),
.B(n_1259),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1319),
.B(n_1311),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1332),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1357),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1319),
.B(n_1311),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1320),
.B(n_1289),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1357),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1356),
.B(n_1295),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1358),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1355),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1341),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1347),
.B(n_1291),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1344),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1353),
.B(n_1292),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1347),
.B(n_1308),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1351),
.B(n_1292),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1346),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1350),
.B(n_1308),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1355),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1350),
.B(n_1293),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1317),
.A2(n_1286),
.B1(n_1312),
.B2(n_1297),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1321),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1349),
.B(n_1312),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1330),
.B(n_1293),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1330),
.B(n_1293),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1330),
.B(n_1296),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1324),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1323),
.B(n_1286),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1340),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1337),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1386),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1385),
.B(n_1316),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1360),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1385),
.B(n_1334),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1361),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1386),
.B(n_1354),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1360),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1383),
.B(n_1296),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1366),
.B(n_1348),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1361),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1359),
.B(n_1345),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_1383),
.B(n_1338),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1361),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1366),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_1380),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1360),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1318),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1370),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1364),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1364),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1373),
.B(n_1315),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1386),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1360),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1368),
.B(n_1336),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1364),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_SL g1413 ( 
.A(n_1381),
.B(n_1338),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1368),
.B(n_1374),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1371),
.B(n_1325),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1359),
.B(n_1345),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1359),
.B(n_1296),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1374),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1374),
.B(n_1335),
.Y(n_1420)
);

AOI32xp33_ASAP7_75t_L g1421 ( 
.A1(n_1378),
.A2(n_1322),
.A3(n_1329),
.B1(n_1328),
.B2(n_1331),
.Y(n_1421)
);

OAI21xp33_ASAP7_75t_L g1422 ( 
.A1(n_1378),
.A2(n_1317),
.B(n_1327),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1370),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1380),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1363),
.B(n_1339),
.Y(n_1425)
);

NAND2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1381),
.B(n_1309),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1422),
.A2(n_1343),
.B1(n_1339),
.B2(n_1342),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1393),
.B(n_1362),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1395),
.B(n_1362),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1392),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1399),
.A2(n_1326),
.B1(n_1333),
.B2(n_1297),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1392),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1390),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1390),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1418),
.Y(n_1435)
);

AOI21xp33_ASAP7_75t_L g1436 ( 
.A1(n_1422),
.A2(n_1300),
.B(n_1372),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1405),
.B(n_1363),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1397),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1389),
.B(n_1362),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1397),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1400),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1395),
.B(n_1377),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1413),
.A2(n_1352),
.B(n_1349),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1418),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1391),
.B(n_1369),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1400),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1406),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1406),
.Y(n_1448)
);

AND2x4_ASAP7_75t_SL g1449 ( 
.A(n_1395),
.B(n_1381),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1394),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1395),
.B(n_1377),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1404),
.B(n_1369),
.Y(n_1452)
);

NOR2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1402),
.B(n_1137),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1407),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1407),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1412),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1420),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1412),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1413),
.B(n_1377),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1394),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1403),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_L g1462 ( 
.A(n_1399),
.B(n_1352),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1403),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1404),
.B(n_1369),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1408),
.B(n_1372),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1417),
.B(n_1382),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1417),
.B(n_1382),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1408),
.B(n_1137),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1425),
.B(n_1372),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1452),
.B(n_1409),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1424),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1449),
.B(n_1398),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1435),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1462),
.B(n_1410),
.Y(n_1474)
);

NOR2x1_ASAP7_75t_L g1475 ( 
.A(n_1453),
.B(n_1443),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1430),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1459),
.B(n_1398),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1436),
.B(n_1421),
.C(n_1401),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1459),
.B(n_1416),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1457),
.B(n_1428),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1435),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1444),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1444),
.Y(n_1483)
);

NOR2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1469),
.B(n_1269),
.Y(n_1484)
);

NOR2x1_ASAP7_75t_L g1485 ( 
.A(n_1468),
.B(n_1388),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1433),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1416),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1466),
.B(n_1423),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1439),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1464),
.B(n_1414),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1433),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1467),
.B(n_1382),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1434),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1427),
.B(n_1410),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1467),
.B(n_1365),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1447),
.B(n_1415),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1430),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1437),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1437),
.B(n_1415),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1432),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1442),
.B(n_1365),
.Y(n_1502)
);

CKINVDCx16_ASAP7_75t_R g1503 ( 
.A(n_1442),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1432),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1438),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1480),
.B(n_1145),
.Y(n_1506)
);

NAND2x1_ASAP7_75t_L g1507 ( 
.A(n_1474),
.B(n_1451),
.Y(n_1507)
);

AOI322xp5_ASAP7_75t_L g1508 ( 
.A1(n_1494),
.A2(n_1431),
.A3(n_1451),
.B1(n_1375),
.B2(n_1426),
.C1(n_1429),
.C2(n_1365),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1476),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1475),
.B(n_1421),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1482),
.B(n_1429),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1476),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1478),
.A2(n_1375),
.B1(n_1376),
.B2(n_1367),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1481),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1498),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1503),
.B(n_1396),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1498),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1494),
.A2(n_1375),
.B1(n_1343),
.B2(n_1387),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1478),
.A2(n_1297),
.B1(n_1296),
.B2(n_1298),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1482),
.B(n_1411),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1501),
.Y(n_1521)
);

NAND2x1_ASAP7_75t_L g1522 ( 
.A(n_1474),
.B(n_1454),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1475),
.A2(n_1456),
.B(n_1455),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1503),
.A2(n_1298),
.B1(n_1440),
.B2(n_1441),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1501),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1505),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1485),
.A2(n_1387),
.B1(n_1371),
.B2(n_1384),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1505),
.Y(n_1528)
);

NOR3xp33_ASAP7_75t_L g1529 ( 
.A(n_1483),
.B(n_1180),
.C(n_1460),
.Y(n_1529)
);

XOR2x2_ASAP7_75t_L g1530 ( 
.A(n_1485),
.B(n_1145),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1473),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1531),
.B(n_1499),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1509),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1510),
.B(n_1499),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1518),
.B(n_1483),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1483),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1530),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1529),
.B(n_1471),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1507),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1515),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1517),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1521),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1518),
.A2(n_1471),
.B1(n_1484),
.B2(n_1488),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1525),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1526),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1483),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1519),
.B(n_1472),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1545),
.B(n_1527),
.Y(n_1552)
);

NAND4xp25_ASAP7_75t_L g1553 ( 
.A(n_1539),
.B(n_1538),
.C(n_1540),
.D(n_1536),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1541),
.A2(n_1527),
.B1(n_1522),
.B2(n_1524),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1538),
.B(n_1489),
.Y(n_1556)
);

O2A1O1Ixp5_ASAP7_75t_L g1557 ( 
.A1(n_1537),
.A2(n_1513),
.B(n_1523),
.C(n_1474),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1549),
.B(n_1477),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_L g1559 ( 
.A1(n_1537),
.A2(n_1508),
.B(n_1528),
.C(n_1504),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1550),
.A2(n_1474),
.B1(n_1477),
.B2(n_1479),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1532),
.B(n_1489),
.Y(n_1561)
);

OAI211xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1533),
.A2(n_1546),
.B(n_1535),
.C(n_1542),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1551),
.A2(n_1504),
.B(n_1496),
.Y(n_1563)
);

AO22x2_ASAP7_75t_L g1564 ( 
.A1(n_1559),
.A2(n_1548),
.B1(n_1534),
.B2(n_1543),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_L g1565 ( 
.A(n_1553),
.B(n_1544),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1558),
.Y(n_1566)
);

NAND3xp33_ASAP7_75t_L g1567 ( 
.A(n_1557),
.B(n_1547),
.C(n_1496),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1563),
.B(n_1486),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1554),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1556),
.Y(n_1570)
);

AOI221xp5_ASAP7_75t_L g1571 ( 
.A1(n_1552),
.A2(n_1497),
.B1(n_1486),
.B2(n_1493),
.C(n_1491),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1561),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1560),
.Y(n_1573)
);

NOR2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1566),
.B(n_1562),
.Y(n_1574)
);

OAI221xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1567),
.A2(n_1555),
.B1(n_1470),
.B2(n_1500),
.C(n_1479),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1565),
.B(n_1491),
.C(n_1486),
.Y(n_1576)
);

XNOR2x2_ASAP7_75t_L g1577 ( 
.A(n_1564),
.B(n_1472),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1573),
.B(n_1487),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1572),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1578),
.A2(n_1564),
.B1(n_1569),
.B2(n_1570),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1577),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1576),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1579),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1574),
.A2(n_1568),
.B1(n_1571),
.B2(n_1484),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1575),
.B(n_1487),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1578),
.A2(n_1491),
.B1(n_1493),
.B2(n_1490),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1581),
.A2(n_1493),
.B1(n_1500),
.B2(n_1497),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1583),
.B(n_1492),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1580),
.A2(n_1490),
.B1(n_1492),
.B2(n_1502),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1582),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1585),
.A2(n_1440),
.B(n_1438),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1588),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1590),
.B(n_1584),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1591),
.Y(n_1594)
);

AOI22x1_ASAP7_75t_L g1595 ( 
.A1(n_1594),
.A2(n_1587),
.B1(n_1145),
.B2(n_1162),
.Y(n_1595)
);

AOI221x1_ASAP7_75t_L g1596 ( 
.A1(n_1595),
.A2(n_1592),
.B1(n_1593),
.B2(n_1586),
.C(n_1589),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1596),
.A2(n_1593),
.B1(n_1162),
.B2(n_1180),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1596),
.A2(n_1450),
.B1(n_1434),
.B2(n_1461),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1597),
.A2(n_1463),
.B(n_1460),
.Y(n_1599)
);

XNOR2xp5_ASAP7_75t_L g1600 ( 
.A(n_1598),
.B(n_1502),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1600),
.A2(n_1495),
.B1(n_1448),
.B2(n_1441),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1599),
.A2(n_1463),
.B(n_1461),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1601),
.A2(n_1458),
.B1(n_1448),
.B2(n_1450),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1603),
.B(n_1602),
.C(n_1458),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_R g1605 ( 
.A1(n_1604),
.A2(n_1213),
.B1(n_1191),
.B2(n_1495),
.C(n_1419),
.Y(n_1605)
);

AOI211xp5_ASAP7_75t_L g1606 ( 
.A1(n_1605),
.A2(n_1131),
.B(n_1209),
.C(n_1208),
.Y(n_1606)
);


endmodule