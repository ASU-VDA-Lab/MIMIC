module fake_jpeg_4340_n_210 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_210);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_32),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_6),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_6),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_28),
.B1(n_19),
.B2(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_72),
.B1(n_27),
.B2(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_54),
.B(n_56),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_16),
.B1(n_28),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_59),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_24),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_62),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_16),
.B1(n_18),
.B2(n_31),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_61),
.Y(n_112)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_73),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_21),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_28),
.B1(n_19),
.B2(n_29),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_76),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_21),
.B1(n_31),
.B2(n_18),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_83),
.B1(n_8),
.B2(n_12),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_26),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_39),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_17),
.Y(n_84)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_18),
.B1(n_27),
.B2(n_17),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_103),
.B1(n_80),
.B2(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_93),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_0),
.C(n_1),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_110),
.C(n_77),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_83),
.B1(n_82),
.B2(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_62),
.B1(n_64),
.B2(n_53),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_48),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_108),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_10),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_3),
.C(n_12),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_129),
.B1(n_102),
.B2(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_121),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_85),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_53),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_63),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_49),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_50),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_66),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_104),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_112),
.A3(n_105),
.B1(n_107),
.B2(n_61),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_157),
.A3(n_153),
.B1(n_125),
.B2(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_96),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_86),
.B1(n_102),
.B2(n_90),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_102),
.B1(n_105),
.B2(n_112),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_49),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_166),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_148),
.B(n_152),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_114),
.B1(n_135),
.B2(n_127),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_168),
.B1(n_144),
.B2(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_132),
.B(n_131),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_174),
.B(n_160),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_124),
.B1(n_128),
.B2(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_122),
.C(n_133),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_171),
.C(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_116),
.C(n_117),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_137),
.A3(n_49),
.B1(n_61),
.B2(n_70),
.C1(n_67),
.C2(n_60),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_154),
.C(n_150),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_88),
.B1(n_87),
.B2(n_61),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_145),
.C(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_165),
.B1(n_144),
.B2(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_171),
.C(n_169),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_166),
.C(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.C(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_159),
.C(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_159),
.C(n_174),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_194),
.C(n_187),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_147),
.C(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_193),
.A2(n_183),
.B1(n_181),
.B2(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_198),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_197),
.B(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_149),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_191),
.B(n_179),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_158),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_207),
.Y(n_210)
);


endmodule