module real_jpeg_5484_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_1),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_1),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_1),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_1),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_1),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_2),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_2),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_3),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_4),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_5),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_59),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_8),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_9),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_9),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_9),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_9),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_9),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_9),
.B(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_11),
.Y(n_200)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_12),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_13),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_13),
.B(n_57),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_13),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_13),
.B(n_269),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_14),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_15),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_15),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_15),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_15),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_205),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_204),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_159),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_19),
.B(n_159),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.C(n_129),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_20),
.B(n_106),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_21),
.B(n_71),
.C(n_91),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.C(n_55),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_22),
.B(n_55),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_29),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_30),
.C(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_28),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_33),
.Y(n_140)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_33),
.Y(n_175)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_34),
.Y(n_228)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_34),
.Y(n_273)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_37),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_38),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_39),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.C(n_50),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_40),
.A2(n_50),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_40),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_44),
.B(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_49),
.Y(n_292)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_101),
.Y(n_100)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_51),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_54),
.B(n_87),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.C(n_66),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_56),
.A2(n_66),
.B1(n_185),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_56),
.Y(n_346)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_60),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_61),
.B(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_62),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_62),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_66),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_66),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_69),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_91),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_81),
.C(n_86),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_72),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_78),
.Y(n_331)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_80),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_80),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_81),
.B(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_93),
.B(n_95),
.C(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_104),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_97),
.A2(n_98),
.B1(n_104),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_98),
.B(n_166),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_98),
.B(n_166),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_104),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_108),
.B(n_109),
.C(n_117),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_110),
.Y(n_163)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_115),
.C(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_127),
.B2(n_128),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_121),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_120),
.A2(n_121),
.B1(n_214),
.B2(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_123),
.C(n_127),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_121),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_123),
.A2(n_126),
.B1(n_148),
.B2(n_149),
.Y(n_320)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_129),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_152),
.C(n_157),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_130),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_146),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_131),
.B(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_135),
.A2(n_146),
.B1(n_147),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_135),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_136),
.A2(n_141),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_136),
.Y(n_317)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_139),
.B(n_316),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_141),
.Y(n_318)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_152),
.B(n_157),
.Y(n_362)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_159),
.Y(n_376)
);

FAx1_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_187),
.CI(n_203),
.CON(n_159),
.SN(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_180),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_169),
.Y(n_258)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_176),
.Y(n_179)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_202),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_201),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_199),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_357),
.B(n_372),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_337),
.B(n_356),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_310),
.B(n_336),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_263),
.B(n_309),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_249),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_211),
.B(n_249),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_223),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_212),
.B(n_224),
.C(n_236),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_219),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_213),
.B(n_220),
.C(n_222),
.Y(n_324)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_236),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.C(n_231),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_239),
.C(n_248),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_262),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_253),
.B1(n_262),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_255),
.B1(n_259),
.B2(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_303),
.B(n_308),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_288),
.B(n_302),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_277),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_274),
.C(n_276),
.Y(n_304)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_296),
.B(n_301),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_300),
.Y(n_301)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_312),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_324),
.C(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_320),
.C(n_321),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_335),
.Y(n_325)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_332),
.B2(n_334),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_334),
.C(n_335),
.Y(n_341)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_355),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_355),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_349),
.B2(n_354),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_350),
.C(n_351),
.Y(n_367)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_344),
.C(n_347),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_348),
.Y(n_342)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_344),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_349),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_368),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_367),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_367),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_364),
.C(n_365),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_368),
.A2(n_374),
.B(n_375),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_370),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);


endmodule