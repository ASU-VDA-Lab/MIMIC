module fake_jpeg_28911_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_30),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_7),
.B(n_8),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_19),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_24),
.B1(n_18),
.B2(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_17),
.B(n_18),
.C(n_24),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_53),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_54),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_19),
.C(n_13),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_27),
.C(n_14),
.Y(n_59)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_31),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_32),
.B1(n_35),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_13),
.B1(n_14),
.B2(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_67),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_34),
.B1(n_38),
.B2(n_21),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_9),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_8),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_40),
.B1(n_55),
.B2(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_43),
.C(n_11),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_66),
.B1(n_65),
.B2(n_60),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_40),
.C(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_82),
.Y(n_104)
);

FAx1_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_72),
.CI(n_67),
.CON(n_91),
.SN(n_91)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_64),
.B1(n_73),
.B2(n_71),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_102),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_75),
.B1(n_83),
.B2(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_104),
.B1(n_91),
.B2(n_88),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_96),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_88),
.B1(n_91),
.B2(n_75),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_100),
.A3(n_98),
.B1(n_105),
.B2(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_114),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_107),
.Y(n_115)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_98),
.A3(n_76),
.B1(n_92),
.B2(n_64),
.C(n_42),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_110),
.B(n_106),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_116),
.C(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_61),
.C(n_71),
.Y(n_121)
);


endmodule