module real_jpeg_23107_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_1),
.A2(n_53),
.B(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_1),
.B(n_42),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_163),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_30),
.C(n_65),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_1),
.B(n_87),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_1),
.A2(n_27),
.B1(n_250),
.B2(n_257),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_43),
.B1(n_46),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_54),
.B1(n_111),
.B2(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_156),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_156),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_38),
.B1(n_43),
.B2(n_46),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_43),
.B1(n_46),
.B2(n_70),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_49),
.B1(n_54),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_10),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_10),
.A2(n_43),
.B1(n_46),
.B2(n_166),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_166),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_166),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_43),
.B1(n_46),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_11),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_89),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_11),
.A2(n_89),
.B1(n_111),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_89),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_13),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_13),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_13),
.A2(n_43),
.B1(n_46),
.B2(n_109),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_109),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_109),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_49),
.B1(n_54),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_14),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_43),
.B1(n_46),
.B2(n_57),
.Y(n_117)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_138),
.B1(n_139),
.B2(n_314),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_18),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_118),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_21),
.B(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_93),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_22),
.A2(n_23),
.B1(n_73),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_59),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_58),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_25),
.A2(n_58),
.B(n_59),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_25),
.A2(n_26),
.B1(n_60),
.B2(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_27),
.A2(n_36),
.B(n_150),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_27),
.A2(n_98),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_27),
.A2(n_33),
.B1(n_247),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_28),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_28),
.A2(n_149),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_28),
.A2(n_246),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_29),
.A2(n_30),
.B1(n_65),
.B2(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_29),
.B(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_31),
.B(n_101),
.Y(n_150)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_32),
.Y(n_99)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_37),
.B(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_51),
.B(n_55),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_40),
.A2(n_108),
.B(n_113),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_40),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_40),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_40),
.A2(n_42),
.B1(n_165),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_40),
.A2(n_42),
.B1(n_108),
.B2(n_173),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_41),
.B(n_52),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_41),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_41),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_46),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_43),
.A2(n_47),
.B(n_162),
.C(n_180),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_43),
.B(n_163),
.CON(n_208),
.SN(n_208)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_45),
.B(n_46),
.C(n_112),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_46),
.A2(n_64),
.A3(n_86),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_50),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_71),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_69),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_71),
.B(n_78),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_61),
.A2(n_106),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_61),
.A2(n_76),
.B(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_61),
.A2(n_106),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_61),
.A2(n_106),
.B1(n_213),
.B2(n_232),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_64),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_63),
.B(n_85),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_64),
.B(n_234),
.Y(n_233)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_77),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_68),
.A2(n_79),
.B(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_68),
.B(n_163),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_73),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_81),
.B(n_92),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_91),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_82),
.A2(n_157),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_82),
.A2(n_91),
.B1(n_155),
.B2(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_82),
.A2(n_132),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_83),
.A2(n_87),
.B1(n_199),
.B2(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_87),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_87),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_91),
.B(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_119),
.CI(n_136),
.CON(n_118),
.SN(n_118)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_93),
.A2(n_94),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_107),
.C(n_114),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_95),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_100),
.A2(n_184),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_107),
.A2(n_114),
.B1(n_115),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_107),
.Y(n_302)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_118),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_307),
.B(n_313),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_294),
.B(n_306),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_200),
.B(n_277),
.C(n_293),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_186),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_169),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_151),
.B1(n_167),
.B2(n_168),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_145),
.B(n_168),
.C(n_169),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_146),
.B(n_147),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_163),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_172),
.B(n_174),
.C(n_178),
.Y(n_291)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_187),
.B(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_190),
.B(n_192),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_195),
.B1(n_196),
.B2(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_272),
.B(n_276),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_226),
.B(n_271),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_205),
.B(n_215),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_212),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_210),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_212),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_223),
.C(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_266),
.B(n_270),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_243),
.B(n_265),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_229),
.B(n_235),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_253),
.B(n_264),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_252),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_263),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_256),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_279),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_291),
.B2(n_292),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_283),
.C(n_292),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_287),
.C(n_290),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_305),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_300),
.B1(n_303),
.B2(n_304),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_304),
.C(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);


endmodule