module real_aes_16404_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_0), .Y(n_550) );
AND2x4_ASAP7_75t_L g851 ( .A(n_1), .B(n_852), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_2), .A2(n_4), .B1(n_275), .B2(n_276), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_3), .A2(n_21), .B1(n_202), .B2(n_211), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_5), .A2(n_51), .B1(n_160), .B2(n_161), .Y(n_159) );
BUFx3_ASAP7_75t_L g501 ( .A(n_6), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_7), .A2(n_15), .B1(n_132), .B2(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g852 ( .A(n_8), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_9), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_10), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_11), .B(n_185), .Y(n_507) );
OR2x2_ASAP7_75t_L g109 ( .A(n_12), .B(n_30), .Y(n_109) );
BUFx2_ASAP7_75t_L g846 ( .A(n_12), .Y(n_846) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_13), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_14), .Y(n_835) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_16), .B(n_167), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_17), .B(n_176), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_18), .A2(n_84), .B1(n_167), .B2(n_211), .Y(n_565) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_19), .A2(n_46), .B(n_145), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_20), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_22), .B(n_202), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_23), .B(n_137), .Y(n_231) );
INVx4_ASAP7_75t_R g184 ( .A(n_24), .Y(n_184) );
AO32x2_ASAP7_75t_L g562 ( .A1(n_25), .A2(n_213), .A3(n_214), .B1(n_563), .B2(n_566), .Y(n_562) );
AO32x1_ASAP7_75t_L g584 ( .A1(n_25), .A2(n_213), .A3(n_214), .B1(n_563), .B2(n_566), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_26), .B(n_202), .Y(n_237) );
INVx1_ASAP7_75t_L g280 ( .A(n_27), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_SL g208 ( .A1(n_28), .A2(n_132), .B(n_136), .C(n_209), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_29), .A2(n_43), .B1(n_132), .B2(n_139), .Y(n_220) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_30), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_31), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_32), .A2(n_50), .B1(n_186), .B2(n_202), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_33), .A2(n_89), .B1(n_139), .B2(n_211), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_34), .B(n_509), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_35), .B(n_531), .Y(n_575) );
INVx1_ASAP7_75t_L g234 ( .A(n_36), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_37), .B(n_132), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_38), .A2(n_66), .B1(n_139), .B2(n_556), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_39), .Y(n_253) );
INVx2_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
INVx1_ASAP7_75t_L g107 ( .A(n_41), .Y(n_107) );
BUFx3_ASAP7_75t_L g117 ( .A(n_41), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_42), .B(n_577), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_44), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_45), .A2(n_83), .B1(n_132), .B2(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_47), .B(n_825), .Y(n_824) );
OAI31xp67_ASAP7_75t_SL g830 ( .A1(n_47), .A2(n_826), .A3(n_828), .B(n_831), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_48), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_49), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_52), .A2(n_77), .B1(n_169), .B2(n_531), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_53), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_54), .A2(n_81), .B1(n_167), .B2(n_211), .Y(n_497) );
INVx1_ASAP7_75t_L g145 ( .A(n_55), .Y(n_145) );
AND2x4_ASAP7_75t_L g147 ( .A(n_56), .B(n_148), .Y(n_147) );
XNOR2xp5_ASAP7_75t_L g118 ( .A(n_57), .B(n_119), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_58), .A2(n_88), .B1(n_139), .B2(n_273), .Y(n_272) );
AO22x1_ASAP7_75t_L g165 ( .A1(n_59), .A2(n_72), .B1(n_166), .B2(n_168), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_60), .B(n_211), .Y(n_506) );
INVx1_ASAP7_75t_L g148 ( .A(n_61), .Y(n_148) );
AND2x2_ASAP7_75t_L g212 ( .A(n_62), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_63), .B(n_213), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_64), .A2(n_157), .B(n_160), .C(n_549), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_65), .B(n_211), .C(n_511), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_67), .A2(n_100), .B1(n_842), .B2(n_853), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_68), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_69), .B(n_160), .Y(n_259) );
AND2x2_ASAP7_75t_L g551 ( .A(n_70), .B(n_190), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_71), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_73), .B(n_202), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_74), .A2(n_94), .B1(n_167), .B2(n_169), .Y(n_533) );
INVx2_ASAP7_75t_L g137 ( .A(n_75), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_76), .B(n_255), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_78), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_79), .B(n_213), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_80), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_82), .B(n_143), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_85), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_86), .A2(n_98), .B1(n_139), .B2(n_186), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_87), .B(n_531), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_90), .B(n_213), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_91), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g486 ( .A(n_91), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_92), .B(n_176), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_93), .A2(n_141), .B(n_160), .C(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g189 ( .A(n_95), .B(n_190), .Y(n_189) );
NAND2xp33_ASAP7_75t_L g258 ( .A(n_96), .B(n_185), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_97), .Y(n_520) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_110), .Y(n_100) );
INVxp67_ASAP7_75t_L g831 ( .A(n_101), .Y(n_831) );
NOR2x1_ASAP7_75t_R g101 ( .A(n_102), .B(n_103), .Y(n_101) );
INVx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx8_ASAP7_75t_R g827 ( .A(n_104), .Y(n_827) );
AND2x6_ASAP7_75t_SL g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_107), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_108), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x1_ASAP7_75t_L g841 ( .A(n_109), .B(n_117), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_118), .B(n_822), .Y(n_110) );
INVx4_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x6_ASAP7_75t_SL g112 ( .A(n_113), .B(n_115), .Y(n_112) );
BUFx3_ASAP7_75t_L g833 ( .A(n_113), .Y(n_833) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_114), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_483), .B1(n_487), .B2(n_821), .Y(n_119) );
INVx2_ASAP7_75t_L g829 ( .A(n_120), .Y(n_829) );
NOR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_397), .Y(n_120) );
NAND4xp75_ASAP7_75t_L g121 ( .A(n_122), .B(n_302), .C(n_344), .D(n_368), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_191), .B(n_239), .C(n_281), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g388 ( .A(n_126), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g482 ( .A(n_126), .B(n_419), .Y(n_482) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_152), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g297 ( .A(n_128), .B(n_249), .Y(n_297) );
AND2x2_ASAP7_75t_L g338 ( .A(n_128), .B(n_299), .Y(n_338) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g245 ( .A(n_129), .B(n_174), .Y(n_245) );
OR2x2_ASAP7_75t_L g263 ( .A(n_129), .B(n_174), .Y(n_263) );
INVx2_ASAP7_75t_L g289 ( .A(n_129), .Y(n_289) );
AND2x2_ASAP7_75t_L g319 ( .A(n_129), .B(n_249), .Y(n_319) );
AND2x2_ASAP7_75t_L g348 ( .A(n_129), .B(n_173), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_129), .B(n_300), .Y(n_384) );
AO31x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_142), .A3(n_146), .B(n_149), .Y(n_129) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B1(n_138), .B2(n_140), .Y(n_130) );
INVx4_ASAP7_75t_L g134 ( .A(n_132), .Y(n_134) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_133), .Y(n_204) );
INVx2_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_134), .A2(n_253), .B(n_254), .C(n_255), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_135), .A2(n_156), .B1(n_219), .B2(n_220), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_135), .A2(n_140), .B1(n_272), .B2(n_274), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_135), .A2(n_136), .B1(n_497), .B2(n_498), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_135), .A2(n_530), .B1(n_532), .B2(n_533), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_135), .A2(n_156), .B1(n_555), .B2(n_557), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_135), .A2(n_575), .B(n_576), .Y(n_574) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_136), .B(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_136), .A2(n_258), .B(n_259), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_136), .A2(n_155), .B(n_165), .C(n_171), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_136), .A2(n_506), .B(n_507), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_136), .A2(n_206), .B1(n_564), .B2(n_565), .Y(n_563) );
BUFx8_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g141 ( .A(n_137), .Y(n_141) );
INVx2_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
INVx1_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_139), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g275 ( .A(n_139), .Y(n_275) );
INVx2_ASAP7_75t_L g509 ( .A(n_139), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_140), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_SL g532 ( .A(n_141), .Y(n_532) );
INVx1_ASAP7_75t_L g547 ( .A(n_141), .Y(n_547) );
INVx2_ASAP7_75t_L g503 ( .A(n_142), .Y(n_503) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
OAI21xp33_ASAP7_75t_L g171 ( .A1(n_143), .A2(n_163), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
INVx2_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
BUFx10_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
BUFx10_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
INVx1_ASAP7_75t_L g278 ( .A(n_147), .Y(n_278) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_147), .A2(n_528), .A3(n_554), .B(n_558), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx2_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
BUFx2_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_151), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_151), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_151), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g361 ( .A(n_152), .B(n_290), .Y(n_361) );
INVx2_ASAP7_75t_L g456 ( .A(n_152), .Y(n_456) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_173), .Y(n_152) );
INVx2_ASAP7_75t_L g244 ( .A(n_153), .Y(n_244) );
AND2x4_ASAP7_75t_L g287 ( .A(n_153), .B(n_174), .Y(n_287) );
AOI21x1_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_164), .B(n_170), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_163), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_156), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_156), .A2(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_162), .B(n_181), .Y(n_180) );
INVxp67_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
INVx3_ASAP7_75t_L g577 ( .A(n_167), .Y(n_577) );
OAI21xp33_ASAP7_75t_SL g230 ( .A1(n_168), .A2(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_169), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_172), .A2(n_199), .B(n_208), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_172), .A2(n_543), .B(n_548), .Y(n_542) );
AND2x2_ASAP7_75t_L g446 ( .A(n_173), .B(n_244), .Y(n_446) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g310 ( .A(n_174), .Y(n_310) );
AND2x2_ASAP7_75t_L g367 ( .A(n_174), .B(n_249), .Y(n_367) );
AND2x2_ASAP7_75t_L g382 ( .A(n_174), .B(n_290), .Y(n_382) );
AND2x2_ASAP7_75t_L g404 ( .A(n_174), .B(n_244), .Y(n_404) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_189), .Y(n_174) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_175), .A2(n_542), .B(n_551), .Y(n_541) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_188), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_183) );
INVx2_ASAP7_75t_L g273 ( .A(n_185), .Y(n_273) );
INVx1_ASAP7_75t_L g524 ( .A(n_186), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_186), .A2(n_202), .B1(n_545), .B2(n_546), .Y(n_544) );
OAI211xp5_ASAP7_75t_SL g451 ( .A1(n_191), .A2(n_452), .B(n_454), .C(n_461), .Y(n_451) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_225), .Y(n_192) );
INVxp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g438 ( .A(n_194), .B(n_374), .Y(n_438) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_215), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_195), .B(n_227), .Y(n_337) );
INVxp67_ASAP7_75t_L g351 ( .A(n_195), .Y(n_351) );
AND2x2_ASAP7_75t_L g371 ( .A(n_195), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_195), .B(n_284), .Y(n_378) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
AOI21x1_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_212), .Y(n_196) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_197), .A2(n_271), .A3(n_277), .B(n_279), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_203), .B(n_206), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
INVx2_ASAP7_75t_L g556 ( .A(n_202), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g276 ( .A(n_204), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g519 ( .A1(n_206), .A2(n_276), .B(n_520), .C(n_521), .Y(n_519) );
BUFx4f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_207), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g511 ( .A(n_207), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_SL g531 ( .A(n_211), .Y(n_531) );
INVx2_ASAP7_75t_L g221 ( .A(n_213), .Y(n_221) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_213), .B(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g238 ( .A(n_214), .B(n_222), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_214), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g517 ( .A(n_214), .Y(n_517) );
BUFx3_ASAP7_75t_L g528 ( .A(n_214), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_214), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g569 ( .A(n_214), .Y(n_569) );
OR2x2_ASAP7_75t_L g312 ( .A(n_215), .B(n_294), .Y(n_312) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g360 ( .A(n_216), .B(n_267), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_216), .B(n_270), .Y(n_366) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g266 ( .A(n_217), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g335 ( .A(n_217), .B(n_270), .Y(n_335) );
BUFx2_ASAP7_75t_L g342 ( .A(n_217), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_217), .B(n_270), .Y(n_422) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_221), .A3(n_222), .B(n_223), .Y(n_217) );
AOI31xp67_ASAP7_75t_L g495 ( .A1(n_221), .A2(n_222), .A3(n_496), .B(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_222), .A2(n_505), .B(n_508), .Y(n_504) );
OAI21x1_ASAP7_75t_L g518 ( .A1(n_222), .A2(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g352 ( .A(n_226), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g481 ( .A(n_226), .B(n_266), .Y(n_481) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g284 ( .A(n_227), .Y(n_284) );
AND2x2_ASAP7_75t_L g295 ( .A(n_227), .B(n_270), .Y(n_295) );
AND2x2_ASAP7_75t_L g341 ( .A(n_227), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g374 ( .A(n_227), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_227), .B(n_285), .Y(n_391) );
AND2x2_ASAP7_75t_L g430 ( .A(n_227), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_235), .B(n_238), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_246), .B(n_264), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_241), .A2(n_409), .B1(n_410), .B2(n_412), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_245), .Y(n_241) );
AND2x2_ASAP7_75t_L g406 ( .A(n_242), .B(n_297), .Y(n_406) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g470 ( .A(n_244), .B(n_290), .Y(n_470) );
AND2x2_ASAP7_75t_L g434 ( .A(n_245), .B(n_329), .Y(n_434) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_262), .Y(n_246) );
OR2x2_ASAP7_75t_L g331 ( .A(n_247), .B(n_308), .Y(n_331) );
OR2x2_ASAP7_75t_L g443 ( .A(n_247), .B(n_263), .Y(n_443) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g306 ( .A(n_248), .Y(n_306) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g290 ( .A(n_249), .Y(n_290) );
BUFx3_ASAP7_75t_L g372 ( .A(n_249), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_257), .B(n_260), .Y(n_251) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_256), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_522) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g440 ( .A(n_263), .B(n_299), .Y(n_440) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x2_ASAP7_75t_L g282 ( .A(n_266), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g323 ( .A(n_266), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g460 ( .A(n_266), .Y(n_460) );
INVx1_ASAP7_75t_L g479 ( .A(n_266), .Y(n_479) );
INVx2_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_267), .B(n_270), .Y(n_343) );
INVx1_ASAP7_75t_L g407 ( .A(n_268), .Y(n_407) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g468 ( .A(n_269), .Y(n_468) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
INVx1_ASAP7_75t_L g375 ( .A(n_270), .Y(n_375) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_277), .A2(n_528), .A3(n_529), .B(n_534), .Y(n_527) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_SL g566 ( .A(n_278), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_286), .B1(n_291), .B2(n_296), .Y(n_281) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
AND2x2_ASAP7_75t_L g326 ( .A(n_284), .B(n_311), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_284), .B(n_294), .Y(n_386) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx3_ASAP7_75t_L g317 ( .A(n_287), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_287), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g411 ( .A(n_287), .B(n_395), .Y(n_411) );
INVx1_ASAP7_75t_L g315 ( .A(n_288), .Y(n_315) );
AOI222xp33_ASAP7_75t_L g325 ( .A1(n_288), .A2(n_326), .B1(n_327), .B2(n_332), .C1(n_338), .C2(n_339), .Y(n_325) );
OAI21xp33_ASAP7_75t_SL g355 ( .A1(n_288), .A2(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g379 ( .A(n_288), .B(n_298), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_288), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OR2x2_ASAP7_75t_L g308 ( .A(n_289), .B(n_300), .Y(n_308) );
INVx1_ASAP7_75t_L g396 ( .A(n_289), .Y(n_396) );
BUFx2_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_293), .B(n_334), .Y(n_363) );
OR2x2_ASAP7_75t_L g475 ( .A(n_293), .B(n_335), .Y(n_475) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g358 ( .A(n_295), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g473 ( .A(n_295), .Y(n_473) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_296), .A2(n_455), .A3(n_457), .B(n_458), .Y(n_454) );
AND2x4_ASAP7_75t_SL g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_297), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_325), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_311), .B(n_313), .Y(n_303) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x6_ASAP7_75t_L g424 ( .A(n_306), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g356 ( .A(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g447 ( .A(n_310), .B(n_384), .Y(n_447) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_312), .A2(n_401), .B1(n_403), .B2(n_405), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_312), .A2(n_373), .B(n_435), .C(n_462), .Y(n_461) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B(n_322), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_317), .B(n_415), .C(n_416), .D(n_418), .Y(n_414) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_319), .B(n_321), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_319), .B(n_404), .Y(n_427) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g393 ( .A(n_324), .B(n_353), .Y(n_393) );
NAND2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_331), .A2(n_475), .B1(n_476), .B2(n_478), .Y(n_474) );
AOI221x1_ASAP7_75t_L g413 ( .A1(n_332), .A2(n_414), .B1(n_420), .B2(n_423), .C(n_426), .Y(n_413) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g353 ( .A(n_335), .Y(n_353) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g365 ( .A(n_337), .B(n_366), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_338), .B(n_419), .Y(n_428) );
O2A1O1Ixp5_ASAP7_75t_L g441 ( .A1(n_339), .A2(n_423), .B(n_442), .C(n_444), .Y(n_441) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx2_ASAP7_75t_L g390 ( .A(n_342), .Y(n_390) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_354), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_346), .A2(n_364), .B1(n_434), .B2(n_435), .C(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g370 ( .A(n_348), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_348), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g469 ( .A(n_348), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2x1_ASAP7_75t_L g448 ( .A(n_351), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g472 ( .A(n_351), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g412 ( .A(n_352), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_361), .B2(n_362), .C1(n_364), .C2(n_367), .Y(n_354) );
INVx1_ASAP7_75t_L g439 ( .A(n_358), .Y(n_439) );
INVx1_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g436 ( .A(n_360), .Y(n_436) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g377 ( .A(n_366), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g431 ( .A(n_366), .Y(n_431) );
AND2x2_ASAP7_75t_L g394 ( .A(n_367), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_387), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B1(n_376), .B2(n_379), .C1(n_380), .C2(n_385), .Y(n_369) );
INVx3_ASAP7_75t_L g419 ( .A(n_372), .Y(n_419) );
BUFx2_ASAP7_75t_L g477 ( .A(n_372), .Y(n_477) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g449 ( .A(n_374), .Y(n_449) );
OR2x2_ASAP7_75t_L g459 ( .A(n_374), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx2_ASAP7_75t_SL g417 ( .A(n_382), .Y(n_417) );
AND2x2_ASAP7_75t_L g462 ( .A(n_383), .B(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_384), .Y(n_415) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g421 ( .A(n_386), .B(n_422), .Y(n_421) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_388), .B(n_392), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
OR2x2_ASAP7_75t_L g478 ( .A(n_391), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g409 ( .A(n_393), .Y(n_409) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g416 ( .A(n_396), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g466 ( .A(n_396), .Y(n_466) );
NAND4xp75_ASAP7_75t_L g397 ( .A(n_398), .B(n_432), .C(n_450), .D(n_463), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_413), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_407), .B(n_408), .Y(n_399) );
INVxp33_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_402), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g425 ( .A(n_404), .Y(n_425) );
AND2x2_ASAP7_75t_L g465 ( .A(n_404), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g435 ( .A(n_407), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp33_ASAP7_75t_SL g444 ( .A1(n_421), .A2(n_445), .B1(n_447), .B2(n_448), .Y(n_444) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_428), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g457 ( .A(n_428), .Y(n_457) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_441), .Y(n_432) );
AOI21xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_439), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_480), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B1(n_469), .B2(n_471), .C(n_474), .Y(n_464) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx4_ASAP7_75t_L g821 ( .A(n_483), .Y(n_821) );
BUFx12f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g840 ( .A(n_485), .B(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g850 ( .A(n_486), .Y(n_850) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_722), .Y(n_487) );
AND4x1_ASAP7_75t_L g488 ( .A(n_489), .B(n_644), .C(n_677), .D(n_708), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_611), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_536), .B1(n_579), .B2(n_589), .C(n_598), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_491), .A2(n_701), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_514), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
INVx2_ASAP7_75t_L g597 ( .A(n_494), .Y(n_597) );
AND2x2_ASAP7_75t_L g607 ( .A(n_494), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g643 ( .A(n_494), .B(n_527), .Y(n_643) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g632 ( .A(n_495), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g618 ( .A(n_502), .B(n_608), .Y(n_618) );
OR2x2_ASAP7_75t_L g727 ( .A(n_502), .B(n_516), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_513), .Y(n_502) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_503), .A2(n_504), .B(n_513), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_512), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_514), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_527), .Y(n_515) );
INVx1_ASAP7_75t_L g592 ( .A(n_516), .Y(n_592) );
INVx2_ASAP7_75t_SL g669 ( .A(n_516), .Y(n_669) );
BUFx2_ASAP7_75t_L g699 ( .A(n_516), .Y(n_699) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_526), .Y(n_516) );
OA21x2_ASAP7_75t_L g608 ( .A1(n_517), .A2(n_518), .B(n_526), .Y(n_608) );
AND2x2_ASAP7_75t_L g591 ( .A(n_527), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g610 ( .A(n_527), .Y(n_610) );
OR2x2_ASAP7_75t_L g630 ( .A(n_527), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g671 ( .A(n_527), .Y(n_671) );
INVx1_ASAP7_75t_L g682 ( .A(n_527), .Y(n_682) );
AND2x2_ASAP7_75t_L g689 ( .A(n_527), .B(n_631), .Y(n_689) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_538), .B(n_560), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_552), .Y(n_538) );
INVx1_ASAP7_75t_L g603 ( .A(n_539), .Y(n_603) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_540), .Y(n_615) );
INVx1_ASAP7_75t_L g624 ( .A(n_540), .Y(n_624) );
INVx1_ASAP7_75t_L g663 ( .A(n_540), .Y(n_663) );
AND2x2_ASAP7_75t_L g693 ( .A(n_540), .B(n_553), .Y(n_693) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g587 ( .A(n_541), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g599 ( .A(n_552), .Y(n_599) );
AND2x4_ASAP7_75t_L g648 ( .A(n_552), .B(n_562), .Y(n_648) );
AND2x2_ASAP7_75t_L g658 ( .A(n_552), .B(n_587), .Y(n_658) );
INVx1_ASAP7_75t_L g719 ( .A(n_552), .Y(n_719) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g605 ( .A(n_553), .B(n_584), .Y(n_605) );
AND2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g639 ( .A(n_553), .B(n_584), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_553), .B(n_567), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_560), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .Y(n_560) );
OR2x2_ASAP7_75t_L g765 ( .A(n_561), .B(n_567), .Y(n_765) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g712 ( .A(n_562), .Y(n_712) );
AND2x2_ASAP7_75t_L g737 ( .A(n_562), .B(n_567), .Y(n_737) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_566), .A2(n_571), .B(n_574), .Y(n_570) );
INVx3_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
AND2x2_ASAP7_75t_L g614 ( .A(n_567), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
INVx1_ASAP7_75t_L g650 ( .A(n_567), .Y(n_650) );
INVx1_ASAP7_75t_L g660 ( .A(n_567), .Y(n_660) );
BUFx2_ASAP7_75t_L g755 ( .A(n_567), .Y(n_755) );
OR2x2_ASAP7_75t_L g783 ( .A(n_567), .B(n_587), .Y(n_783) );
INVxp67_ASAP7_75t_L g800 ( .A(n_567), .Y(n_800) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_578), .Y(n_568) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_585), .Y(n_580) );
AND2x4_ASAP7_75t_L g613 ( .A(n_581), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_581), .B(n_693), .Y(n_774) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g601 ( .A(n_583), .B(n_588), .Y(n_601) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
INVx1_ASAP7_75t_L g749 ( .A(n_583), .Y(n_749) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g662 ( .A(n_584), .Y(n_662) );
AND2x2_ASAP7_75t_L g676 ( .A(n_585), .B(n_639), .Y(n_676) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
OR2x2_ASAP7_75t_L g696 ( .A(n_587), .B(n_662), .Y(n_696) );
INVx1_ASAP7_75t_L g759 ( .A(n_587), .Y(n_759) );
AND2x2_ASAP7_75t_L g702 ( .A(n_588), .B(n_648), .Y(n_702) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
AND2x2_ASAP7_75t_L g705 ( .A(n_591), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
AND2x2_ASAP7_75t_L g609 ( .A(n_594), .B(n_610), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_594), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g628 ( .A(n_595), .Y(n_628) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g707 ( .A(n_596), .B(n_632), .Y(n_707) );
AND2x2_ASAP7_75t_L g670 ( .A(n_597), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g741 ( .A(n_597), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_602), .C(n_606), .Y(n_598) );
INVx1_ASAP7_75t_L g733 ( .A(n_600), .Y(n_733) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g729 ( .A(n_601), .B(n_693), .Y(n_729) );
INVx1_ASAP7_75t_L g820 ( .A(n_601), .Y(n_820) );
INVx1_ASAP7_75t_L g785 ( .A(n_602), .Y(n_785) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g818 ( .A(n_603), .B(n_737), .Y(n_818) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g635 ( .A(n_605), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g790 ( .A(n_605), .B(n_755), .Y(n_790) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVxp67_ASAP7_75t_L g680 ( .A(n_607), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_607), .B(n_642), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_607), .B(n_609), .Y(n_772) );
INVx1_ASAP7_75t_L g655 ( .A(n_608), .Y(n_655) );
INVx2_ASAP7_75t_SL g620 ( .A(n_610), .Y(n_620) );
OR2x2_ASAP7_75t_L g649 ( .A(n_610), .B(n_650), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_616), .B1(n_621), .B2(n_626), .C(n_633), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_SL g657 ( .A(n_613), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g685 ( .A(n_615), .Y(n_685) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g742 ( .A(n_618), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_618), .B(n_620), .Y(n_780) );
OR2x2_ASAP7_75t_L g762 ( .A(n_619), .B(n_752), .Y(n_762) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g731 ( .A(n_620), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g778 ( .A(n_620), .B(n_707), .Y(n_778) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g713 ( .A(n_623), .B(n_636), .Y(n_713) );
BUFx2_ASAP7_75t_L g739 ( .A(n_623), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_627), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g642 ( .A(n_628), .Y(n_642) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g715 ( .A(n_630), .Y(n_715) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B(n_640), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g692 ( .A(n_636), .Y(n_692) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_636), .Y(n_695) );
OR2x2_ASAP7_75t_L g805 ( .A(n_636), .B(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g766 ( .A(n_637), .Y(n_766) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
AND2x2_ASAP7_75t_L g801 ( .A(n_639), .B(n_674), .Y(n_801) );
INVx2_ASAP7_75t_SL g806 ( .A(n_639), .Y(n_806) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx2_ASAP7_75t_L g688 ( .A(n_642), .Y(n_688) );
AND2x4_ASAP7_75t_L g664 ( .A(n_643), .B(n_653), .Y(n_664) );
INVx2_ASAP7_75t_L g728 ( .A(n_643), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_643), .B(n_669), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_643), .B(n_699), .Y(n_815) );
AOI221x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_651), .B1(n_656), .B2(n_664), .C(n_665), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx2_ASAP7_75t_L g784 ( .A(n_647), .Y(n_784) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_647), .A2(n_792), .B(n_794), .Y(n_791) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g673 ( .A(n_648), .B(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g704 ( .A(n_648), .Y(n_704) );
AND2x4_ASAP7_75t_L g758 ( .A(n_648), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g718 ( .A(n_650), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g763 ( .A1(n_652), .A2(n_761), .A3(n_764), .B1(n_766), .B2(n_767), .Y(n_763) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_653), .B(n_670), .Y(n_786) );
AND2x2_ASAP7_75t_L g802 ( .A(n_653), .B(n_682), .Y(n_802) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_657), .B(n_659), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_658), .B(n_800), .Y(n_799) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_659), .A2(n_735), .B(n_738), .C(n_740), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g683 ( .A(n_661), .Y(n_683) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_672), .B(n_675), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_666), .A2(n_701), .B(n_703), .Y(n_700) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_669), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_673), .A2(n_746), .B1(n_750), .B2(n_751), .Y(n_745) );
AND2x2_ASAP7_75t_L g812 ( .A(n_673), .B(n_800), .Y(n_812) );
NOR2xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_700), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_683), .B1(n_684), .B2(n_686), .C(n_690), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g788 ( .A1(n_679), .A2(n_789), .B(n_790), .Y(n_788) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g771 ( .A(n_685), .B(n_737), .Y(n_771) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AOI31xp33_ASAP7_75t_L g708 ( .A1(n_688), .A2(n_709), .A3(n_714), .B(n_716), .Y(n_708) );
AND2x2_ASAP7_75t_L g808 ( .A(n_688), .B(n_715), .Y(n_808) );
AND2x2_ASAP7_75t_L g697 ( .A(n_689), .B(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_689), .Y(n_761) );
INVx1_ASAP7_75t_L g795 ( .A(n_689), .Y(n_795) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_694), .B(n_697), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx2_ASAP7_75t_L g721 ( .A(n_693), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_693), .B(n_820), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_694), .A2(n_777), .B(n_779), .Y(n_776) );
NOR2x1p5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_696), .A2(n_711), .B(n_718), .C(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g730 ( .A(n_699), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g750 ( .A(n_699), .B(n_706), .Y(n_750) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g732 ( .A(n_707), .Y(n_732) );
INVx1_ASAP7_75t_L g768 ( .A(n_707), .Y(n_768) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_713), .A2(n_730), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g789 ( .A(n_713), .Y(n_789) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_775), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_743), .C(n_753), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_729), .B1(n_730), .B2(n_733), .C(n_734), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_731), .A2(n_798), .B1(n_801), .B2(n_802), .Y(n_797) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
OR2x2_ASAP7_75t_L g794 ( .A(n_742), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g793 ( .A(n_748), .Y(n_793) );
INVx2_ASAP7_75t_L g773 ( .A(n_750), .Y(n_773) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI211xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B(n_763), .C(n_769), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_760), .B(n_762), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g764 ( .A(n_759), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g807 ( .A(n_764), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND4xp75_ASAP7_75t_L g775 ( .A(n_776), .B(n_787), .C(n_796), .D(n_809), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_785), .B2(n_786), .Y(n_779) );
NAND2x1_ASAP7_75t_SL g781 ( .A(n_782), .B(n_784), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_803), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B(n_808), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B1(n_813), .B2(n_816), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVxp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
A2O1A1O1Ixp25_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_828), .B(n_830), .C(n_832), .D(n_834), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
INVx4_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
INVx6_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
BUFx10_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx3_ASAP7_75t_L g855 ( .A(n_842), .Y(n_855) );
AND2x4_ASAP7_75t_L g842 ( .A(n_843), .B(n_847), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
NOR2x1p5_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
CKINVDCx14_ASAP7_75t_R g853 ( .A(n_854), .Y(n_853) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
endmodule