module fake_jpeg_220_n_675 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_675);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_675;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_19),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_60),
.B(n_61),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_62),
.Y(n_172)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_65),
.B(n_67),
.Y(n_161)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_71),
.Y(n_164)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_73),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_75),
.B(n_81),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_82),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_0),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_20),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_89),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g156 ( 
.A(n_92),
.Y(n_156)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_40),
.B(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_100),
.Y(n_158)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_3),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_104),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_105),
.Y(n_231)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_54),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_112),
.B(n_116),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_25),
.Y(n_114)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_54),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_117),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_37),
.Y(n_173)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx16f_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_45),
.B(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_123),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_3),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_130),
.B(n_73),
.Y(n_193)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_36),
.B(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_4),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_26),
.B1(n_52),
.B2(n_23),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_137),
.A2(n_140),
.B1(n_224),
.B2(n_225),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_84),
.A2(n_27),
.B1(n_48),
.B2(n_32),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_92),
.A2(n_31),
.B1(n_27),
.B2(n_48),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_141),
.A2(n_177),
.B1(n_181),
.B2(n_210),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_31),
.B1(n_23),
.B2(n_52),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_148),
.A2(n_141),
.B(n_181),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_21),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_152),
.B(n_154),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_101),
.B(n_21),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_32),
.B1(n_48),
.B2(n_53),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_157),
.A2(n_162),
.B1(n_168),
.B2(n_171),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_59),
.A2(n_56),
.B1(n_53),
.B2(n_46),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_90),
.A2(n_32),
.B1(n_46),
.B2(n_43),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_74),
.A2(n_56),
.B1(n_43),
.B2(n_37),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_68),
.A2(n_36),
.B1(n_26),
.B2(n_34),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_178),
.A2(n_205),
.B(n_15),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_120),
.A2(n_34),
.B1(n_25),
.B2(n_29),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_62),
.B(n_4),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_186),
.B(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_193),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_93),
.A2(n_34),
.B1(n_25),
.B2(n_29),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_189),
.A2(n_196),
.B1(n_201),
.B2(n_213),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_99),
.B(n_127),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_79),
.A2(n_34),
.B1(n_29),
.B2(n_7),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_117),
.B(n_5),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_197),
.B(n_199),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_5),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_88),
.A2(n_34),
.B1(n_7),
.B2(n_8),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_96),
.B(n_131),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_203),
.B(n_206),
.Y(n_286)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_214),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_110),
.A2(n_6),
.B(n_8),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_131),
.B(n_6),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_6),
.C(n_8),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_211),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_77),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_103),
.B(n_9),
.C(n_10),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_109),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_113),
.B(n_12),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_217),
.B(n_205),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_83),
.B(n_12),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_219),
.B(n_228),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_95),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_70),
.A2(n_13),
.B1(n_15),
.B2(n_78),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_115),
.B(n_13),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_107),
.B1(n_119),
.B2(n_111),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_232),
.A2(n_249),
.B1(n_255),
.B2(n_269),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_234),
.Y(n_351)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g342 ( 
.A(n_235),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_167),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_237),
.B(n_238),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_161),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_239),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_240),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_241),
.B(n_244),
.Y(n_343)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_173),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_245),
.B(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_140),
.A2(n_98),
.B1(n_105),
.B2(n_128),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_247),
.A2(n_254),
.B1(n_307),
.B2(n_293),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_172),
.A2(n_73),
.B1(n_118),
.B2(n_122),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

AO22x2_ASAP7_75t_L g254 ( 
.A1(n_195),
.A2(n_97),
.B1(n_64),
.B2(n_118),
.Y(n_254)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_254),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_172),
.A2(n_15),
.B1(n_97),
.B2(n_219),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_164),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_256),
.B(n_261),
.Y(n_359)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_166),
.Y(n_258)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_133),
.B(n_135),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_262),
.B(n_263),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_165),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_151),
.B(n_163),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_265),
.B(n_270),
.Y(n_373)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_266),
.Y(n_366)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_268),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_175),
.A2(n_146),
.B1(n_179),
.B2(n_176),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_169),
.B(n_145),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g272 ( 
.A(n_136),
.Y(n_272)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_194),
.Y(n_273)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_136),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_274),
.B(n_275),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_216),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_216),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_277),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_278),
.A2(n_300),
.B1(n_311),
.B2(n_314),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_158),
.B(n_143),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_280),
.Y(n_336)
);

OR2x4_ASAP7_75t_L g281 ( 
.A(n_177),
.B(n_210),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_281),
.A2(n_306),
.B(n_254),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_139),
.B(n_218),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_290),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_138),
.B(n_150),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_227),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_285),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_156),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_289),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_227),
.B(n_231),
.Y(n_290)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_146),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_291),
.A2(n_302),
.B1(n_304),
.B2(n_312),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_159),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_292),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_153),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_293),
.B(n_296),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_149),
.B(n_147),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g344 ( 
.A(n_294),
.B(n_316),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_171),
.B(n_231),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_153),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_195),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_149),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_298),
.Y(n_377)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_190),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_301),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_180),
.B(n_147),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_160),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_174),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_190),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_168),
.A2(n_157),
.B(n_192),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_215),
.B(n_202),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_308),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_196),
.A2(n_220),
.B(n_180),
.C(n_202),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_215),
.B(n_174),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_309),
.B(n_310),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_184),
.B(n_142),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_200),
.B(n_226),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_184),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_200),
.Y(n_313)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_182),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_142),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_315),
.A2(n_239),
.B1(n_240),
.B2(n_292),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_226),
.B(n_144),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_281),
.A2(n_144),
.B(n_182),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_324),
.A2(n_349),
.B(n_352),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_257),
.B1(n_295),
.B2(n_287),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_328),
.B1(n_329),
.B2(n_331),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_308),
.B1(n_286),
.B2(n_309),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_306),
.A2(n_233),
.B1(n_301),
.B2(n_310),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_297),
.B1(n_253),
.B2(n_277),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_332),
.A2(n_364),
.B1(n_276),
.B2(n_313),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_286),
.A2(n_279),
.B1(n_248),
.B2(n_303),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_334),
.A2(n_337),
.B1(n_347),
.B2(n_370),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_279),
.A2(n_248),
.B1(n_303),
.B2(n_251),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_278),
.A2(n_271),
.B1(n_251),
.B2(n_236),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_271),
.A2(n_254),
.B(n_294),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_271),
.A2(n_254),
.B(n_294),
.Y(n_352)
);

AOI32xp33_ASAP7_75t_L g353 ( 
.A1(n_256),
.A2(n_238),
.A3(n_241),
.B1(n_237),
.B2(n_263),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_353),
.A2(n_260),
.B(n_259),
.C(n_304),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_250),
.B(n_246),
.C(n_284),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_347),
.C(n_348),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_293),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_271),
.A2(n_275),
.B1(n_312),
.B2(n_302),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_315),
.A2(n_268),
.B1(n_252),
.B2(n_258),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_371),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_336),
.B(n_242),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_379),
.B(n_389),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_380),
.Y(n_442)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_266),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_387),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx8_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_296),
.Y(n_387)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_388),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_356),
.B(n_243),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_359),
.B(n_298),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_390),
.B(n_397),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_319),
.Y(n_391)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_392),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_362),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_394),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_413),
.C(n_387),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_334),
.B(n_267),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_356),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_398),
.B(n_409),
.Y(n_458)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_399),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_419),
.B(n_422),
.Y(n_432)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_325),
.A2(n_264),
.B1(n_299),
.B2(n_273),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_402),
.A2(n_404),
.B1(n_420),
.B2(n_332),
.Y(n_437)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_403),
.Y(n_455)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_405),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_327),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_410),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_235),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_365),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_289),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_291),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_412),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_337),
.B(n_343),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_416),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_338),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_417),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_328),
.A2(n_364),
.B1(n_324),
.B2(n_352),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_418),
.A2(n_344),
.B1(n_330),
.B2(n_317),
.Y(n_462)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_375),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_373),
.B(n_355),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_344),
.Y(n_441)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_318),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_423),
.A2(n_424),
.B(n_426),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_351),
.B(n_348),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

OA22x2_ASAP7_75t_L g445 ( 
.A1(n_425),
.A2(n_339),
.B1(n_360),
.B2(n_370),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_321),
.B(n_317),
.Y(n_426)
);

NOR2x1p5_ASAP7_75t_SL g436 ( 
.A(n_382),
.B(n_386),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_417),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_404),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_390),
.Y(n_478)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_445),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_450),
.C(n_468),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_367),
.B(n_349),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_449),
.A2(n_454),
.B(n_457),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_396),
.B(n_321),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_427),
.A2(n_367),
.B(n_361),
.Y(n_454)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_400),
.A2(n_339),
.B(n_338),
.C(n_333),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_456),
.A2(n_397),
.B(n_380),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_380),
.A2(n_317),
.B(n_333),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_467),
.B1(n_383),
.B2(n_423),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_384),
.B(n_344),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_465),
.B(n_419),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_418),
.A2(n_326),
.B1(n_358),
.B2(n_378),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_415),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_484),
.Y(n_509)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_394),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_477),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_475),
.A2(n_507),
.B(n_508),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_476),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_453),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_488),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_436),
.B(n_393),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_479),
.B(n_485),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g480 ( 
.A1(n_467),
.A2(n_383),
.B1(n_402),
.B2(n_407),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_480),
.A2(n_491),
.B1(n_500),
.B2(n_503),
.Y(n_518)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_482),
.A2(n_452),
.B1(n_440),
.B2(n_444),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_392),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_381),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_457),
.Y(n_512)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_410),
.C(n_326),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_492),
.C(n_496),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_434),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_490),
.B(n_495),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_395),
.C(n_399),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_433),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_493),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_430),
.B(n_388),
.Y(n_494)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_494),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_439),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_401),
.C(n_405),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_497),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_430),
.B(n_422),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_499),
.A2(n_501),
.B(n_502),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_439),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_429),
.B(n_428),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_416),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_432),
.A2(n_358),
.B1(n_403),
.B2(n_385),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_466),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_505),
.A2(n_431),
.B1(n_481),
.B2(n_487),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_438),
.B(n_425),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_L g517 ( 
.A1(n_506),
.A2(n_456),
.B(n_446),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_462),
.A2(n_391),
.B1(n_385),
.B2(n_414),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_442),
.A2(n_378),
.B(n_377),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_512),
.B(n_523),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_468),
.C(n_435),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_515),
.B(n_525),
.C(n_528),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_517),
.A2(n_479),
.B(n_485),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_498),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_519),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_498),
.A2(n_432),
.B1(n_437),
.B2(n_458),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_507),
.Y(n_563)
);

XNOR2x1_ASAP7_75t_L g523 ( 
.A(n_489),
.B(n_442),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_483),
.B(n_435),
.C(n_446),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_486),
.B(n_461),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_526),
.B(n_536),
.Y(n_567)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_527),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_492),
.B(n_496),
.C(n_488),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_440),
.C(n_461),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_538),
.C(n_540),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_534),
.A2(n_506),
.B(n_473),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_482),
.A2(n_452),
.B1(n_469),
.B2(n_445),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_535),
.A2(n_543),
.B1(n_503),
.B2(n_482),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_469),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_452),
.C(n_443),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_484),
.B(n_377),
.C(n_433),
.Y(n_540)
);

XNOR2x1_ASAP7_75t_L g542 ( 
.A(n_475),
.B(n_445),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_542),
.B(n_532),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_474),
.A2(n_445),
.B1(n_455),
.B2(n_463),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_476),
.B(n_376),
.C(n_369),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_544),
.B(n_508),
.C(n_505),
.Y(n_554)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_511),
.Y(n_546)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_546),
.Y(n_597)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_516),
.Y(n_548)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_548),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_497),
.Y(n_550)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_550),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_SL g584 ( 
.A(n_552),
.B(n_536),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_557),
.C(n_559),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_513),
.B(n_491),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_513),
.B(n_525),
.C(n_528),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_558),
.A2(n_563),
.B1(n_529),
.B2(n_571),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_515),
.B(n_494),
.C(n_493),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_523),
.B(n_470),
.C(n_499),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_560),
.B(n_566),
.C(n_544),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_531),
.B(n_502),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_564),
.Y(n_583)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_562),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_512),
.B(n_472),
.C(n_471),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_534),
.A2(n_535),
.B1(n_514),
.B2(n_519),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_568),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_520),
.B(n_351),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_569),
.B(n_572),
.Y(n_591)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_570),
.B(n_571),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_510),
.B(n_455),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_526),
.B(n_350),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_530),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_570),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_532),
.A2(n_463),
.B(n_368),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_575),
.Y(n_594)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_541),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_517),
.B(n_414),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_576),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_563),
.A2(n_518),
.B1(n_551),
.B2(n_547),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_577),
.A2(n_586),
.B1(n_537),
.B2(n_542),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_567),
.B(n_545),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_578),
.B(n_584),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_581),
.B(n_408),
.Y(n_614)
);

FAx1_ASAP7_75t_SL g587 ( 
.A(n_560),
.B(n_509),
.CI(n_524),
.CON(n_587),
.SN(n_587)
);

FAx1_ASAP7_75t_SL g610 ( 
.A(n_587),
.B(n_545),
.CI(n_540),
.CON(n_610),
.SN(n_610)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_557),
.B(n_549),
.C(n_555),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_588),
.B(n_592),
.Y(n_604)
);

A2O1A1O1Ixp25_ASAP7_75t_L g590 ( 
.A1(n_566),
.A2(n_509),
.B(n_559),
.C(n_553),
.D(n_529),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_590),
.A2(n_556),
.B(n_572),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_549),
.B(n_553),
.C(n_567),
.Y(n_592)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_593),
.Y(n_616)
);

INVx13_ASAP7_75t_L g598 ( 
.A(n_565),
.Y(n_598)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_598),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_538),
.C(n_554),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_573),
.C(n_546),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_594),
.Y(n_603)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_603),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_605),
.A2(n_608),
.B(n_618),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_552),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_614),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_590),
.A2(n_574),
.B(n_564),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_609),
.B(n_622),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_610),
.B(n_611),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_586),
.A2(n_562),
.B1(n_533),
.B2(n_459),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_613),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_600),
.B(n_451),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_578),
.B(n_601),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_615),
.B(n_619),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_408),
.C(n_376),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_617),
.B(n_620),
.C(n_585),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_SL g618 ( 
.A1(n_596),
.A2(n_451),
.B(n_459),
.C(n_368),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_577),
.B(n_369),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_579),
.B(n_320),
.C(n_354),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_579),
.B(n_323),
.Y(n_621)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_621),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_323),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_625),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_603),
.B(n_583),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_604),
.B(n_580),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_628),
.B(n_631),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_616),
.A2(n_580),
.B1(n_595),
.B2(n_582),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_592),
.C(n_596),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_632),
.B(n_633),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_617),
.B(n_584),
.C(n_591),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_611),
.B(n_582),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_634),
.B(n_602),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_606),
.B(n_587),
.C(n_593),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_636),
.B(n_637),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_587),
.C(n_589),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_623),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_640),
.B(n_643),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_639),
.A2(n_612),
.B(n_619),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_641),
.A2(n_650),
.B(n_629),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_635),
.B(n_607),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_638),
.B(n_597),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_646),
.B(n_647),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_636),
.B(n_615),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_630),
.A2(n_589),
.B1(n_618),
.B2(n_610),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_648),
.B(n_627),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_637),
.A2(n_610),
.B(n_618),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_634),
.A2(n_618),
.B1(n_602),
.B2(n_598),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_651),
.A2(n_319),
.B1(n_354),
.B2(n_340),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_652),
.B(n_632),
.Y(n_656)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_653),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_655),
.A2(n_658),
.B(n_659),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_656),
.B(n_657),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_642),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_644),
.A2(n_633),
.B(n_624),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_645),
.B(n_626),
.C(n_629),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g667 ( 
.A(n_660),
.B(n_651),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_652),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_665),
.A2(n_666),
.B(n_667),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_661),
.A2(n_649),
.B(n_650),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_663),
.A2(n_654),
.B(n_641),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_669),
.A2(n_670),
.B(n_662),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_664),
.A2(n_340),
.B(n_350),
.Y(n_670)
);

BUFx24_ASAP7_75t_SL g673 ( 
.A(n_671),
.Y(n_673)
);

AOI321xp33_ASAP7_75t_SL g672 ( 
.A1(n_668),
.A2(n_342),
.A3(n_357),
.B1(n_665),
.B2(n_667),
.C(n_669),
.Y(n_672)
);

FAx1_ASAP7_75t_SL g674 ( 
.A(n_673),
.B(n_672),
.CI(n_357),
.CON(n_674),
.SN(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_342),
.Y(n_675)
);


endmodule