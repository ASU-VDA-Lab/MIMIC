module real_jpeg_28852_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_329, n_5, n_4, n_1, n_328, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_329;
input n_5;
input n_4;
input n_1;
input n_328;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_29),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_2),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_2),
.A2(n_39),
.B1(n_58),
.B2(n_60),
.Y(n_321)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_44),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_29),
.B1(n_33),
.B2(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_4),
.A2(n_53),
.B1(n_65),
.B2(n_66),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_4),
.A2(n_53),
.B1(n_58),
.B2(n_60),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_58),
.B1(n_60),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_89),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_5),
.A2(n_44),
.B1(n_46),
.B2(n_89),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_5),
.A2(n_29),
.B1(n_33),
.B2(n_89),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_6),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_62),
.B(n_66),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_58),
.B1(n_60),
.B2(n_94),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_6),
.B(n_64),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_6),
.A2(n_46),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_46),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_83),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_6),
.A2(n_27),
.B1(n_220),
.B2(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_6),
.A2(n_65),
.B(n_236),
.Y(n_235)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_81),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_8),
.A2(n_44),
.B1(n_46),
.B2(n_81),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_8),
.A2(n_29),
.B1(n_33),
.B2(n_81),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_9),
.A2(n_34),
.B1(n_44),
.B2(n_46),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_34),
.B1(n_65),
.B2(n_66),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_9),
.A2(n_34),
.B1(n_58),
.B2(n_60),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_10),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_44),
.B1(n_46),
.B2(n_57),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_57),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_29),
.B1(n_33),
.B2(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_58),
.B1(n_60),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_12),
.A2(n_29),
.B1(n_33),
.B2(n_70),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_12),
.A2(n_44),
.B1(n_46),
.B2(n_70),
.Y(n_240)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_15),
.A2(n_29),
.B1(n_33),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_15),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_15),
.A2(n_44),
.B1(n_46),
.B2(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_104),
.Y(n_301)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_17),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_17),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_17),
.A2(n_43),
.B1(n_58),
.B2(n_60),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_17),
.A2(n_29),
.B1(n_33),
.B2(n_43),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_309),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_278),
.A3(n_305),
.B1(n_307),
.B2(n_308),
.C(n_328),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_126),
.A3(n_149),
.B1(n_272),
.B2(n_277),
.C(n_329),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_22),
.A2(n_273),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_107),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_23),
.B(n_107),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_84),
.C(n_101),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_24),
.B(n_101),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_25),
.B(n_55),
.C(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_26),
.B(n_40),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_27),
.A2(n_35),
.B1(n_38),
.B2(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_27),
.A2(n_35),
.B(n_103),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_27),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_27),
.A2(n_37),
.B1(n_214),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_27),
.A2(n_208),
.B1(n_209),
.B2(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_28),
.A2(n_32),
.B1(n_36),
.B2(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_28),
.A2(n_36),
.B1(n_97),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_28),
.A2(n_36),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_29),
.B(n_49),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_29),
.B(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_33),
.A2(n_46),
.A3(n_51),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g209 ( 
.A(n_36),
.Y(n_209)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_37),
.B(n_94),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_42),
.A2(n_113),
.B1(n_116),
.B2(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_46),
.B1(n_75),
.B2(n_78),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_44),
.A2(n_65),
.A3(n_78),
.B1(n_237),
.B2(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_46),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_47),
.A2(n_48),
.B1(n_115),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_47),
.A2(n_48),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_47),
.A2(n_48),
.B1(n_194),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_47),
.A2(n_48),
.B1(n_161),
.B2(n_262),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_47),
.A2(n_48),
.B(n_136),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_48),
.B(n_94),
.Y(n_221)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_71),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_61),
.B1(n_64),
.B2(n_69),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_68),
.B(n_94),
.C(n_95),
.Y(n_93)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_61),
.A2(n_64),
.B1(n_69),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_61),
.A2(n_64),
.B1(n_88),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_61),
.A2(n_64),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_74),
.B(n_76),
.C(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_74),
.Y(n_76)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_66),
.B(n_94),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_82),
.B1(n_83),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_72),
.A2(n_83),
.B1(n_157),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_72),
.A2(n_83),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_72),
.A2(n_83),
.B1(n_287),
.B2(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_77),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_73),
.A2(n_77),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_73),
.A2(n_77),
.B1(n_99),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_73),
.A2(n_77),
.B1(n_169),
.B2(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_73),
.A2(n_77),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_78),
.Y(n_246)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_84),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.C(n_98),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_85),
.B(n_98),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_90),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_86),
.A2(n_90),
.B1(n_143),
.B2(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_86),
.A2(n_90),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_92),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_96),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_125),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_119),
.C(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_113),
.A2(n_116),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_118),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_117),
.A2(n_141),
.B(n_144),
.Y(n_292)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_119),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_122),
.CI(n_124),
.CON(n_119),
.SN(n_119)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_122),
.C(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_127),
.B(n_128),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_147),
.B2(n_148),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_131),
.B(n_138),
.C(n_148),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_135),
.B(n_137),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_135),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_134),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_137),
.B(n_280),
.CI(n_292),
.CON(n_279),
.SN(n_279)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_147),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_179),
.C(n_184),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_173),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_151),
.B(n_173),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_164),
.C(n_165),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_152),
.B(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_159),
.C(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_164),
.Y(n_270)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_172),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_171),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_180),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_181),
.B(n_182),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_266),
.B(n_271),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_252),
.B(n_265),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_230),
.B(n_251),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_210),
.B(n_229),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_199),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_217),
.B(n_228),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_216),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_222),
.B(n_227),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_232),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_243),
.B1(n_249),
.B2(n_250),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_242),
.C(n_250),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_254),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_261),
.C(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_260),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_293),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_279),
.B(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_293),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_291),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_282),
.B1(n_295),
.B2(n_303),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_285),
.C(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_303),
.C(n_304),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_290),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_296),
.C(n_300),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_304),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_300),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_324),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);


endmodule