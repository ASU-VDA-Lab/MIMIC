module real_aes_130_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g224 ( .A(n_0), .B(n_139), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_1), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g130 ( .A(n_2), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_3), .B(n_123), .Y(n_122) );
NAND2xp33_ASAP7_75t_SL g209 ( .A(n_4), .B(n_129), .Y(n_209) );
INVx1_ASAP7_75t_L g200 ( .A(n_5), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_6), .B(n_143), .Y(n_474) );
INVx1_ASAP7_75t_L g517 ( .A(n_7), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g772 ( .A(n_8), .Y(n_772) );
AND2x2_ASAP7_75t_L g117 ( .A(n_9), .B(n_118), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_10), .Y(n_531) );
INVx2_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_12), .Y(n_424) );
INVx1_ASAP7_75t_L g482 ( .A(n_13), .Y(n_482) );
AOI221x1_ASAP7_75t_L g203 ( .A1(n_14), .A2(n_132), .B1(n_204), .B2(n_206), .C(n_208), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_15), .B(n_123), .Y(n_190) );
INVx1_ASAP7_75t_L g428 ( .A(n_16), .Y(n_428) );
INVx1_ASAP7_75t_L g480 ( .A(n_17), .Y(n_480) );
INVx1_ASAP7_75t_SL g467 ( .A(n_18), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_19), .B(n_124), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_20), .A2(n_132), .B(n_137), .Y(n_131) );
AOI221xp5_ASAP7_75t_SL g214 ( .A1(n_21), .A2(n_38), .B1(n_123), .B2(n_132), .C(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_22), .B(n_139), .Y(n_138) );
AOI33xp33_ASAP7_75t_L g497 ( .A1(n_23), .A2(n_52), .A3(n_176), .B1(n_183), .B2(n_498), .B3(n_499), .Y(n_497) );
AOI22x1_ASAP7_75t_R g755 ( .A1(n_24), .A2(n_36), .B1(n_756), .B2(n_757), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_24), .Y(n_757) );
INVx1_ASAP7_75t_L g525 ( .A(n_25), .Y(n_525) );
OR2x2_ASAP7_75t_L g120 ( .A(n_26), .B(n_92), .Y(n_120) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_26), .A2(n_92), .B(n_119), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_27), .B(n_141), .Y(n_194) );
INVxp67_ASAP7_75t_L g202 ( .A(n_28), .Y(n_202) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_29), .A2(n_105), .B1(n_765), .B2(n_776), .C1(n_796), .C2(n_798), .Y(n_104) );
AND2x2_ASAP7_75t_L g163 ( .A(n_29), .B(n_153), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g780 ( .A1(n_29), .A2(n_89), .B1(n_781), .B2(n_782), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_29), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_30), .B(n_174), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_31), .A2(n_132), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_32), .B(n_141), .Y(n_216) );
AND2x2_ASAP7_75t_L g129 ( .A(n_33), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g133 ( .A(n_33), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g182 ( .A(n_33), .Y(n_182) );
OR2x6_ASAP7_75t_L g426 ( .A(n_34), .B(n_427), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_35), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_36), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_37), .B(n_174), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_39), .A2(n_143), .B1(n_207), .B2(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_40), .B(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_41), .A2(n_82), .B1(n_132), .B2(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_42), .B(n_124), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_43), .B(n_139), .Y(n_161) );
XOR2xp5_ASAP7_75t_L g431 ( .A(n_44), .B(n_432), .Y(n_431) );
AOI22x1_ASAP7_75t_SL g788 ( .A1(n_44), .A2(n_67), .B1(n_789), .B2(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_44), .Y(n_789) );
XNOR2x2_ASAP7_75t_SL g754 ( .A(n_45), .B(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_46), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_47), .B(n_170), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_48), .B(n_124), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_49), .Y(n_444) );
AND2x2_ASAP7_75t_L g227 ( .A(n_50), .B(n_153), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_51), .B(n_153), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_53), .B(n_124), .Y(n_509) );
INVx1_ASAP7_75t_L g126 ( .A(n_54), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_54), .Y(n_136) );
AND2x2_ASAP7_75t_L g510 ( .A(n_55), .B(n_153), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_56), .A2(n_74), .B1(n_174), .B2(n_180), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_57), .B(n_174), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_58), .B(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_59), .B(n_207), .Y(n_533) );
AOI21xp5_ASAP7_75t_SL g454 ( .A1(n_60), .A2(n_180), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g154 ( .A(n_61), .B(n_153), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_62), .B(n_141), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_63), .B(n_139), .Y(n_150) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_64), .B(n_118), .Y(n_195) );
INVx1_ASAP7_75t_L g477 ( .A(n_65), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_66), .A2(n_132), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_67), .Y(n_790) );
INVx1_ASAP7_75t_L g508 ( .A(n_68), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_69), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_70), .B(n_170), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_71), .A2(n_180), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g134 ( .A(n_72), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_73), .B(n_174), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_75), .B(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g469 ( .A(n_76), .B(n_206), .Y(n_469) );
INVx1_ASAP7_75t_L g478 ( .A(n_77), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_78), .A2(n_180), .B(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_79), .A2(n_169), .B(n_180), .C(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_80), .B(n_123), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_81), .A2(n_85), .B1(n_123), .B2(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g429 ( .A(n_83), .Y(n_429) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_84), .B(n_206), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_86), .A2(n_180), .B1(n_495), .B2(n_496), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_87), .B(n_139), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_88), .B(n_139), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_89), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g753 ( .A(n_90), .B(n_754), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_91), .A2(n_132), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g456 ( .A(n_93), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_94), .B(n_141), .Y(n_149) );
AND2x2_ASAP7_75t_L g501 ( .A(n_95), .B(n_206), .Y(n_501) );
OAI22xp33_ASAP7_75t_SL g786 ( .A1(n_96), .A2(n_787), .B1(n_788), .B2(n_791), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_96), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_97), .A2(n_523), .B(n_524), .C(n_526), .Y(n_522) );
INVxp67_ASAP7_75t_L g205 ( .A(n_98), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_99), .B(n_123), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_100), .B(n_141), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_101), .A2(n_132), .B(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g773 ( .A(n_102), .Y(n_773) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_102), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_103), .B(n_124), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_753), .B(n_758), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OAI22x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_421), .B1(n_430), .B2(n_751), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g760 ( .A(n_109), .Y(n_760) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_343), .Y(n_109) );
NOR3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_267), .C(n_317), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_247), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_186), .B(n_228), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_164), .Y(n_114) );
INVx1_ASAP7_75t_SL g353 ( .A(n_115), .Y(n_353) );
AOI32xp33_ASAP7_75t_L g384 ( .A1(n_115), .A2(n_366), .A3(n_385), .B1(n_386), .B2(n_387), .Y(n_384) );
AND2x2_ASAP7_75t_L g386 ( .A(n_115), .B(n_243), .Y(n_386) );
AND2x4_ASAP7_75t_SL g115 ( .A(n_116), .B(n_144), .Y(n_115) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_116), .Y(n_165) );
INVx5_ASAP7_75t_L g246 ( .A(n_116), .Y(n_246) );
OR2x2_ASAP7_75t_L g253 ( .A(n_116), .B(n_245), .Y(n_253) );
INVx2_ASAP7_75t_L g258 ( .A(n_116), .Y(n_258) );
AND2x2_ASAP7_75t_L g270 ( .A(n_116), .B(n_145), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_116), .B(n_155), .Y(n_275) );
OR2x2_ASAP7_75t_L g282 ( .A(n_116), .B(n_167), .Y(n_282) );
AND2x4_ASAP7_75t_L g291 ( .A(n_116), .B(n_156), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_SL g333 ( .A1(n_116), .A2(n_249), .B(n_284), .C(n_322), .Y(n_333) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x4_ASAP7_75t_L g143 ( .A(n_119), .B(n_120), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_131), .B(n_143), .Y(n_121) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g210 ( .A(n_124), .Y(n_210) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
AND2x6_ASAP7_75t_L g139 ( .A(n_125), .B(n_134), .Y(n_139) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g141 ( .A(n_127), .B(n_136), .Y(n_141) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx5_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_129), .Y(n_526) );
AND2x2_ASAP7_75t_L g135 ( .A(n_130), .B(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
BUFx3_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
INVx2_ASAP7_75t_L g184 ( .A(n_134), .Y(n_184) );
AND2x4_ASAP7_75t_L g180 ( .A(n_135), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_142), .Y(n_137) );
INVxp67_ASAP7_75t_L g481 ( .A(n_139), .Y(n_481) );
INVxp67_ASAP7_75t_L g483 ( .A(n_141), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_142), .A2(n_149), .B(n_150), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_142), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_142), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_142), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_142), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_142), .A2(n_447), .B(n_448), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_142), .A2(n_450), .B(n_456), .C(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_142), .A2(n_450), .B(n_467), .C(n_468), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_142), .B(n_143), .Y(n_484) );
INVx1_ASAP7_75t_L g495 ( .A(n_142), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_142), .A2(n_450), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_142), .A2(n_450), .B(n_517), .C(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_143), .B(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_143), .B(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_143), .B(n_205), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g208 ( .A(n_143), .B(n_209), .C(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_143), .A2(n_454), .B(n_458), .Y(n_453) );
INVx3_ASAP7_75t_SL g283 ( .A(n_144), .Y(n_283) );
AND2x2_ASAP7_75t_L g329 ( .A(n_144), .B(n_246), .Y(n_329) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_155), .Y(n_144) );
AND2x2_ASAP7_75t_L g166 ( .A(n_145), .B(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g260 ( .A(n_145), .B(n_156), .Y(n_260) );
AND2x2_ASAP7_75t_L g264 ( .A(n_145), .B(n_243), .Y(n_264) );
INVx1_ASAP7_75t_L g290 ( .A(n_145), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_145), .B(n_156), .Y(n_312) );
INVx2_ASAP7_75t_L g316 ( .A(n_145), .Y(n_316) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_145), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_145), .B(n_246), .Y(n_393) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_152), .B(n_154), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_152), .A2(n_157), .B(n_163), .Y(n_156) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_152), .A2(n_157), .B(n_163), .Y(n_245) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_152), .A2(n_463), .B(n_469), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_153), .Y(n_152) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_153), .A2(n_214), .B(n_218), .Y(n_213) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g327 ( .A(n_156), .B(n_167), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g337 ( .A(n_165), .Y(n_337) );
NAND2xp33_ASAP7_75t_SL g362 ( .A(n_165), .B(n_254), .Y(n_362) );
AND2x2_ASAP7_75t_L g404 ( .A(n_166), .B(n_246), .Y(n_404) );
AND2x2_ASAP7_75t_L g315 ( .A(n_167), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g378 ( .A(n_167), .Y(n_378) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_168), .Y(n_243) );
AOI21x1_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_185), .Y(n_168) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_169), .A2(n_493), .B(n_501), .Y(n_492) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_169), .A2(n_493), .B(n_501), .Y(n_541) );
INVx2_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_170), .A2(n_190), .B(n_191), .Y(n_189) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_170), .A2(n_515), .B(n_519), .Y(n_514) );
BUFx4f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx3_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_179), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_174), .A2(n_180), .B1(n_199), .B2(n_201), .Y(n_198) );
INVx1_ASAP7_75t_L g534 ( .A(n_174), .Y(n_534) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_178), .Y(n_174) );
INVx1_ASAP7_75t_L g442 ( .A(n_175), .Y(n_442) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
OR2x6_ASAP7_75t_L g450 ( .A(n_176), .B(n_184), .Y(n_450) );
INVxp33_ASAP7_75t_L g498 ( .A(n_176), .Y(n_498) );
INVx1_ASAP7_75t_L g443 ( .A(n_178), .Y(n_443) );
INVxp67_ASAP7_75t_L g532 ( .A(n_180), .Y(n_532) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g499 ( .A(n_183), .Y(n_499) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_186), .A2(n_269), .B1(n_371), .B2(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_211), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_187), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_187), .B(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_196), .Y(n_187) );
INVx2_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
OR2x2_ASAP7_75t_L g238 ( .A(n_188), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_188), .B(n_251), .Y(n_256) );
AND2x4_ASAP7_75t_SL g266 ( .A(n_188), .B(n_197), .Y(n_266) );
OR2x2_ASAP7_75t_L g273 ( .A(n_188), .B(n_213), .Y(n_273) );
OR2x2_ASAP7_75t_L g285 ( .A(n_188), .B(n_197), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_188), .B(n_213), .Y(n_299) );
INVx1_ASAP7_75t_L g304 ( .A(n_188), .Y(n_304) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_188), .Y(n_322) );
AND2x2_ASAP7_75t_L g385 ( .A(n_188), .B(n_305), .Y(n_385) );
INVx2_ASAP7_75t_L g389 ( .A(n_188), .Y(n_389) );
OR2x2_ASAP7_75t_L g396 ( .A(n_188), .B(n_286), .Y(n_396) );
OR2x2_ASAP7_75t_L g418 ( .A(n_188), .B(n_419), .Y(n_418) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_195), .Y(n_188) );
AND2x2_ASAP7_75t_L g235 ( .A(n_196), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_196), .B(n_219), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_196), .B(n_295), .Y(n_357) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
AND2x4_ASAP7_75t_L g305 ( .A(n_197), .B(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_197), .B(n_250), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_197), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_197), .B(n_239), .Y(n_398) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_203), .Y(n_197) );
INVx3_ASAP7_75t_L g503 ( .A(n_206), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_206), .A2(n_503), .B1(n_522), .B2(n_527), .Y(n_521) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AOI21x1_ASAP7_75t_L g220 ( .A1(n_207), .A2(n_221), .B(n_227), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_207), .B(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_210), .A2(n_450), .B1(n_477), .B2(n_478), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_210), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g265 ( .A(n_211), .B(n_266), .Y(n_265) );
AO221x1_ASAP7_75t_L g339 ( .A1(n_211), .A2(n_254), .B1(n_285), .B2(n_340), .C(n_341), .Y(n_339) );
OAI322xp33_ASAP7_75t_L g391 ( .A1(n_211), .A2(n_311), .A3(n_392), .B1(n_394), .B2(n_395), .C1(n_396), .C2(n_397), .Y(n_391) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_219), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx3_ASAP7_75t_L g233 ( .A(n_213), .Y(n_233) );
INVx2_ASAP7_75t_L g239 ( .A(n_213), .Y(n_239) );
AND2x2_ASAP7_75t_L g251 ( .A(n_213), .B(n_219), .Y(n_251) );
INVx1_ASAP7_75t_L g296 ( .A(n_213), .Y(n_296) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_213), .Y(n_352) );
INVx1_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
OR2x2_ASAP7_75t_L g286 ( .A(n_219), .B(n_239), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_219), .Y(n_306) );
INVx1_ASAP7_75t_L g359 ( .A(n_219), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_219), .B(n_389), .Y(n_388) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_226), .Y(n_221) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI21xp33_ASAP7_75t_SL g229 ( .A1(n_230), .A2(n_237), .B(n_240), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_230), .A2(n_269), .B1(n_271), .B2(n_275), .C(n_276), .Y(n_268) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
NOR2x1p5_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g355 ( .A(n_234), .Y(n_355) );
INVx1_ASAP7_75t_SL g274 ( .A(n_235), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_235), .A2(n_380), .B(n_382), .Y(n_379) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_236), .Y(n_279) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_239), .Y(n_342) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
OAI211xp5_ASAP7_75t_L g317 ( .A1(n_242), .A2(n_318), .B(n_323), .C(n_334), .Y(n_317) );
OR2x2_ASAP7_75t_L g407 ( .A(n_242), .B(n_312), .Y(n_407) );
AND2x2_ASAP7_75t_L g409 ( .A(n_242), .B(n_275), .Y(n_409) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g249 ( .A(n_243), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g311 ( .A(n_243), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g349 ( .A(n_243), .B(n_316), .Y(n_349) );
OA33x2_ASAP7_75t_L g356 ( .A1(n_243), .A2(n_273), .A3(n_357), .B1(n_358), .B2(n_360), .B3(n_362), .Y(n_356) );
OR2x2_ASAP7_75t_L g367 ( .A(n_243), .B(n_352), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_243), .B(n_291), .Y(n_381) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g269 ( .A(n_245), .B(n_270), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_245), .A2(n_275), .B1(n_319), .B2(n_320), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g358 ( .A(n_246), .B(n_326), .C(n_359), .Y(n_358) );
AOI322xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_252), .A3(n_254), .B1(n_255), .B2(n_257), .C1(n_261), .C2(n_265), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g354 ( .A(n_250), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_251), .A2(n_266), .B(n_310), .C(n_313), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_252), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
NAND4xp25_ASAP7_75t_SL g373 ( .A(n_253), .B(n_282), .C(n_374), .D(n_376), .Y(n_373) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g263 ( .A(n_258), .Y(n_263) );
OR2x2_ASAP7_75t_L g308 ( .A(n_258), .B(n_260), .Y(n_308) );
AND2x2_ASAP7_75t_L g377 ( .A(n_259), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g382 ( .A(n_263), .B(n_377), .Y(n_382) );
BUFx2_ASAP7_75t_L g375 ( .A(n_264), .Y(n_375) );
INVx1_ASAP7_75t_SL g405 ( .A(n_265), .Y(n_405) );
AND2x4_ASAP7_75t_L g341 ( .A(n_266), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g394 ( .A(n_266), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_287), .C(n_309), .Y(n_267) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_SL g331 ( .A(n_273), .Y(n_331) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_273), .A2(n_400), .B(n_401), .C(n_410), .Y(n_399) );
OR2x2_ASAP7_75t_L g321 ( .A(n_274), .B(n_322), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B1(n_283), .B2(n_284), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_278), .B(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_281), .B(n_338), .Y(n_420) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g395 ( .A(n_282), .B(n_283), .Y(n_395) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g340 ( .A(n_286), .Y(n_340) );
AOI222xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B1(n_297), .B2(n_301), .C1(n_302), .C2(n_307), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_290), .Y(n_301) );
AND2x2_ASAP7_75t_L g348 ( .A(n_291), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_291), .A2(n_364), .B1(n_369), .B2(n_373), .Y(n_363) );
INVx2_ASAP7_75t_SL g416 ( .A(n_291), .Y(n_416) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g372 ( .A(n_296), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_296), .B(n_359), .Y(n_419) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g332 ( .A(n_300), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_302), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g370 ( .A(n_304), .Y(n_370) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_305), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g413 ( .A(n_305), .B(n_342), .Y(n_413) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g338 ( .A(n_312), .Y(n_338) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g417 ( .A(n_315), .Y(n_417) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B(n_330), .C(n_333), .Y(n_323) );
AND2x2_ASAP7_75t_SL g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g368 ( .A(n_330), .Y(n_368) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NOR3xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_383), .C(n_399), .Y(n_343) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_363), .C(n_379), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B1(n_353), .B2(n_354), .C(n_356), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_368), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g392 ( .A(n_378), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g400 ( .A(n_382), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_390), .Y(n_383) );
INVx2_ASAP7_75t_L g406 ( .A(n_385), .Y(n_406) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g397 ( .A(n_388), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_408), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_418), .B2(n_420), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
CKINVDCx11_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_423), .A2(n_431), .B1(n_751), .B2(n_760), .Y(n_759) );
OR2x6_ASAP7_75t_SL g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AND2x6_ASAP7_75t_SL g752 ( .A(n_424), .B(n_426), .Y(n_752) );
OR2x2_ASAP7_75t_L g764 ( .A(n_424), .B(n_426), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_424), .B(n_425), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AO22x1_ASAP7_75t_L g784 ( .A1(n_432), .A2(n_785), .B1(n_786), .B2(n_792), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_432), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g432 ( .A(n_433), .B(n_602), .C(n_668), .D(n_731), .Y(n_432) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_565), .Y(n_433) );
OR3x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_535), .C(n_562), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_470), .B(n_490), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_459), .Y(n_437) );
AND2x2_ASAP7_75t_L g665 ( .A(n_438), .B(n_635), .Y(n_665) );
INVx1_ASAP7_75t_L g738 ( .A(n_438), .Y(n_738) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_451), .Y(n_438) );
INVx2_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_439), .Y(n_553) );
AND2x2_ASAP7_75t_L g557 ( .A(n_439), .B(n_473), .Y(n_557) );
AND2x4_ASAP7_75t_L g573 ( .A(n_439), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g577 ( .A(n_439), .Y(n_577) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_445), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .C(n_444), .Y(n_441) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g523 ( .A(n_450), .Y(n_523) );
AND2x2_ASAP7_75t_L g471 ( .A(n_451), .B(n_472), .Y(n_471) );
INVx4_ASAP7_75t_L g554 ( .A(n_451), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_451), .B(n_544), .Y(n_558) );
INVx2_ASAP7_75t_L g572 ( .A(n_451), .Y(n_572) );
AND2x4_ASAP7_75t_L g576 ( .A(n_451), .B(n_577), .Y(n_576) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_451), .Y(n_611) );
OR2x2_ASAP7_75t_L g617 ( .A(n_451), .B(n_462), .Y(n_617) );
NOR2x1_ASAP7_75t_SL g646 ( .A(n_451), .B(n_473), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_451), .B(n_720), .Y(n_748) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AND2x2_ASAP7_75t_L g645 ( .A(n_459), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2x1_ASAP7_75t_L g679 ( .A(n_460), .B(n_472), .Y(n_679) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g486 ( .A(n_462), .Y(n_486) );
INVx2_ASAP7_75t_L g545 ( .A(n_462), .Y(n_545) );
AND2x2_ASAP7_75t_L g568 ( .A(n_462), .B(n_473), .Y(n_568) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_462), .Y(n_595) );
INVx1_ASAP7_75t_L g636 ( .A(n_462), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_485), .Y(n_470) );
AND2x2_ASAP7_75t_L g648 ( .A(n_471), .B(n_543), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_472), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g715 ( .A(n_472), .Y(n_715) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g574 ( .A(n_473), .Y(n_574) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_484), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_479) );
OAI211xp5_ASAP7_75t_SL g651 ( .A1(n_485), .A2(n_652), .B(n_656), .C(n_662), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_487), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g698 ( .A(n_487), .Y(n_698) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g620 ( .A(n_489), .B(n_574), .Y(n_620) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_511), .Y(n_490) );
AOI32xp33_ASAP7_75t_L g656 ( .A1(n_491), .A2(n_640), .A3(n_657), .B1(n_658), .B2(n_660), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
INVx2_ASAP7_75t_L g582 ( .A(n_492), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_492), .B(n_514), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_494), .B(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g594 ( .A(n_502), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_502), .B(n_520), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_502), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_502), .Y(n_712) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_510), .Y(n_502) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_503), .A2(n_504), .B(n_510), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OR2x2_ASAP7_75t_L g613 ( .A(n_511), .B(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g564 ( .A(n_512), .B(n_538), .Y(n_564) );
AND2x2_ASAP7_75t_L g713 ( .A(n_512), .B(n_711), .Y(n_713) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g550 ( .A(n_514), .Y(n_550) );
AND2x4_ASAP7_75t_L g589 ( .A(n_514), .B(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g623 ( .A(n_514), .Y(n_623) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_514), .Y(n_631) );
AND2x2_ASAP7_75t_L g640 ( .A(n_514), .B(n_520), .Y(n_640) );
INVx1_ASAP7_75t_L g724 ( .A(n_514), .Y(n_724) );
INVx2_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
INVx1_ASAP7_75t_L g588 ( .A(n_520), .Y(n_588) );
INVx1_ASAP7_75t_L g655 ( .A(n_520), .Y(n_655) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B1(n_533), .B2(n_534), .Y(n_528) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI32xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_546), .A3(n_551), .B1(n_555), .B2(n_559), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_537), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_538), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g639 ( .A(n_538), .B(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g664 ( .A(n_538), .Y(n_664) );
AND2x2_ASAP7_75t_L g745 ( .A(n_538), .B(n_587), .Y(n_745) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g560 ( .A(n_540), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g659 ( .A(n_540), .B(n_582), .Y(n_659) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_540), .B(n_561), .Y(n_681) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_540), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
INVx1_ASAP7_75t_L g614 ( .A(n_541), .Y(n_614) );
AND2x2_ASAP7_75t_L g629 ( .A(n_541), .B(n_561), .Y(n_629) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g657 ( .A(n_543), .B(n_646), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_543), .B(n_576), .Y(n_727) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_544), .Y(n_696) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_545), .Y(n_678) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g579 ( .A(n_548), .B(n_580), .Y(n_579) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_548), .B(n_664), .Y(n_663) );
NOR2xp67_ASAP7_75t_SL g750 ( .A(n_548), .B(n_688), .Y(n_750) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g607 ( .A(n_550), .B(n_561), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_551), .B(n_617), .Y(n_675) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_552), .B(n_568), .Y(n_641) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_554), .B(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g706 ( .A(n_554), .B(n_577), .Y(n_706) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_554), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_555), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
OR2x2_ASAP7_75t_L g677 ( .A(n_556), .B(n_678), .Y(n_677) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_556), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g666 ( .A(n_557), .B(n_611), .Y(n_666) );
INVxp33_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_560), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g740 ( .A(n_560), .B(n_622), .Y(n_740) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_583), .Y(n_565) );
OAI21xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B(n_578), .Y(n_566) );
AND2x2_ASAP7_75t_L g701 ( .A(n_568), .B(n_576), .Y(n_701) );
NAND2xp33_ASAP7_75t_R g569 ( .A(n_570), .B(n_575), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g743 ( .A(n_572), .Y(n_743) );
INVx4_ASAP7_75t_L g601 ( .A(n_573), .Y(n_601) );
INVx1_ASAP7_75t_L g720 ( .A(n_574), .Y(n_720) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g714 ( .A(n_576), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_SL g718 ( .A(n_576), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_579), .A2(n_644), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g608 ( .A(n_582), .B(n_594), .Y(n_608) );
AND2x2_ASAP7_75t_L g622 ( .A(n_582), .B(n_623), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_591), .B(n_596), .C(n_599), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g670 ( .A(n_586), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g598 ( .A(n_587), .Y(n_598) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g658 ( .A(n_588), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g667 ( .A(n_588), .B(n_589), .Y(n_667) );
INVx1_ASAP7_75t_L g699 ( .A(n_588), .Y(n_699) );
AND2x4_ASAP7_75t_L g680 ( .A(n_589), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g702 ( .A(n_589), .B(n_593), .Y(n_702) );
AND2x2_ASAP7_75t_L g710 ( .A(n_589), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g685 ( .A(n_593), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_593), .B(n_607), .Y(n_687) );
AND2x2_ASAP7_75t_L g690 ( .A(n_593), .B(n_640), .Y(n_690) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_594), .B(n_655), .Y(n_704) );
AND2x2_ASAP7_75t_L g632 ( .A(n_595), .B(n_620), .Y(n_632) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g728 ( .A(n_598), .B(n_608), .Y(n_728) );
BUFx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_600), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g612 ( .A(n_601), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_601), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_642), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_626), .Y(n_603) );
OAI222xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_609), .B1(n_613), .B2(n_615), .C1(n_618), .C2(n_621), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_SL g619 ( .A(n_611), .B(n_620), .Y(n_619) );
OR2x6_ASAP7_75t_L g691 ( .A(n_611), .B(n_661), .Y(n_691) );
NAND5xp2_ASAP7_75t_L g694 ( .A(n_611), .B(n_614), .C(n_630), .D(n_695), .E(n_697), .Y(n_694) );
NAND2x1_ASAP7_75t_L g730 ( .A(n_612), .B(n_616), .Y(n_730) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_617), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_619), .A2(n_710), .B1(n_713), .B2(n_714), .Y(n_709) );
INVx2_ASAP7_75t_L g661 ( .A(n_620), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_620), .B(n_636), .Y(n_673) );
INVx3_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g653 ( .A(n_622), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g686 ( .A(n_622), .Y(n_686) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g649 ( .A(n_625), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_627), .B(n_638), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_632), .B(n_633), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g637 ( .A(n_629), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_632), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x4_ASAP7_75t_SL g719 ( .A(n_636), .B(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_651), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g688 ( .A(n_659), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_662) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_692), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .C(n_682), .Y(n_669) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OA21x2_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_680), .Y(n_674) );
NAND2xp33_ASAP7_75t_SL g676 ( .A(n_677), .B(n_679), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_689), .B(n_691), .Y(n_682) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_687), .C(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_686), .A2(n_726), .B1(n_728), .B2(n_729), .Y(n_725) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_716), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g693 ( .A(n_694), .B(n_700), .C(n_707), .D(n_709), .Y(n_693) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g705 ( .A(n_696), .B(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g736 ( .A(n_699), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_703), .B2(n_705), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_705), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_721), .B(n_725), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_746), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B(n_737), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_741), .B2(n_744), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
CKINVDCx11_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_753), .A2(n_759), .B(n_761), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
BUFx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_774), .Y(n_767) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_SL g769 ( .A(n_770), .B(n_773), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_SL g797 ( .A(n_771), .B(n_773), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_771), .A2(n_802), .B(n_805), .Y(n_801) );
INVx1_ASAP7_75t_SL g795 ( .A(n_774), .Y(n_795) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx3_ASAP7_75t_L g778 ( .A(n_775), .Y(n_778) );
BUFx2_ASAP7_75t_L g806 ( .A(n_775), .Y(n_806) );
OAI21x1_ASAP7_75t_SL g776 ( .A1(n_777), .A2(n_779), .B(n_794), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .B1(n_784), .B2(n_793), .Y(n_779) );
INVx1_ASAP7_75t_L g793 ( .A(n_780), .Y(n_793) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g792 ( .A(n_786), .Y(n_792) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
CKINVDCx11_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
CKINVDCx8_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
endmodule