module real_aes_4894_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_1106;
wire n_618;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_1067;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1123;
wire n_549;
wire n_376;
wire n_694;
wire n_491;
wire n_571;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1053;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_1115;
wire n_725;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1103;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1105;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1097;
wire n_500;
wire n_601;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
INVx1_ASAP7_75t_L g633 ( .A(n_0), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_1), .A2(n_298), .B1(n_510), .B2(n_610), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_2), .A2(n_193), .B1(n_431), .B2(n_433), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_3), .A2(n_255), .B1(n_404), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_4), .A2(n_238), .B1(n_521), .B2(n_842), .Y(n_841) );
AOI21xp33_ASAP7_75t_SL g785 ( .A1(n_5), .A2(n_786), .B(n_787), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_6), .A2(n_297), .B1(n_456), .B2(n_462), .Y(n_811) );
AO22x1_ASAP7_75t_L g821 ( .A1(n_7), .A2(n_199), .B1(n_472), .B2(n_473), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_8), .A2(n_230), .B1(n_531), .B2(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g849 ( .A(n_9), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_10), .A2(n_177), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_11), .A2(n_117), .B1(n_454), .B2(n_478), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_12), .A2(n_39), .B1(n_439), .B2(n_545), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_13), .A2(n_282), .B1(n_540), .B2(n_802), .Y(n_801) );
AOI21xp33_ASAP7_75t_SL g496 ( .A1(n_14), .A2(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g641 ( .A(n_15), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_16), .A2(n_185), .B1(n_465), .B2(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_17), .B(n_342), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_18), .A2(n_153), .B1(n_505), .B2(n_506), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_19), .A2(n_259), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_20), .A2(n_162), .B1(n_531), .B2(n_541), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_21), .A2(n_113), .B1(n_459), .B2(n_461), .Y(n_1114) );
AOI21xp33_ASAP7_75t_L g584 ( .A1(n_22), .A2(n_585), .B(n_586), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_23), .A2(n_293), .B1(n_836), .B2(n_837), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_24), .A2(n_281), .B1(n_431), .B2(n_434), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_25), .A2(n_250), .B1(n_551), .B2(n_610), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_26), .A2(n_245), .B1(n_596), .B2(n_597), .C(n_598), .Y(n_595) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_27), .Y(n_342) );
INVx1_ASAP7_75t_L g480 ( .A(n_28), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_29), .A2(n_69), .B1(n_334), .B2(n_360), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_30), .A2(n_227), .B1(n_876), .B2(n_878), .Y(n_904) );
AO22x1_ASAP7_75t_L g687 ( .A1(n_31), .A2(n_134), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_32), .A2(n_738), .B(n_739), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_33), .A2(n_37), .B1(n_513), .B2(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g587 ( .A(n_34), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_35), .A2(n_130), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_36), .A2(n_197), .B1(n_459), .B2(n_461), .Y(n_1091) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_38), .A2(n_165), .B1(n_876), .B2(n_878), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_40), .A2(n_290), .B1(n_880), .B2(n_898), .Y(n_908) );
AO22x2_ASAP7_75t_L g624 ( .A1(n_41), .A2(n_625), .B1(n_630), .B2(n_650), .Y(n_624) );
INVxp33_ASAP7_75t_SL g649 ( .A(n_41), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_42), .A2(n_176), .B1(n_869), .B2(n_871), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_43), .A2(n_112), .B1(n_520), .B2(n_521), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_44), .A2(n_53), .B1(n_861), .B2(n_866), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_45), .A2(n_295), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g672 ( .A(n_46), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_47), .A2(n_93), .B1(n_607), .B2(n_615), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_48), .A2(n_684), .B(n_687), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_49), .A2(n_208), .B1(n_551), .B2(n_703), .Y(n_702) );
AOI22x1_ASAP7_75t_L g828 ( .A1(n_50), .A2(n_829), .B1(n_830), .B2(n_850), .Y(n_828) );
INVx1_ASAP7_75t_L g850 ( .A(n_50), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_51), .B(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_52), .A2(n_270), .B1(n_434), .B2(n_545), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_54), .A2(n_64), .B1(n_694), .B2(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g668 ( .A(n_55), .Y(n_668) );
OA22x2_ASAP7_75t_L g348 ( .A1(n_56), .A2(n_136), .B1(n_342), .B2(n_346), .Y(n_348) );
INVx1_ASAP7_75t_L g379 ( .A(n_56), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_57), .A2(n_100), .B1(n_335), .B2(n_552), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_58), .A2(n_187), .B1(n_551), .B2(n_610), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_59), .A2(n_310), .B1(n_439), .B2(n_607), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_60), .A2(n_242), .B1(n_880), .B2(n_881), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_61), .A2(n_71), .B1(n_540), .B2(n_725), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_62), .A2(n_97), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_63), .A2(n_145), .B1(n_698), .B2(n_699), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_65), .A2(n_207), .B1(n_367), .B2(n_439), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_66), .A2(n_120), .B1(n_513), .B2(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g500 ( .A(n_67), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_68), .A2(n_292), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_70), .A2(n_164), .B1(n_513), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_72), .A2(n_212), .B1(n_472), .B2(n_473), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_73), .A2(n_148), .B1(n_465), .B2(n_466), .Y(n_658) );
INVx1_ASAP7_75t_L g986 ( .A(n_74), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_75), .A2(n_194), .B1(n_466), .B2(n_476), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_76), .A2(n_121), .B1(n_541), .B2(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g390 ( .A(n_77), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_78), .A2(n_308), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_79), .A2(n_252), .B1(n_544), .B2(n_607), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_80), .B(n_152), .Y(n_322) );
INVx1_ASAP7_75t_L g345 ( .A(n_80), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_80), .A2(n_136), .B(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_81), .A2(n_195), .B1(n_469), .B2(n_475), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_82), .A2(n_264), .B1(n_334), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_83), .A2(n_299), .B1(n_579), .B2(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_84), .A2(n_188), .B1(n_465), .B2(n_468), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_85), .B(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_86), .A2(n_155), .B1(n_513), .B2(n_612), .Y(n_628) );
INVxp33_ASAP7_75t_L g890 ( .A(n_87), .Y(n_890) );
INVx1_ASAP7_75t_L g865 ( .A(n_88), .Y(n_865) );
AND2x4_ASAP7_75t_L g870 ( .A(n_88), .B(n_231), .Y(n_870) );
INVx1_ASAP7_75t_L g526 ( .A(n_89), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_90), .A2(n_106), .B1(n_692), .B2(n_745), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_91), .A2(n_276), .B1(n_465), .B2(n_466), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_92), .A2(n_225), .B1(n_459), .B2(n_461), .Y(n_812) );
INVx1_ASAP7_75t_L g449 ( .A(n_94), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_95), .A2(n_239), .B1(n_367), .B2(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_96), .A2(n_274), .B1(n_416), .B2(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_98), .A2(n_137), .B1(n_456), .B2(n_802), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_99), .A2(n_149), .B1(n_615), .B2(n_753), .Y(n_840) );
XOR2x2_ASAP7_75t_L g734 ( .A(n_101), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_102), .B(n_454), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_103), .A2(n_139), .B1(n_505), .B2(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g863 ( .A(n_104), .Y(n_863) );
AND2x4_ASAP7_75t_L g867 ( .A(n_104), .B(n_318), .Y(n_867) );
INVx1_ASAP7_75t_SL g877 ( .A(n_104), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_105), .A2(n_233), .B1(n_433), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_107), .A2(n_302), .B1(n_551), .B2(n_610), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_108), .A2(n_202), .B1(n_880), .B2(n_881), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_109), .A2(n_213), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_110), .A2(n_260), .B1(n_513), .B2(n_515), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_111), .A2(n_114), .B1(n_424), .B2(n_427), .Y(n_845) );
OAI22x1_ASAP7_75t_L g330 ( .A1(n_115), .A2(n_331), .B1(n_411), .B2(n_445), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_115), .B(n_332), .C(n_382), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_116), .A2(n_143), .B1(n_691), .B2(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_118), .A2(n_201), .B1(n_761), .B2(n_1087), .Y(n_1086) );
XOR2x2_ASAP7_75t_L g680 ( .A(n_119), .B(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_119), .A2(n_235), .B1(n_869), .B2(n_871), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_122), .B(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_123), .A2(n_261), .B1(n_521), .B2(n_761), .Y(n_792) );
INVx1_ASAP7_75t_L g772 ( .A(n_124), .Y(n_772) );
AO22x1_ASAP7_75t_L g819 ( .A1(n_125), .A2(n_243), .B1(n_468), .B2(n_469), .Y(n_819) );
INVx1_ASAP7_75t_L g732 ( .A(n_126), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_127), .A2(n_291), .B1(n_468), .B2(n_469), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_128), .A2(n_275), .B1(n_367), .B2(n_372), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_129), .A2(n_150), .B1(n_548), .B2(n_1089), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_131), .A2(n_296), .B1(n_360), .B2(n_510), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_132), .A2(n_262), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_133), .A2(n_306), .B1(n_861), .B2(n_866), .Y(n_860) );
INVx1_ASAP7_75t_L g359 ( .A(n_135), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_135), .B(n_181), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_135), .B(n_377), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_136), .B(n_241), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_138), .A2(n_178), .B1(n_472), .B2(n_473), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_140), .A2(n_142), .B1(n_876), .B2(n_878), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_141), .A2(n_256), .B1(n_544), .B2(n_545), .Y(n_543) );
XNOR2x1_ASAP7_75t_L g1083 ( .A(n_142), .B(n_1084), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_142), .A2(n_1106), .B1(n_1108), .B2(n_1123), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_144), .A2(n_279), .B1(n_404), .B2(n_579), .Y(n_776) );
INVx1_ASAP7_75t_L g569 ( .A(n_146), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_147), .A2(n_280), .B1(n_468), .B2(n_469), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_151), .A2(n_311), .B1(n_372), .B2(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_152), .B(n_352), .Y(n_351) );
AO22x1_ASAP7_75t_L g820 ( .A1(n_154), .A2(n_265), .B1(n_475), .B2(n_476), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_156), .A2(n_219), .B1(n_521), .B2(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_157), .B(n_686), .Y(n_784) );
XOR2x2_ASAP7_75t_SL g756 ( .A(n_158), .B(n_757), .Y(n_756) );
XOR2x2_ASAP7_75t_L g823 ( .A(n_158), .B(n_757), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_159), .A2(n_229), .B1(n_544), .B2(n_545), .Y(n_1093) );
AOI21xp33_ASAP7_75t_SL g533 ( .A1(n_160), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g767 ( .A(n_161), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_163), .A2(n_300), .B1(n_511), .B2(n_551), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_166), .A2(n_478), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_167), .A2(n_304), .B1(n_424), .B2(n_427), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_168), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g740 ( .A(n_169), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_170), .A2(n_226), .B1(n_895), .B2(n_898), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_171), .B(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_172), .A2(n_232), .B1(n_880), .B2(n_881), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_173), .A2(n_288), .B1(n_540), .B2(n_541), .Y(n_539) );
NAND2xp33_ASAP7_75t_L g452 ( .A(n_174), .B(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_175), .A2(n_234), .B1(n_518), .B2(n_548), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g1115 ( .A1(n_179), .A2(n_200), .B1(n_456), .B2(n_462), .Y(n_1115) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_180), .A2(n_286), .B1(n_416), .B2(n_847), .C(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g343 ( .A(n_181), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g909 ( .A1(n_182), .A2(n_183), .B1(n_876), .B2(n_878), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_184), .A2(n_283), .B1(n_551), .B2(n_610), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_186), .A2(n_211), .B1(n_475), .B2(n_476), .Y(n_660) );
INVx1_ASAP7_75t_L g536 ( .A(n_189), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_190), .A2(n_244), .B1(n_548), .B2(n_608), .Y(n_795) );
INVx1_ASAP7_75t_L g639 ( .A(n_191), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_192), .A2(n_196), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_198), .A2(n_268), .B1(n_424), .B2(n_427), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_203), .A2(n_263), .B1(n_596), .B2(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_204), .A2(n_216), .B1(n_414), .B2(n_419), .Y(n_413) );
XNOR2x2_ASAP7_75t_L g807 ( .A(n_205), .B(n_808), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_206), .A2(n_1109), .B1(n_1110), .B2(n_1122), .Y(n_1108) );
CKINVDCx5p33_ASAP7_75t_R g1109 ( .A(n_206), .Y(n_1109) );
INVx1_ASAP7_75t_L g771 ( .A(n_209), .Y(n_771) );
AOI21xp5_ASAP7_75t_SL g666 ( .A1(n_210), .A2(n_478), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g635 ( .A(n_214), .Y(n_635) );
INVx1_ASAP7_75t_L g987 ( .A(n_215), .Y(n_987) );
INVx1_ASAP7_75t_L g489 ( .A(n_217), .Y(n_489) );
INVx1_ASAP7_75t_L g1098 ( .A(n_218), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_220), .A2(n_223), .B1(n_439), .B2(n_442), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_221), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_222), .A2(n_246), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_224), .A2(n_305), .B1(n_513), .B2(n_615), .Y(n_722) );
INVx1_ASAP7_75t_L g768 ( .A(n_228), .Y(n_768) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_231), .Y(n_323) );
AND2x4_ASAP7_75t_L g864 ( .A(n_231), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_SL g653 ( .A(n_232), .Y(n_653) );
INVx1_ASAP7_75t_L g670 ( .A(n_236), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_237), .A2(n_269), .B1(n_392), .B2(n_419), .Y(n_844) );
INVx1_ASAP7_75t_L g774 ( .A(n_240), .Y(n_774) );
INVx1_ASAP7_75t_L g357 ( .A(n_241), .Y(n_357) );
INVxp67_ASAP7_75t_L g401 ( .A(n_241), .Y(n_401) );
INVxp67_ASAP7_75t_R g780 ( .A(n_247), .Y(n_780) );
INVx1_ASAP7_75t_L g805 ( .A(n_247), .Y(n_805) );
INVx2_ASAP7_75t_L g318 ( .A(n_248), .Y(n_318) );
INVx1_ASAP7_75t_L g674 ( .A(n_249), .Y(n_674) );
INVx1_ASAP7_75t_L g892 ( .A(n_251), .Y(n_892) );
INVx1_ASAP7_75t_L g402 ( .A(n_253), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_254), .B(n_462), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g1094 ( .A1(n_257), .A2(n_271), .B1(n_1095), .B2(n_1096), .C(n_1097), .Y(n_1094) );
INVx1_ASAP7_75t_L g815 ( .A(n_258), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_266), .A2(n_287), .B1(n_468), .B2(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g644 ( .A(n_267), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_272), .A2(n_278), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g896 ( .A(n_273), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_277), .B(n_689), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_284), .A2(n_383), .B(n_389), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_285), .A2(n_294), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g664 ( .A(n_289), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_290), .Y(n_592) );
AOI21xp33_ASAP7_75t_SL g477 ( .A1(n_301), .A2(n_478), .B(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_303), .A2(n_309), .B1(n_534), .B2(n_800), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_307), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_324), .B(n_853), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_316), .B(n_1103), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_316), .B(n_1104), .Y(n_1107) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OA21x2_ASAP7_75t_L g1124 ( .A1(n_317), .A2(n_877), .B(n_1125), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g862 ( .A(n_318), .B(n_863), .Y(n_862) );
AND3x4_ASAP7_75t_L g876 ( .A(n_318), .B(n_864), .C(n_877), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_319), .B(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_320), .A2(n_408), .B(n_409), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g1104 ( .A(n_323), .Y(n_1104) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_709), .B2(n_710), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
XNOR2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_621), .Y(n_326) );
XOR2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_484), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OA22x2_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_446), .B1(n_447), .B2(n_483), .Y(n_329) );
INVx2_ASAP7_75t_L g483 ( .A(n_330), .Y(n_483) );
AND4x1_ASAP7_75t_L g445 ( .A(n_332), .B(n_382), .C(n_412), .D(n_429), .Y(n_445) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_366), .Y(n_332) );
BUFx4f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_337), .Y(n_510) );
BUFx12f_ASAP7_75t_L g551 ( .A(n_337), .Y(n_551) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_349), .Y(n_337) );
AND2x2_ASAP7_75t_L g363 ( .A(n_338), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g368 ( .A(n_338), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g440 ( .A(n_338), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g472 ( .A(n_338), .B(n_349), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_338), .B(n_364), .Y(n_473) );
AND2x4_ASAP7_75t_L g475 ( .A(n_338), .B(n_369), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_338), .B(n_436), .Y(n_476) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_347), .Y(n_338) );
AND2x2_ASAP7_75t_L g418 ( .A(n_339), .B(n_348), .Y(n_418) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_348), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
NAND2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx2_ASAP7_75t_L g346 ( .A(n_342), .Y(n_346) );
INVx3_ASAP7_75t_L g352 ( .A(n_342), .Y(n_352) );
NAND2xp33_ASAP7_75t_L g358 ( .A(n_342), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g381 ( .A(n_342), .Y(n_381) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_342), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_343), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_345), .A2(n_381), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g399 ( .A(n_348), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g417 ( .A(n_349), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g422 ( .A(n_349), .B(n_388), .Y(n_422) );
AND2x4_ASAP7_75t_L g456 ( .A(n_349), .B(n_388), .Y(n_456) );
AND2x4_ASAP7_75t_L g461 ( .A(n_349), .B(n_418), .Y(n_461) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .Y(n_349) );
INVx2_ASAP7_75t_L g365 ( .A(n_350), .Y(n_365) );
AND2x4_ASAP7_75t_L g369 ( .A(n_350), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g395 ( .A(n_350), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g437 ( .A(n_350), .B(n_371), .Y(n_437) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_352), .B(n_357), .Y(n_356) );
INVxp67_ASAP7_75t_L g377 ( .A(n_352), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_353), .B(n_376), .C(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g364 ( .A(n_354), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g371 ( .A(n_355), .Y(n_371) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g834 ( .A(n_361), .Y(n_834) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx5_ASAP7_75t_L g511 ( .A(n_363), .Y(n_511) );
BUFx3_ASAP7_75t_L g552 ( .A(n_363), .Y(n_552) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_363), .Y(n_610) );
AND2x2_ASAP7_75t_L g387 ( .A(n_364), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g426 ( .A(n_364), .B(n_418), .Y(n_426) );
AND2x4_ASAP7_75t_L g428 ( .A(n_364), .B(n_375), .Y(n_428) );
AND2x2_ASAP7_75t_L g454 ( .A(n_364), .B(n_388), .Y(n_454) );
AND2x4_ASAP7_75t_L g459 ( .A(n_364), .B(n_375), .Y(n_459) );
AND2x2_ASAP7_75t_L g478 ( .A(n_364), .B(n_418), .Y(n_478) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx12f_ASAP7_75t_L g548 ( .A(n_368), .Y(n_548) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_368), .Y(n_607) );
AND2x4_ASAP7_75t_L g374 ( .A(n_369), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g432 ( .A(n_369), .B(n_388), .Y(n_432) );
AND2x4_ASAP7_75t_L g468 ( .A(n_369), .B(n_388), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_369), .B(n_375), .Y(n_469) );
AND2x2_ASAP7_75t_L g514 ( .A(n_369), .B(n_388), .Y(n_514) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g515 ( .A(n_373), .Y(n_515) );
INVx1_ASAP7_75t_L g549 ( .A(n_373), .Y(n_549) );
INVx4_ASAP7_75t_L g615 ( .A(n_373), .Y(n_615) );
INVx2_ASAP7_75t_L g707 ( .A(n_373), .Y(n_707) );
INVx4_ASAP7_75t_L g764 ( .A(n_373), .Y(n_764) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_373), .Y(n_1089) );
INVx8_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g444 ( .A(n_375), .B(n_441), .Y(n_444) );
AND2x4_ASAP7_75t_L g466 ( .A(n_375), .B(n_441), .Y(n_466) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g775 ( .A(n_385), .Y(n_775) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g583 ( .A(n_386), .Y(n_583) );
INVx2_ASAP7_75t_L g597 ( .A(n_386), .Y(n_597) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g495 ( .A(n_387), .Y(n_495) );
BUFx3_ASAP7_75t_L g731 ( .A(n_387), .Y(n_731) );
AND2x4_ASAP7_75t_L g435 ( .A(n_388), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g465 ( .A(n_388), .B(n_441), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_402), .B2(n_403), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g506 ( .A(n_393), .Y(n_506) );
INVx2_ASAP7_75t_L g688 ( .A(n_393), .Y(n_688) );
INVx4_ASAP7_75t_L g725 ( .A(n_393), .Y(n_725) );
INVx2_ASAP7_75t_L g802 ( .A(n_393), .Y(n_802) );
INVx5_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g532 ( .A(n_394), .Y(n_532) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_394), .Y(n_579) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_399), .Y(n_394) );
AND2x4_ASAP7_75t_L g462 ( .A(n_395), .B(n_399), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g408 ( .A(n_397), .Y(n_408) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx4_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_405), .B(n_815), .Y(n_814) );
INVx4_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g588 ( .A(n_406), .Y(n_588) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_407), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_429), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_423), .Y(n_412) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g498 ( .A(n_417), .Y(n_498) );
BUFx3_ASAP7_75t_L g531 ( .A(n_417), .Y(n_531) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_417), .Y(n_596) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g747 ( .A(n_420), .Y(n_747) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g581 ( .A(n_421), .Y(n_581) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g505 ( .A(n_422), .Y(n_505) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_422), .Y(n_540) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_SL g1095 ( .A(n_425), .Y(n_1095) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_426), .Y(n_534) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_426), .Y(n_585) );
BUFx3_ASAP7_75t_L g602 ( .A(n_426), .Y(n_602) );
INVx2_ASAP7_75t_L g729 ( .A(n_426), .Y(n_729) );
BUFx3_ASAP7_75t_L g692 ( .A(n_427), .Y(n_692) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_428), .Y(n_541) );
INVx3_ASAP7_75t_L g604 ( .A(n_428), .Y(n_604) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_438), .Y(n_429) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx4f_ASAP7_75t_L g1087 ( .A(n_432), .Y(n_1087) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx12f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_435), .Y(n_520) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_435), .Y(n_612) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_435), .Y(n_761) );
BUFx3_ASAP7_75t_L g842 ( .A(n_435), .Y(n_842) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g441 ( .A(n_437), .Y(n_441) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_440), .Y(n_518) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_440), .Y(n_544) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_440), .Y(n_608) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx5_ASAP7_75t_L g545 ( .A(n_443), .Y(n_545) );
INVx2_ASAP7_75t_L g573 ( .A(n_443), .Y(n_573) );
INVx2_ASAP7_75t_L g613 ( .A(n_443), .Y(n_613) );
INVx6_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx12f_ASAP7_75t_L g521 ( .A(n_444), .Y(n_521) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
XNOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NOR2x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_463), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .C(n_460), .Y(n_451) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g665 ( .A(n_454), .Y(n_665) );
INVx1_ASAP7_75t_L g675 ( .A(n_456), .Y(n_675) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_458), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g671 ( .A(n_461), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g463 ( .A(n_464), .B(n_467), .C(n_470), .D(n_477), .Y(n_463) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_481), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_481), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g648 ( .A(n_481), .Y(n_648) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g502 ( .A(n_482), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_482), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_SL g689 ( .A(n_482), .Y(n_689) );
INVx1_ASAP7_75t_L g743 ( .A(n_482), .Y(n_743) );
BUFx6f_ASAP7_75t_L g1099 ( .A(n_482), .Y(n_1099) );
XNOR2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_563), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_522), .B1(n_559), .B2(n_561), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g562 ( .A(n_487), .Y(n_562) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
XNOR2x1_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
NOR4xp75_ASAP7_75t_L g490 ( .A(n_491), .B(n_503), .C(n_508), .D(n_516), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
INVx2_ASAP7_75t_L g686 ( .A(n_494), .Y(n_686) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g646 ( .A(n_495), .Y(n_646) );
INVx2_ASAP7_75t_L g640 ( .A(n_497), .Y(n_640) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g786 ( .A(n_498), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_501), .B(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
BUFx2_ASAP7_75t_L g695 ( .A(n_505), .Y(n_695) );
INVx2_ASAP7_75t_L g769 ( .A(n_505), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_512), .Y(n_508) );
BUFx3_ASAP7_75t_L g703 ( .A(n_511), .Y(n_703) );
BUFx3_ASAP7_75t_L g701 ( .A(n_513), .Y(n_701) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx8_ASAP7_75t_L g753 ( .A(n_514), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_517), .B(n_519), .Y(n_516) );
INVx1_ASAP7_75t_L g838 ( .A(n_518), .Y(n_838) );
BUFx3_ASAP7_75t_L g699 ( .A(n_521), .Y(n_699) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_527), .B(n_553), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_525), .B(n_539), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
NOR2xp67_ASAP7_75t_L g527 ( .A(n_528), .B(n_542), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_537), .C(n_539), .Y(n_528) );
INVx1_ASAP7_75t_L g557 ( .A(n_529), .Y(n_557) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_533), .Y(n_529) );
BUFx2_ASAP7_75t_L g694 ( .A(n_531), .Y(n_694) );
INVxp67_ASAP7_75t_L g741 ( .A(n_532), .Y(n_741) );
BUFx3_ASAP7_75t_L g691 ( .A(n_534), .Y(n_691) );
INVxp67_ASAP7_75t_L g555 ( .A(n_537), .Y(n_555) );
INVx3_ASAP7_75t_L g642 ( .A(n_540), .Y(n_642) );
INVx1_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .C(n_547), .D(n_550), .Y(n_542) );
BUFx12f_ASAP7_75t_L g836 ( .A(n_548), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_589), .B1(n_616), .B2(n_619), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g620 ( .A(n_568), .Y(n_620) );
XNOR2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_577), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .C(n_575), .D(n_576), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .C(n_582), .D(n_584), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_588), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g618 ( .A(n_591), .Y(n_618) );
XNOR2x1_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_605), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_600), .C(n_601), .Y(n_594) );
INVx2_ASAP7_75t_L g634 ( .A(n_602), .Y(n_634) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g637 ( .A(n_604), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_604), .A2(n_634), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx3_ASAP7_75t_L g800 ( .A(n_604), .Y(n_800) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_606), .B(n_609), .C(n_611), .D(n_614), .Y(n_605) );
BUFx2_ASAP7_75t_SL g705 ( .A(n_607), .Y(n_705) );
BUFx3_ASAP7_75t_L g698 ( .A(n_608), .Y(n_698) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI22x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_679), .B1(n_680), .B2(n_708), .Y(n_622) );
INVx2_ASAP7_75t_L g708 ( .A(n_623), .Y(n_708) );
AO22x2_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_651), .B1(n_677), .B2(n_678), .Y(n_623) );
INVx2_ASAP7_75t_L g678 ( .A(n_624), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_625), .B(n_631), .Y(n_650) );
AND4x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .C(n_628), .D(n_629), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_649), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_638), .C(n_643), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_635), .B2(n_636), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_640), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_766) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_647), .Y(n_643) );
INVxp67_ASAP7_75t_L g738 ( .A(n_645), .Y(n_738) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_649), .A2(n_894), .B1(n_896), .B2(n_897), .Y(n_893) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
XNOR2x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_653), .B(n_654), .Y(n_677) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_662), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_669), .C(n_673), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_666), .Y(n_663) );
INVx2_ASAP7_75t_L g1096 ( .A(n_665), .Y(n_1096) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B(n_676), .Y(n_673) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_696), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_690), .C(n_693), .Y(n_682) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND4xp25_ASAP7_75t_SL g696 ( .A(n_697), .B(n_700), .C(n_702), .D(n_704), .Y(n_696) );
BUFx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_754), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AO22x2_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_733), .B2(n_734), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
XOR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_732), .Y(n_716) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_723), .Y(n_717) );
NAND4xp25_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .C(n_721), .D(n_722), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .C(n_727), .D(n_730), .Y(n_723) );
INVx3_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g745 ( .A(n_729), .Y(n_745) );
BUFx3_ASAP7_75t_L g847 ( .A(n_731), .Y(n_847) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_748), .Y(n_735) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_744), .C(n_746), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_742), .Y(n_739) );
NAND4xp25_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .C(n_751), .D(n_752), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_825), .B1(n_851), .B2(n_852), .Y(n_754) );
INVx1_ASAP7_75t_L g851 ( .A(n_755), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_777), .B1(n_822), .B2(n_824), .Y(n_755) );
AND2x4_ASAP7_75t_L g757 ( .A(n_758), .B(n_765), .Y(n_757) );
AND4x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .C(n_762), .D(n_763), .Y(n_758) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_770), .C(n_773), .Y(n_765) );
OAI21xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B(n_776), .Y(n_773) );
INVx2_ASAP7_75t_L g824 ( .A(n_777), .Y(n_824) );
OA22x2_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_806), .B2(n_807), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI21x1_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B(n_803), .Y(n_779) );
NOR4xp75_ASAP7_75t_L g781 ( .A(n_782), .B(n_789), .C(n_793), .D(n_797), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g803 ( .A(n_783), .B(n_790), .C(n_794), .D(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AND2x2_ASAP7_75t_L g804 ( .A(n_798), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_816), .Y(n_808) );
AND4x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .C(n_812), .D(n_813), .Y(n_809) );
NOR4xp25_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .C(n_820), .D(n_821), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g852 ( .A(n_825), .Y(n_852) );
BUFx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NAND4xp75_ASAP7_75t_L g830 ( .A(n_831), .B(n_839), .C(n_843), .D(n_846), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_1076), .B1(n_1077), .B2(n_1101), .C(n_1105), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_948), .B(n_989), .C(n_1032), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_918), .C(n_925), .Y(n_855) );
AOI222xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_885), .B1(n_899), .B2(n_906), .C1(n_910), .C2(n_915), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_857), .B(n_907), .Y(n_1045) );
AND2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_872), .Y(n_857) );
INVx1_ASAP7_75t_L g900 ( .A(n_858), .Y(n_900) );
NAND2xp5_ASAP7_75t_SL g922 ( .A(n_858), .B(n_923), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_858), .B(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g939 ( .A(n_858), .Y(n_939) );
INVx2_ASAP7_75t_L g951 ( .A(n_858), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_858), .B(n_913), .Y(n_961) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_858), .Y(n_969) );
AND2x2_ASAP7_75t_L g994 ( .A(n_858), .B(n_982), .Y(n_994) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_858), .B(n_886), .Y(n_1024) );
NOR2x1_ASAP7_75t_L g1035 ( .A(n_858), .B(n_924), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_858), .B(n_887), .Y(n_1043) );
NAND2xp5_ASAP7_75t_SL g1063 ( .A(n_858), .B(n_1064), .Y(n_1063) );
INVx4_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_859), .B(n_902), .Y(n_911) );
OR2x2_ASAP7_75t_L g927 ( .A(n_859), .B(n_928), .Y(n_927) );
AND2x2_ASAP7_75t_L g933 ( .A(n_859), .B(n_887), .Y(n_933) );
AND2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_868), .Y(n_859) );
INVx3_ASAP7_75t_L g889 ( .A(n_861), .Y(n_889) );
AND2x4_ASAP7_75t_L g861 ( .A(n_862), .B(n_864), .Y(n_861) );
AND2x2_ASAP7_75t_L g869 ( .A(n_862), .B(n_870), .Y(n_869) );
AND2x2_ASAP7_75t_L g880 ( .A(n_862), .B(n_870), .Y(n_880) );
AND2x4_ASAP7_75t_L g895 ( .A(n_862), .B(n_870), .Y(n_895) );
AND2x4_ASAP7_75t_L g866 ( .A(n_864), .B(n_867), .Y(n_866) );
AND2x4_ASAP7_75t_L g878 ( .A(n_864), .B(n_867), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_864), .B(n_867), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g1125 ( .A(n_864), .Y(n_1125) );
AND2x2_ASAP7_75t_L g871 ( .A(n_867), .B(n_870), .Y(n_871) );
AND2x2_ASAP7_75t_L g881 ( .A(n_867), .B(n_870), .Y(n_881) );
AND2x4_ASAP7_75t_L g898 ( .A(n_867), .B(n_870), .Y(n_898) );
AND2x2_ASAP7_75t_L g940 ( .A(n_872), .B(n_928), .Y(n_940) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_872), .B(n_914), .Y(n_1029) );
INVx1_ASAP7_75t_L g1068 ( .A(n_872), .Y(n_1068) );
AND2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_882), .Y(n_872) );
AND2x2_ASAP7_75t_L g906 ( .A(n_873), .B(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g913 ( .A(n_873), .B(n_914), .Y(n_913) );
OR2x2_ASAP7_75t_L g924 ( .A(n_873), .B(n_882), .Y(n_924) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OR2x2_ASAP7_75t_L g954 ( .A(n_874), .B(n_882), .Y(n_954) );
AND2x2_ASAP7_75t_L g960 ( .A(n_874), .B(n_882), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_874), .B(n_914), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_874), .B(n_907), .Y(n_1018) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_879), .Y(n_874) );
INVx1_ASAP7_75t_L g936 ( .A(n_882), .Y(n_936) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_882), .B(n_928), .Y(n_1073) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_885), .B(n_920), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_885), .B(n_942), .Y(n_971) );
NOR2xp33_ASAP7_75t_L g1066 ( .A(n_885), .B(n_1067), .Y(n_1066) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g902 ( .A(n_887), .Y(n_902) );
AND2x2_ASAP7_75t_L g956 ( .A(n_887), .B(n_903), .Y(n_956) );
OR2x2_ASAP7_75t_L g966 ( .A(n_887), .B(n_903), .Y(n_966) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_887), .B(n_1051), .Y(n_1050) );
OR2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_893), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g985 ( .A1(n_889), .A2(n_891), .B1(n_986), .B2(n_987), .C(n_988), .Y(n_985) );
BUFx2_ASAP7_75t_L g1076 ( .A(n_891), .Y(n_1076) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVxp67_ASAP7_75t_L g1041 ( .A(n_899), .Y(n_1041) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_900), .B(n_917), .Y(n_978) );
OAI322xp33_ASAP7_75t_L g926 ( .A1(n_901), .A2(n_923), .A3(n_927), .B1(n_930), .B2(n_931), .C1(n_932), .C2(n_934), .Y(n_926) );
OAI211xp5_ASAP7_75t_SL g948 ( .A1(n_901), .A2(n_949), .B(n_955), .C(n_972), .Y(n_948) );
INVx1_ASAP7_75t_L g1015 ( .A(n_901), .Y(n_1015) );
OR2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
AND2x2_ASAP7_75t_L g975 ( .A(n_902), .B(n_964), .Y(n_975) );
AND2x2_ASAP7_75t_L g980 ( .A(n_902), .B(n_903), .Y(n_980) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_902), .B(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1054 ( .A(n_902), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_903), .Y(n_917) );
INVx2_ASAP7_75t_L g930 ( .A(n_903), .Y(n_930) );
OR2x2_ASAP7_75t_L g997 ( .A(n_903), .B(n_944), .Y(n_997) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_903), .B(n_945), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_903), .B(n_944), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_903), .B(n_943), .Y(n_1075) );
AND2x2_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_906), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g1005 ( .A(n_906), .B(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g914 ( .A(n_907), .Y(n_914) );
INVx1_ASAP7_75t_SL g929 ( .A(n_907), .Y(n_929) );
OR2x2_ASAP7_75t_L g953 ( .A(n_907), .B(n_954), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_907), .B(n_923), .Y(n_974) );
AND2x2_ASAP7_75t_L g982 ( .A(n_907), .B(n_936), .Y(n_982) );
OR2x2_ASAP7_75t_L g1007 ( .A(n_907), .B(n_924), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_907), .B(n_1035), .Y(n_1034) );
AND2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_911), .B(n_1018), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_912), .A2(n_922), .B1(n_1011), .B2(n_1013), .C(n_1016), .Y(n_1010) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
NOR2x1_ASAP7_75t_R g921 ( .A(n_914), .B(n_922), .Y(n_921) );
AND2x2_ASAP7_75t_L g935 ( .A(n_914), .B(n_936), .Y(n_935) );
AND2x2_ASAP7_75t_L g959 ( .A(n_914), .B(n_960), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_914), .B(n_1047), .Y(n_1046) );
OAI322xp33_ASAP7_75t_L g1004 ( .A1(n_915), .A2(n_938), .A3(n_969), .B1(n_997), .B2(n_1005), .C1(n_1008), .C2(n_1009), .Y(n_1004) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_917), .B(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVxp67_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
OAI21xp5_ASAP7_75t_SL g1028 ( .A1(n_923), .A2(n_1029), .B(n_1030), .Y(n_1028) );
INVx3_ASAP7_75t_SL g923 ( .A(n_924), .Y(n_923) );
OAI21xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_937), .B(n_941), .Y(n_925) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_927), .B(n_1068), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_928), .B(n_960), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_928), .B(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_930), .A2(n_931), .B1(n_992), .B2(n_993), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_930), .A2(n_995), .B1(n_1053), .B2(n_1055), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_930), .B(n_933), .Y(n_1071) );
O2A1O1Ixp33_ASAP7_75t_L g967 ( .A1(n_931), .A2(n_968), .B(n_970), .C(n_971), .Y(n_967) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NOR2xp67_ASAP7_75t_SL g1053 ( .A(n_938), .B(n_1054), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_938), .B(n_1056), .Y(n_1055) );
NAND2xp67_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_939), .B(n_960), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_939), .B(n_956), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_940), .A2(n_956), .B1(n_957), .B2(n_962), .C(n_967), .Y(n_955) );
INVx1_ASAP7_75t_L g1008 ( .A(n_940), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1014 ( .A(n_941), .B(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_942), .A2(n_1051), .B1(n_1058), .B2(n_1059), .C(n_1069), .Y(n_1057) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g964 ( .A(n_945), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
INVx1_ASAP7_75t_L g999 ( .A(n_951), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_951), .B(n_953), .Y(n_1003) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1021 ( .A(n_954), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_954), .B(n_1048), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_961), .Y(n_957) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_958), .A2(n_997), .B1(n_1070), .B2(n_1072), .C(n_1074), .Y(n_1069) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_959), .B(n_1015), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_959), .B(n_968), .Y(n_1058) );
INVx1_ASAP7_75t_L g1048 ( .A(n_960), .Y(n_1048) );
INVx1_ASAP7_75t_L g1009 ( .A(n_962), .Y(n_1009) );
AND2x2_ASAP7_75t_L g962 ( .A(n_963), .B(n_965), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_963), .A2(n_973), .B1(n_975), .B2(n_976), .C(n_983), .Y(n_972) );
INVx2_ASAP7_75t_L g995 ( .A(n_963), .Y(n_995) );
BUFx3_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_964), .B(n_966), .Y(n_1012) );
INVx2_ASAP7_75t_L g1025 ( .A(n_964), .Y(n_1025) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_969), .B(n_980), .Y(n_992) );
INVx1_ASAP7_75t_L g1002 ( .A(n_971), .Y(n_1002) );
OAI21xp33_ASAP7_75t_L g1074 ( .A1(n_973), .A2(n_1017), .B(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_979), .B2(n_981), .Y(n_976) );
A2O1A1Ixp33_ASAP7_75t_L g1059 ( .A1(n_979), .A2(n_1060), .B(n_1061), .C(n_1065), .Y(n_1059) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AOI211xp5_ASAP7_75t_L g1019 ( .A1(n_984), .A2(n_1020), .B(n_1022), .C(n_1026), .Y(n_1019) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
NAND4xp25_ASAP7_75t_L g989 ( .A(n_990), .B(n_1001), .C(n_1019), .D(n_1028), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_995), .B(n_996), .Y(n_990) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g1061 ( .A(n_994), .B(n_1062), .Y(n_1061) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_999), .B(n_1000), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_1000), .B(n_1029), .Y(n_1039) );
AOI211xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1003), .B(n_1004), .C(n_1010), .Y(n_1001) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVxp67_ASAP7_75t_SL g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1018), .Y(n_1064) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1025), .B(n_1043), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1029), .Y(n_1060) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND3xp33_ASAP7_75t_SL g1032 ( .A(n_1033), .B(n_1052), .C(n_1057), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_1034), .A2(n_1036), .B1(n_1038), .B2(n_1040), .C(n_1044), .Y(n_1033) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_SL g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
AOI21xp33_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1046), .B(n_1049), .Y(n_1044) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1054), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1054), .B(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NOR2x1_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1092), .Y(n_1084) );
NAND4xp25_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .C(n_1090), .D(n_1091), .Y(n_1085) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .C(n_1100), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1099), .Y(n_1097) );
CKINVDCx16_ASAP7_75t_R g1101 ( .A(n_1102), .Y(n_1101) );
BUFx3_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVxp67_ASAP7_75t_SL g1122 ( .A(n_1110), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1117), .Y(n_1111) );
NAND4xp25_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .C(n_1115), .D(n_1116), .Y(n_1112) );
NAND4xp25_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1119), .C(n_1120), .D(n_1121), .Y(n_1117) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
endmodule