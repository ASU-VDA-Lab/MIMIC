module real_aes_4687_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_0), .A2(n_19), .B1(n_281), .B2(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_1), .A2(n_65), .B1(n_352), .B2(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_3), .A2(n_21), .B1(n_167), .B2(n_169), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_4), .A2(n_20), .B1(n_340), .B2(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g325 ( .A(n_5), .Y(n_325) );
INVx1_ASAP7_75t_L g103 ( .A(n_6), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_6), .B(n_48), .Y(n_122) );
INVxp67_ASAP7_75t_L g165 ( .A(n_6), .Y(n_165) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_46), .B(n_251), .Y(n_250) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_7), .A2(n_46), .B(n_251), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g99 ( .A(n_8), .B(n_88), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_9), .B(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_9), .Y(n_649) );
INVx1_ASAP7_75t_SL g322 ( .A(n_10), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_11), .B(n_343), .Y(n_342) );
BUFx3_ASAP7_75t_L g206 ( .A(n_12), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_13), .A2(n_79), .B1(n_80), .B2(n_655), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_13), .Y(n_655) );
O2A1O1Ixp5_ASAP7_75t_L g275 ( .A1(n_14), .A2(n_227), .B(n_276), .C(n_279), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_15), .B(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_16), .Y(n_88) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_17), .Y(n_197) );
INVx1_ASAP7_75t_L g92 ( .A(n_18), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_18), .B(n_47), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_22), .A2(n_26), .B1(n_355), .B2(n_368), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_23), .A2(n_45), .B1(n_290), .B2(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_24), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_24), .Y(n_663) );
INVx2_ASAP7_75t_L g377 ( .A(n_25), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_27), .B(n_294), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_28), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_29), .A2(n_319), .B(n_320), .C(n_323), .Y(n_318) );
INVx1_ASAP7_75t_L g254 ( .A(n_30), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_31), .A2(n_43), .B1(n_132), .B2(n_137), .Y(n_131) );
INVx2_ASAP7_75t_L g292 ( .A(n_32), .Y(n_292) );
INVx1_ASAP7_75t_L g251 ( .A(n_33), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_34), .A2(n_37), .B1(n_155), .B2(n_157), .Y(n_154) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_35), .Y(n_217) );
AND2x4_ASAP7_75t_L g231 ( .A(n_35), .B(n_215), .Y(n_231) );
AND2x4_ASAP7_75t_L g304 ( .A(n_35), .B(n_215), .Y(n_304) );
INVx2_ASAP7_75t_L g384 ( .A(n_36), .Y(n_384) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_38), .Y(n_229) );
INVx1_ASAP7_75t_SL g280 ( .A(n_39), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_40), .A2(n_64), .B1(n_145), .B2(n_151), .Y(n_144) );
OA22x2_ASAP7_75t_L g86 ( .A1(n_41), .A2(n_48), .B1(n_87), .B2(n_88), .Y(n_86) );
INVx1_ASAP7_75t_L g129 ( .A(n_41), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_42), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_44), .A2(n_70), .B1(n_178), .B2(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g105 ( .A(n_47), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_47), .B(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_47), .Y(n_209) );
OAI21xp33_ASAP7_75t_L g141 ( .A1(n_48), .A2(n_58), .B(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_49), .A2(n_281), .B(n_323), .C(n_386), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_50), .Y(n_192) );
AOI221x1_ASAP7_75t_SL g82 ( .A1(n_51), .A2(n_52), .B1(n_83), .B2(n_106), .C(n_113), .Y(n_82) );
INVx1_ASAP7_75t_L g247 ( .A(n_53), .Y(n_247) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_54), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_55), .B(n_340), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_56), .B(n_314), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_57), .A2(n_248), .B(n_381), .C(n_383), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g425 ( .A1(n_57), .A2(n_248), .B(n_381), .C(n_383), .Y(n_425) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_58), .B(n_69), .Y(n_123) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_59), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_60), .A2(n_68), .B1(n_244), .B2(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_61), .Y(n_224) );
BUFx5_ASAP7_75t_L g245 ( .A(n_61), .Y(n_245) );
INVx1_ASAP7_75t_L g284 ( .A(n_61), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_62), .B(n_262), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_63), .A2(n_72), .B1(n_173), .B2(n_175), .Y(n_172) );
INVx2_ASAP7_75t_SL g215 ( .A(n_66), .Y(n_215) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_67), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_69), .B(n_98), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_71), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_SL g372 ( .A(n_73), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_74), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g406 ( .A(n_75), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g291 ( .A(n_76), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_201), .B1(n_218), .B2(n_232), .C(n_647), .Y(n_77) );
OAI22xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_80), .B1(n_183), .B2(n_184), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_79), .A2(n_80), .B1(n_649), .B2(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_81), .Y(n_80) );
NAND4xp75_ASAP7_75t_L g81 ( .A(n_82), .B(n_130), .C(n_153), .D(n_171), .Y(n_81) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AND2x4_ASAP7_75t_L g84 ( .A(n_85), .B(n_95), .Y(n_84) );
AND2x4_ASAP7_75t_L g168 ( .A(n_85), .B(n_111), .Y(n_168) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_89), .Y(n_85) );
AND2x2_ASAP7_75t_L g110 ( .A(n_86), .B(n_90), .Y(n_110) );
INVx1_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
AND2x2_ASAP7_75t_L g163 ( .A(n_86), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g93 ( .A(n_87), .B(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
NAND2xp33_ASAP7_75t_L g91 ( .A(n_88), .B(n_92), .Y(n_91) );
INVx3_ASAP7_75t_L g98 ( .A(n_88), .Y(n_98) );
NAND2xp33_ASAP7_75t_L g104 ( .A(n_88), .B(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_88), .Y(n_120) );
INVx1_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
AND2x4_ASAP7_75t_L g147 ( .A(n_89), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_91), .B(n_93), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_92), .B(n_129), .Y(n_128) );
INVxp67_ASAP7_75t_L g210 ( .A(n_92), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_94), .A2(n_142), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g156 ( .A(n_95), .B(n_110), .Y(n_156) );
AND2x4_ASAP7_75t_L g174 ( .A(n_95), .B(n_147), .Y(n_174) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_100), .Y(n_95) );
INVx2_ASAP7_75t_L g112 ( .A(n_96), .Y(n_112) );
OR2x2_ASAP7_75t_L g135 ( .A(n_96), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g149 ( .A(n_96), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g160 ( .A(n_96), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_99), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_98), .B(n_103), .Y(n_102) );
INVxp67_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
NAND3xp33_ASAP7_75t_L g124 ( .A(n_99), .B(n_125), .C(n_127), .Y(n_124) );
AND2x4_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x4_ASAP7_75t_L g133 ( .A(n_110), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g179 ( .A(n_110), .B(n_149), .Y(n_179) );
AND2x4_ASAP7_75t_L g170 ( .A(n_111), .B(n_140), .Y(n_170) );
AND2x2_ASAP7_75t_L g176 ( .A(n_111), .B(n_147), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_121), .B(n_124), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_120), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_126), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g140 ( .A(n_127), .B(n_141), .Y(n_140) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_129), .Y(n_211) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_144), .Y(n_130) );
BUFx12f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g150 ( .A(n_136), .Y(n_150) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx6_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_143), .Y(n_139) );
AND2x4_ASAP7_75t_L g182 ( .A(n_140), .B(n_149), .Y(n_182) );
AND2x4_ASAP7_75t_L g152 ( .A(n_143), .B(n_147), .Y(n_152) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_166), .Y(n_153) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_163), .Y(n_159) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
BUFx8_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_177), .Y(n_171) );
BUFx12f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx8_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
XOR2xp5_ASAP7_75t_SL g184 ( .A(n_185), .B(n_195), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_193), .B2(n_194), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_186), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_187), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B1(n_198), .B2(n_199), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_197), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_200), .B(n_290), .Y(n_386) );
BUFx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_212), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g652 ( .A(n_205), .B(n_212), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .C(n_211), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_216), .Y(n_212) );
OR2x2_ASAP7_75t_L g657 ( .A(n_213), .B(n_217), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_213), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_213), .B(n_216), .Y(n_661) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_230), .Y(n_218) );
OA21x2_ASAP7_75t_L g659 ( .A1(n_219), .A2(n_660), .B(n_661), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_225), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_222), .A2(n_289), .B1(n_291), .B2(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_223), .Y(n_319) );
INVx2_ASAP7_75t_L g399 ( .A(n_223), .Y(n_399) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx6_ASAP7_75t_L g257 ( .A(n_224), .Y(n_257) );
INVx2_ASAP7_75t_L g263 ( .A(n_224), .Y(n_263) );
INVx3_ASAP7_75t_L g315 ( .A(n_224), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_227), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_227), .B(n_401), .Y(n_400) );
INVx4_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_229), .Y(n_248) );
INVx4_ASAP7_75t_L g264 ( .A(n_229), .Y(n_264) );
INVxp67_ASAP7_75t_L g287 ( .A(n_229), .Y(n_287) );
INVx3_ASAP7_75t_L g323 ( .A(n_229), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_230), .B(n_350), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_230), .B(n_405), .Y(n_422) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
INVx1_ASAP7_75t_L g295 ( .A(n_231), .Y(n_295) );
AND2x2_ASAP7_75t_L g404 ( .A(n_231), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR3x1_ASAP7_75t_L g234 ( .A(n_235), .B(n_502), .C(n_570), .Y(n_234) );
NAND3xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_433), .C(n_468), .Y(n_235) );
AOI31xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_344), .A3(n_373), .B(n_387), .Y(n_236) );
OAI21xp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_271), .B(n_299), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_238), .B(n_271), .Y(n_512) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g608 ( .A(n_239), .B(n_472), .Y(n_608) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g542 ( .A(n_240), .B(n_301), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_258), .B(n_265), .Y(n_240) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_241), .A2(n_258), .B(n_265), .Y(n_413) );
NAND3x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_249), .C(n_252), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_246), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_245), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
INVx2_ASAP7_75t_L g340 ( .A(n_245), .Y(n_340) );
INVx2_ASAP7_75t_L g352 ( .A(n_245), .Y(n_352) );
INVx1_ASAP7_75t_L g382 ( .A(n_245), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_248), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g316 ( .A(n_248), .Y(n_316) );
INVx2_ASAP7_75t_SL g357 ( .A(n_248), .Y(n_357) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_249), .A2(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g298 ( .A(n_250), .Y(n_298) );
INVx1_ASAP7_75t_L g378 ( .A(n_250), .Y(n_378) );
BUFx3_ASAP7_75t_L g407 ( .A(n_250), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g260 ( .A(n_255), .Y(n_260) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g278 ( .A(n_257), .Y(n_278) );
INVx2_ASAP7_75t_L g321 ( .A(n_257), .Y(n_321) );
INVx1_ASAP7_75t_L g338 ( .A(n_257), .Y(n_338) );
O2A1O1Ixp5_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_260), .B(n_261), .C(n_264), .Y(n_258) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
INVx2_ASAP7_75t_L g335 ( .A(n_264), .Y(n_335) );
INVx2_ASAP7_75t_L g341 ( .A(n_266), .Y(n_341) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_267), .A2(n_329), .B(n_342), .Y(n_328) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_269), .B(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g343 ( .A(n_269), .Y(n_343) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx3_ASAP7_75t_L g294 ( .A(n_270), .Y(n_294) );
INVx4_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g326 ( .A(n_273), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_SL g471 ( .A(n_273), .Y(n_471) );
AND2x2_ASAP7_75t_L g538 ( .A(n_273), .B(n_412), .Y(n_538) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g440 ( .A(n_274), .Y(n_440) );
INVx3_ASAP7_75t_L g467 ( .A(n_274), .Y(n_467) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_285), .B(n_296), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g356 ( .A(n_284), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_288), .B(n_293), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_286), .A2(n_351), .B1(n_354), .B2(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_290), .B(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx3_ASAP7_75t_L g405 ( .A(n_294), .Y(n_405) );
NOR4xp25_ASAP7_75t_L g379 ( .A(n_297), .B(n_303), .C(n_380), .D(n_385), .Y(n_379) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_298), .B(n_372), .Y(n_371) );
NAND2x1_ASAP7_75t_SL g299 ( .A(n_300), .B(n_326), .Y(n_299) );
AOI211xp5_ASAP7_75t_L g435 ( .A1(n_300), .A2(n_436), .B(n_438), .C(n_441), .Y(n_435) );
AND2x2_ASAP7_75t_L g504 ( .A(n_300), .B(n_480), .Y(n_504) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g432 ( .A(n_301), .B(n_412), .Y(n_432) );
INVx1_ASAP7_75t_L g458 ( .A(n_301), .Y(n_458) );
INVx2_ASAP7_75t_L g465 ( .A(n_301), .Y(n_465) );
OR2x2_ASAP7_75t_L g501 ( .A(n_301), .B(n_412), .Y(n_501) );
AO31x2_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_309), .A3(n_317), .B(n_324), .Y(n_301) );
NOR2x1_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B(n_316), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_316), .A2(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx3_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
BUFx2_ASAP7_75t_L g499 ( .A(n_326), .Y(n_499) );
AND2x2_ASAP7_75t_L g630 ( .A(n_326), .B(n_432), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_326), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g414 ( .A(n_327), .Y(n_414) );
AND2x2_ASAP7_75t_L g481 ( .A(n_327), .B(n_413), .Y(n_481) );
AND2x2_ASAP7_75t_L g546 ( .A(n_327), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI21x1_ASAP7_75t_L g437 ( .A1(n_329), .A2(n_342), .B(n_392), .Y(n_437) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_336), .B(n_341), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_335), .Y(n_330) );
INVx1_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_341), .B(n_347), .Y(n_370) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g461 ( .A(n_345), .Y(n_461) );
OR2x2_ASAP7_75t_L g629 ( .A(n_345), .B(n_495), .Y(n_629) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_360), .Y(n_345) );
AND2x2_ASAP7_75t_L g483 ( .A(n_346), .B(n_453), .Y(n_483) );
INVx1_ASAP7_75t_L g515 ( .A(n_346), .Y(n_515) );
AOI21x1_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_358), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OA21x2_ASAP7_75t_L g391 ( .A1(n_359), .A2(n_392), .B(n_393), .Y(n_391) );
AND2x2_ASAP7_75t_L g390 ( .A(n_360), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g420 ( .A(n_360), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g492 ( .A(n_361), .Y(n_492) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g453 ( .A(n_362), .Y(n_453) );
AOI21x1_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B(n_371), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_370), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_369), .B(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_374), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g394 ( .A(n_375), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g448 ( .A(n_375), .Y(n_448) );
AND2x4_ASAP7_75t_L g484 ( .A(n_375), .B(n_418), .Y(n_484) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_375), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_375), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_379), .Y(n_375) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_376), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g392 ( .A(n_378), .Y(n_392) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_385), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_408), .B1(n_415), .B2(n_428), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_388), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_394), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_390), .B(n_447), .Y(n_463) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
INVx1_ASAP7_75t_L g475 ( .A(n_391), .Y(n_475) );
INVx1_ASAP7_75t_L g586 ( .A(n_391), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_391), .B(n_395), .Y(n_623) );
AOI211xp5_ASAP7_75t_SL g503 ( .A1(n_394), .A2(n_504), .B(n_505), .C(n_516), .Y(n_503) );
AND2x2_ASAP7_75t_L g590 ( .A(n_394), .B(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g569 ( .A(n_395), .Y(n_569) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_SL g419 ( .A(n_396), .Y(n_419) );
AO31x2_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .A3(n_404), .B(n_406), .Y(n_396) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_409), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g456 ( .A(n_411), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g443 ( .A(n_413), .B(n_437), .Y(n_443) );
BUFx2_ASAP7_75t_SL g431 ( .A(n_414), .Y(n_431) );
INVx1_ASAP7_75t_L g521 ( .A(n_414), .Y(n_521) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_414), .Y(n_539) );
AND2x2_ASAP7_75t_L g635 ( .A(n_414), .B(n_465), .Y(n_635) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_416), .B(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_416), .A2(n_634), .B1(n_636), .B2(n_637), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_416), .B(n_558), .Y(n_638) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
OR2x2_ASAP7_75t_L g477 ( .A(n_417), .B(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g460 ( .A(n_418), .B(n_421), .Y(n_460) );
INVx1_ASAP7_75t_L g495 ( .A(n_418), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_418), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2x1_ASAP7_75t_L g452 ( .A(n_419), .B(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g478 ( .A(n_420), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_420), .B(n_451), .Y(n_523) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_421), .B(n_453), .Y(n_531) );
OA21x2_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B(n_427), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x6_ASAP7_75t_L g472 ( .A(n_431), .B(n_457), .Y(n_472) );
AND2x2_ASAP7_75t_L g438 ( .A(n_432), .B(n_439), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_432), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_432), .B(n_594), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_444), .B(n_454), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g466 ( .A(n_437), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g541 ( .A(n_437), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g643 ( .A(n_437), .B(n_547), .Y(n_643) );
AND2x2_ASAP7_75t_L g637 ( .A(n_439), .B(n_443), .Y(n_637) );
INVx2_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g594 ( .A(n_440), .Y(n_594) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g558 ( .A(n_443), .B(n_458), .Y(n_558) );
AND2x4_ASAP7_75t_L g562 ( .A(n_443), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g627 ( .A(n_443), .B(n_614), .Y(n_627) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
AND2x2_ASAP7_75t_L g527 ( .A(n_447), .B(n_450), .Y(n_527) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_448), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g577 ( .A(n_448), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NOR2x1p5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
INVx1_ASAP7_75t_L g543 ( .A(n_451), .Y(n_543) );
INVx2_ASAP7_75t_L g592 ( .A(n_451), .Y(n_592) );
INVx1_ASAP7_75t_L g566 ( .A(n_453), .Y(n_566) );
AO22x1_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_459), .B1(n_462), .B2(n_464), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_455), .A2(n_525), .B1(n_532), .B2(n_537), .C(n_540), .Y(n_524) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_458), .B(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_458), .Y(n_581) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AND2x2_ASAP7_75t_L g536 ( .A(n_460), .B(n_483), .Y(n_536) );
AND2x2_ASAP7_75t_L g636 ( .A(n_460), .B(n_565), .Y(n_636) );
AND2x2_ASAP7_75t_L g644 ( .A(n_460), .B(n_592), .Y(n_644) );
AND2x4_ASAP7_75t_L g610 ( .A(n_461), .B(n_484), .Y(n_610) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g557 ( .A(n_465), .Y(n_557) );
INVx1_ASAP7_75t_L g563 ( .A(n_465), .Y(n_563) );
INVx1_ASAP7_75t_L g597 ( .A(n_465), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_465), .B(n_547), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_465), .B(n_481), .Y(n_615) );
INVx1_ASAP7_75t_L g488 ( .A(n_466), .Y(n_488) );
INVx2_ASAP7_75t_L g547 ( .A(n_467), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_467), .B(n_557), .Y(n_556) );
AOI211xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_473), .B(n_479), .C(n_485), .Y(n_468) );
NOR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g480 ( .A(n_471), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g508 ( .A(n_471), .Y(n_508) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_471), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_471), .B(n_580), .Y(n_619) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g560 ( .A(n_475), .Y(n_560) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g513 ( .A(n_478), .B(n_514), .Y(n_513) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_478), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
AND2x2_ASAP7_75t_L g507 ( .A(n_481), .B(n_508), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_482), .B(n_574), .C(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_483), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_484), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_491), .Y(n_534) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
OAI22xp33_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_489), .B1(n_496), .B2(n_498), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g578 ( .A(n_492), .Y(n_578) );
AND2x2_ASAP7_75t_L g604 ( .A(n_492), .B(n_515), .Y(n_604) );
INVx1_ASAP7_75t_L g626 ( .A(n_492), .Y(n_626) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_494), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g603 ( .A(n_495), .B(n_604), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g575 ( .A(n_501), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_524), .C(n_550), .Y(n_502) );
OAI22xp33_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_509), .B1(n_512), .B2(n_513), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
INVx1_ASAP7_75t_L g530 ( .A(n_514), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_522), .Y(n_516) );
INVxp33_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_521), .B(n_538), .Y(n_602) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g553 ( .A(n_523), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_529), .A2(n_584), .B1(n_612), .B2(n_615), .Y(n_611) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_530), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_536), .A2(n_640), .B1(n_643), .B2(n_644), .Y(n_639) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_543), .B(n_544), .C(n_548), .Y(n_540) );
OR2x2_ASAP7_75t_L g544 ( .A(n_542), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g634 ( .A(n_547), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_554), .B1(n_558), .B2(n_559), .C(n_561), .Y(n_550) );
AND2x2_ASAP7_75t_L g631 ( .A(n_551), .B(n_601), .Y(n_631) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_562), .A2(n_601), .B1(n_603), .B2(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g642 ( .A(n_563), .Y(n_642) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g584 ( .A(n_569), .B(n_585), .Y(n_584) );
NAND3xp33_ASAP7_75t_SL g570 ( .A(n_571), .B(n_587), .C(n_616), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B1(n_581), .B2(n_582), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_574), .A2(n_618), .B(n_620), .Y(n_617) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g599 ( .A(n_585), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_606), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_593), .B1(n_595), .B2(n_598), .C(n_600), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_631), .C(n_632), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_627), .B1(n_628), .B2(n_630), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND4xp25_ASAP7_75t_SL g632 ( .A(n_633), .B(n_638), .C(n_639), .D(n_645), .Y(n_632) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_643), .Y(n_646) );
OAI222xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B1(n_653), .B2(n_656), .C1(n_658), .C2(n_662), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_649), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_663), .Y(n_662) );
endmodule