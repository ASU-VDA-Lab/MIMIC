module fake_jpeg_21424_n_67 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_33),
.B1(n_29),
.B2(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_41),
.B1(n_37),
.B2(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_1),
.B1(n_7),
.B2(n_10),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_12),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_34),
.B1(n_32),
.B2(n_5),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_34),
.B(n_3),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_51),
.B(n_53),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_34),
.B1(n_3),
.B2(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_11),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_56),
.C(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_53),
.B(n_54),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_61),
.B(n_57),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_55),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_44),
.A3(n_48),
.B1(n_19),
.B2(n_20),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_66),
.B(n_23),
.Y(n_67)
);


endmodule